// Benchmark "c5315" written by ABC on Thu Mar  5 01:07:35 2020

module c5315 ( 
    G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
    G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
    G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
    G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140,
    G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173,
    G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209,
    G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251,
    G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293,
    G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338,
    G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389,
    G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523,
    G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691,
    G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717,
    G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34,
    G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76,
    G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103,
    G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
    G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137,
    G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170,
    G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206,
    G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248,
    G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292,
    G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335,
    G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386,
    G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514,
    G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690,
    G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552,
    G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire G4114, G2825, G3547, G3549, G3551, G3553, G633, G814, G816, G844,
    G846, G852, G1502, G1528, G1552, G1609, G1633, G1697, G1698, G1701,
    G2179, G2203, G2226, G2281, G2304, G2361, G2370, G2382, G2393, G2405,
    G2418, G2442, G2476, G2500, G2533, G2537, G2541, G2545, G2549, G2553,
    G2557, G2561, G2627, G2631, G2635, G2639, G2643, G2647, G2651, G2655,
    G2721, G2734, G2816, G2822, G2826, G2828, G2882, G2886, G2890, G2894,
    G2898, G2902, G2948, G2952, G2956, G2960, G2964, G2968, G3024, G3028,
    G3032, G3036, G3040, G3044, G3048, G3052, G3092, G3105, G3175, G3176,
    G3181, G3204, G3208, G3212, G3216, G3220, G3224, G3256, G3260, G3264,
    G3268, G3272, G3276, G3302, G3314, G3354, G3358, G3362, G3366, G3370,
    G3374, G3378, G3382, G3440, G3554, G3555, G3556, G3558, G3582, G3616,
    G3628, G3660, G3684, G3721, G3728, G3737, G3757, G3795, G3815, G3972,
    G3991, G4030, G4049, G4110, G4119, G4127, G4135, G4143, G4151, G4159,
    G4167, G4175, G4183, G4188, G4276, G4284, G4292, G4300, G4308, G4316,
    G4324, G4332, G4340, G4631, G4639, G4647, G4655, G4663, G4671, G4676,
    G4764, G4772, G4780, G4788, G4796, G4804, G5082, G5085, G5090, G5093,
    G5098, G5101, G5108, G5111, G5332, G5335, G5340, G5343, G5348, G5351,
    G5356, G5359, G5369, G2979, G2999, G1580, G1586, G1592, G1598, G1604,
    G1668, G1674, G1680, G1686, G2254, G2260, G2266, G2272, G2278, G2339,
    G2345, G2351, G2357, G711, G721, G726, G731, G736, G741, G746, G751,
    G756, G761, G766, G771, G776, G781, G786, G791, G796, G801, G806,
    G3734, G842, G858, G881, G4123, G4131, G4139, G4147, G4155, G4163,
    G4171, G4179, G4187, G4194, G4282, G4290, G4298, G4306, G4314, G4322,
    G4330, G4338, G4346, G1526, G1540, G1564, G1606, G1621, G1645, G1661,
    G1688, G4635, G4643, G4651, G4659, G4667, G4675, G4682, G4770, G4778,
    G4786, G4794, G4802, G4810, G2202, G2215, G2238, G2279, G2293, G2316,
    G2332, G2430, G2454, G2488, G2512, G2536, G2540, G2544, G2548, G2552,
    G2556, G2560, G2564, G2566, G2572, G2578, G2584, G2590, G2595, G2600,
    G2605, G2630, G2634, G2638, G2642, G2646, G2650, G2654, G2658, G2660,
    G2666, G2672, G2678, G2684, G2689, G2694, G2699, G2728, G2741, G2748,
    G2750, G2752, G2754, G2756, G2758, G2760, G2762, G2764, G2766, G2827,
    G2838, G2847, G2885, G2889, G2893, G2897, G2901, G2905, G2906, G2909,
    G2913, G2918, G2922, G2927, G2951, G2955, G2959, G2963, G2967, G2971,
    G2973, G2980, G2982, G2988, G2994, G3001, G3006, G3027, G3031, G3035,
    G3039, G3043, G3047, G3051, G3055, G3056, G3060, G3064, G3068, G3073,
    G3078, G3083, G3088, G3099, G3112, G3119, G3121, G3123, G3125, G3126,
    G3128, G3130, G3132, G3134, G3136, G3187, G3193, G3196, G3199, G3202,
    G3207, G3211, G3215, G3219, G3223, G3227, G3228, G3232, G3234, G3238,
    G3243, G3247, G3249, G3253, G3259, G3263, G3267, G3271, G3275, G3279,
    G3280, G3283, G3287, G3292, G3295, G3299, G3305, G3306, G3310, G3317,
    G3318, G3322, G3326, G3333, G3357, G3361, G3365, G3369, G3373, G3377,
    G3381, G3385, G3386, G3390, G3394, G3398, G3403, G3408, G3413, G3418,
    G5088, G5089, G5096, G5097, G3489, G3493, G3570, G3594, G3622, G3632,
    G3637, G3640, G3643, G3646, G3672, G3696, G3745, G3765, G3803, G3823,
    G5338, G5339, G5346, G5347, G5354, G5355, G3979, G3998, G4037, G4056,
    G4094, G5104, G5105, G5114, G5115, G5362, G5363, G5366, G5373, G2568,
    G2574, G2580, G2586, G2592, G2597, G2602, G2607, G2662, G2668, G2674,
    G2680, G2686, G2691, G2696, G2701, G2907, G2910, G2914, G2920, G2924,
    G2929, G2975, G2984, G2990, G2996, G3003, G3008, G3015, G3057, G3061,
    G3065, G3069, G3075, G3080, G3085, G3090, G3229, G3233, G3235, G3239,
    G3244, G3250, G3254, G3281, G3284, G3288, G3293, G3296, G3300, G3327,
    G3334, G3387, G3391, G3395, G3399, G3405, G3410, G3415, G3420, G3422,
    G3423, G3431, G3432, G3895, G3896, G3904, G3905, G3913, G3914, G5106,
    G5107, G5116, G5117, G5364, G5365, G2880, G2881, G1579, G1585, G1591,
    G1597, G1603, G1667, G1673, G1679, G1685, G2876, G2877, G2253, G2259,
    G2265, G2271, G2277, G2338, G2344, G2350, G2356, G2868, G2869, G710,
    G2872, G2873, G720, G725, G730, G735, G740, G745, G750, G755, G760,
    G765, G770, G775, G780, G785, G790, G795, G800, G805, G841, G857, G880,
    G1660, G2331, G2569, G2575, G2581, G2587, G2593, G2598, G2603, G2608,
    G2663, G2669, G2675, G2681, G2687, G2692, G2697, G2702, G2747, G2749,
    G2751, G2753, G2755, G2757, G2759, G2761, G2763, G2765, G2857, G2908,
    G2911, G2915, G2925, G2930, G2933, G2976, G2985, G2991, G2997, G3004,
    G3009, G3058, G3062, G3066, G3070, G3076, G3081, G3086, G3091, G3118,
    G3120, G3122, G3124, G3127, G3129, G3131, G3133, G3135, G3147, G3192,
    G3195, G3198, G3201, G3230, G3236, G3240, G3245, G3251, G3255, G3282,
    G3285, G3289, G3297, G3301, G3309, G3313, G3321, G3325, G3328, G3329,
    G3335, G3336, G3341, G3345, G3388, G3392, G3396, G3400, G3406, G3411,
    G3416, G3421, G3424, G3433, G3492, G3496, G3780, G3783, G3786, G3789,
    G3838, G3841, G3844, G3847, G3897, G3906, G3915, G4011, G4014, G4017,
    G4020, G4023, G4069, G4072, G4075, G4078, G4081, G5206, G5209, G5307,
    G5322, G5372, G5375, G5399, G2813, G3197, G3200, G3203, G3194, G2570,
    G2576, G2582, G2588, G2664, G2670, G2676, G2682, G2767, G2772, G2776,
    G2780, G2784, G2788, G2794, G2798, G2802, G2912, G2916, G2936, G2977,
    G2986, G2992, G3059, G3063, G3067, G3071, G3137, G3139, G3143, G3151,
    G3155, G3161, G3165, G3167, G3231, G3237, G3241, G3286, G3290, G3330,
    G3337, G3342, G3346, G3348, G3352, G3389, G3393, G3397, G3401, G3845,
    G5126, G5178, G5325, G5374, G2810, G635, G2878, G2879, G2874, G2875,
    G703, G2866, G2867, G2870, G2871, G716, G819, G1789, G2036, G2611,
    G2615, G2619, G2623, G2705, G2709, G2713, G2717, G2939, G2942, G2945,
    G3012, G3018, G3021, G3331, G3338, G3343, G3347, G3428, G3437, G3514,
    G3836, G3852, G5311, G3901, G3910, G3934, G3938, G4652, G4783, G5137,
    G5212, G5213, G5260, G5263, G5268, G5271, G5276, G5279, G5289, G5296,
    G5299, G5304, G5312, G5315, G5328, G5396, G5403, G1286, G2809, G597,
    G1031, G637, G671, G705, G713, G1046, G1064, G1071, G1097, G1111,
    G1128, G1145, G1160, G1301, G1318, G1324, G1341, G1359, G1382, G1404,
    G1412, G1704, G1712, G1724, G1742, G1749, G1775, G1806, G1823, G1829,
    G1837, G1958, G1966, G1978, G1995, G2001, G2018, G2059, G2081, G2089,
    G2106, G3170, G3332, G3339, G5132, G5184, G3853, G3874, G4076, G4116,
    G4124, G4132, G4140, G4148, G4156, G4164, G4172, G4180, G4228, G4279,
    G4287, G4295, G4303, G4311, G4319, G4327, G4335, G4343, G4348, G4464,
    G4628, G4636, G4644, G4660, G4668, G4716, G4767, G4775, G4791, G4799,
    G4807, G4812, G5118, G5121, G5129, G5134, G5142, G5145, G5152, G5155,
    G5162, G5165, G5170, G5173, G5181, G5186, G5189, G5196, G5199, G5214,
    G5215, G5329, G5330, G2807, G2808, G2811, G2812, G2814, G2626, G2622,
    G2618, G2614, G2720, G2716, G2712, G2708, G3731, G4658, G1777, G2019,
    G4787, G3350, G3353, G5141, G3513, G3516, G3517, G3778, G3781, G3784,
    G3787, G3839, G3842, G5266, G5267, G5274, G5275, G5302, G5303, G5310,
    G3891, G3937, G3941, G3955, G3958, G4009, G4012, G4015, G4018, G4067,
    G4070, G4073, G4079, G5239, G5282, G5283, G5293, G5318, G5319, G5331,
    G5402, G5405, G595, G596, G607, G608, G1845, G1846, G2115, G2116,
    G4122, G1022, G4130, G1033, G4138, G1051, G4146, G1079, G4154, G1088,
    G4162, G1099, G4170, G1115, G4178, G1133, G4186, G1151, G4234, G1276,
    G4283, G1287, G4291, G1305, G4299, G1330, G4307, G1342, G4315, G1363,
    G4323, G1388, G4331, G1420, G4339, G1428, G4347, G4634, G1729, G4642,
    G1757, G4650, G1766, G1776, G4666, G1793, G4674, G1811, G1849, G1852,
    G1875, G4722, G1982, G4771, G2007, G4779, G2020, G2040, G4795, G2065,
    G4803, G2097, G4811, G2119, G2122, G5124, G5125, G3452, G5133, G5140,
    G3462, G5168, G5169, G5176, G5177, G3484, G5185, G3515, G3518, G3857,
    G3860, G3861, G3869, G3870, G3878, G3881, G3882, G3890, G3954, G3957,
    G4021, G4099, G4236, G4354, G4406, G4470, G4552, G4679, G4687, G4695,
    G4703, G4711, G4724, G4818, G4855, G4865, G4870, G4913, G4923, G4951,
    G5006, G5039, G5148, G5149, G5158, G5159, G5192, G5193, G5202, G5203,
    G5284, G5285, G5320, G5321, G5386, G5404, G609, G1021, G1032, G1050,
    G1078, G1087, G1098, G1114, G1132, G1150, G1277, G1288, G1306, G1331,
    G1343, G1364, G1389, G1421, G1429, G1728, G1756, G1765, G1778, G1792,
    G1810, G1983, G2008, G2021, G2041, G2066, G2098, G3443, G3444, G3453,
    G3461, G3466, G3467, G3475, G3476, G3485, G5243, G3862, G3871, G3883,
    G3892, G3956, G3959, G4756, G5150, G5151, G5160, G5161, G5194, G5195,
    G5204, G5205, G5236, G5286, G5379, G5389, G5425, G1023, G1034, G1052,
    G1080, G1089, G1100, G1116, G1134, G1152, G4242, G1278, G1289, G1307,
    G1332, G1344, G1365, G1390, G1422, G1430, G1730, G1758, G1767, G1794,
    G1812, G1876, G4683, G4691, G4699, G4707, G4715, G4730, G1984, G2009,
    G2042, G2067, G2099, G4869, G4927, G3445, G3454, G3463, G3468, G3477,
    G3486, G4103, G4412, G4558, G4859, G4876, G4917, G4955, G5012, G5043,
    G5216, G5219, G5226, G5229, G5392, G5422, G1866, G1877, G4762, G2142,
    G2146, G5242, G3532, G3866, G3887, G3918, G3922, G3926, G3930, G5429,
    G4104, G4743, G4991, G5001, G5292, G5295, G5383, G5393, G5394, G1439,
    G1440, G1441, G1847, G1168, G1169, G1170, G2117, G1086, G1166, G1171,
    G1172, G1173, G1174, G1175, G1176, G1177, G1178, G1179, G1181, G1182,
    G1183, G1184, G1188, G1189, G1190, G1191, G1192, G1193, G1194, G1195,
    G1196, G1197, G1437, G1442, G1443, G1444, G1445, G1446, G1447, G1451,
    G1454, G1455, G1456, G1457, G1465, G1466, G1467, G1468, G1469, G1470,
    G1471, G1472, G1473, G1474, G1475, G1476, G1477, G1481, G1482, G1764,
    G1843, G1850, G1851, G1853, G1854, G1855, G1856, G1857, G1859, G1860,
    G1861, G1862, G1867, G1868, G1869, G1870, G1871, G1872, G1873, G1874,
    G1878, G2113, G2120, G2121, G2123, G2124, G2128, G2131, G2132, G2133,
    G2134, G2143, G2144, G2145, G2147, G2148, G2149, G2150, G2151, G2152,
    G2153, G2154, G2158, G2159, G3449, G3458, G3472, G3481, G3497, G3501,
    G3505, G3509, G3531, G5428, G3967, G4191, G4199, G4207, G4215, G4223,
    G4231, G4239, G4247, G4255, G4263, G4271, G4371, G4381, G4391, G4401,
    G4429, G4439, G4449, G4459, G4497, G4507, G4517, G4527, G4537, G4547,
    G4585, G4595, G4605, G4615, G4719, G4727, G4735, G4751, G4759, G4835,
    G4845, G4893, G4903, G4961, G4971, G4981, G5049, G5059, G5069, G5222,
    G5223, G5232, G5233, G5294, G5395, G589, G616, G619, G627, G1185,
    G1448, G1458, G1478, G1863, G4747, G2125, G2135, G2155, G4995, G5005,
    G3533, G3921, G3925, G3929, G3933, G3943, G3946, G3949, G3952, G3966,
    G4107, G4196, G4204, G4212, G4220, G4244, G4252, G4260, G4268, G4361,
    G4419, G4467, G4487, G4555, G4575, G4684, G4692, G4700, G4708, G4732,
    G4740, G4748, G4825, G4883, G4928, G4941, G5009, G5029, G5224, G5225,
    G5234, G5235, G5376, G5417, G576, G1198, G4195, G4203, G4211, G4219,
    G4227, G1217, G4235, G1221, G4243, G1224, G4251, G4259, G4267, G4275,
    G1453, G4405, G4463, G4541, G4551, G1895, G4723, G1899, G4731, G1902,
    G4739, G4755, G1929, G4763, G2130, G3500, G3504, G3508, G3512, G3520,
    G3523, G3526, G3529, G3837, G3942, G3945, G3948, G3951, G3968, G4375,
    G4385, G4395, G4433, G4443, G4453, G4501, G4511, G4521, G4531, G4619,
    G4589, G4599, G4609, G4839, G4849, G4897, G4907, G4965, G4975, G4985,
    G5073, G5053, G5063, G5247, G5255, G590, G617, G620, G628, G3535,
    G1199, G4202, G1204, G4210, G1207, G4218, G1211, G4226, G1214, G1218,
    G1222, G1225, G4250, G1237, G4258, G1242, G4266, G1247, G4274, G1252,
    G1462, G4690, G1882, G4698, G1885, G4706, G1889, G4714, G1892, G1896,
    G1900, G1903, G4738, G1915, G4746, G1920, G4754, G1925, G1930, G2139,
    G3519, G3522, G3525, G3528, G3848, G3944, G3947, G3950, G3953, G5421,
    G4111, G4112, G4351, G4365, G4409, G4423, G4471, G4472, G4477, G4491,
    G4559, G4560, G4565, G4579, G4815, G4829, G4873, G4887, G4931, G4934,
    G4945, G5013, G5014, G5019, G5033, G5382, G5385, G3970, G1200, G1203,
    G1206, G1210, G1213, G1219, G1223, G1236, G1241, G1246, G1251, G1881,
    G1884, G1888, G1891, G1897, G1901, G1914, G1919, G1924, G1931, G3521,
    G3524, G3527, G3530, G5251, G5259, G4113, G4473, G4561, G5015, G5384,
    G5406, G5414, G1664, G2335, G718, G855, G1205, G1208, G1212, G1215,
    G1220, G1231, G1238, G1243, G1248, G1253, G1272, G1483, G1883, G1886,
    G1890, G1893, G1898, G1909, G1916, G1921, G1926, G1953, G2160, G4355,
    G4356, G4413, G4414, G4474, G4481, G4562, G4569, G4819, G4820, G4877,
    G4878, G4935, G4936, G5016, G5023, G5244, G5252, G5409, G566, G577,
    G3733, G1209, G1216, G1257, G1262, G1267, G1887, G1894, G1935, G1943,
    G1948, G3779, G3840, G5412, G5420, G3964, G4357, G4415, G4821, G4879,
    G4937, G567, G568, G569, G570, G578, G579, G580, G1256, G1261, G1266,
    G1271, G1486, G1934, G1942, G1947, G1952, G2163, G5250, G3537, G5258,
    G3542, G3782, G3785, G3788, G3790, G3843, G3846, G3849, G3960, G5413,
    G3963, G4010, G4068, G4358, G4416, G4480, G4483, G4568, G4571, G4822,
    G4880, G4938, G5022, G5025, G1258, G1263, G1268, G1273, G1936, G1944,
    G1949, G1954, G3536, G3541, G3791, G3792, G3793, G3850, G3851, G3961,
    G3965, G4024, G4082, G4482, G4570, G5024, G1666, G1670, G2337, G2341,
    G719, G758, G798, G856, G3538, G3543, G3962, G4364, G4367, G4422,
    G4425, G4484, G4572, G4828, G4831, G4886, G4889, G4944, G4947, G5026,
    G571, G572, G573, G574, G581, G582, G583, G584, G1576, G1578, G659,
    G1672, G1676, G1678, G1682, G1684, G2250, G2252, G691, G2343, G2347,
    G2349, G2353, G2355, G743, G744, G748, G749, G753, G754, G759, G783,
    G784, G788, G789, G793, G794, G799, G3735, G3835, G3651, G4013, G4016,
    G4019, G4022, G4071, G4074, G4077, G4080, G4096, G4366, G4424, G4830,
    G4888, G4946, G640, G662, G665, G668, G674, G694, G697, G700, G817,
    G839, G3540, G3545, G3777, G3648, G4025, G4026, G4027, G4028, G4083,
    G4084, G4085, G4086, G4368, G4426, G4490, G4493, G4578, G4581, G4832,
    G4890, G4948, G5032, G5035, G811, G812, G853, G878, G4492, G4580,
    G5034, G1582, G1584, G1588, G1590, G1594, G1596, G1600, G1602, G2256,
    G2258, G2262, G2264, G2268, G2270, G2274, G2276, G708, G709, G723,
    G724, G728, G729, G733, G734, G738, G739, G768, G769, G773, G774, G778,
    G779, G4374, G4377, G4432, G4435, G4494, G4582, G4838, G4841, G4896,
    G4899, G4954, G4957, G5036, G643, G646, G649, G652, G677, G680, G683,
    G686, G4376, G4434, G4840, G4898, G4956, G4378, G4436, G4500, G4503,
    G4588, G4591, G4842, G4900, G4958, G5042, G5045, G4502, G4590, G5044,
    G4384, G4387, G4442, G4445, G4504, G4592, G4848, G4851, G4906, G4909,
    G4964, G4967, G5046, G4386, G4444, G4850, G4908, G4966, G4388, G4446,
    G4510, G4513, G4598, G4601, G4852, G4910, G4968, G5052, G5055, G4512,
    G4600, G5054, G4394, G4397, G4452, G4455, G4514, G4602, G4858, G4861,
    G4916, G4919, G4974, G4977, G5056, G4396, G4454, G4860, G4918, G4976,
    G4398, G4456, G4520, G4523, G4608, G4611, G4862, G4920, G4978, G5062,
    G5065, G4522, G4610, G5064, G4404, G1488, G4462, G1493, G4868, G2165,
    G4926, G2170, G4524, G4612, G4984, G4987, G5066, G1487, G1492, G2164,
    G2169, G4986, G1489, G1494, G2166, G2171, G4530, G4533, G4618, G4543,
    G4988, G5072, G4997, G4532, G4542, G4996, G1513, G1514, G1515, G1516,
    G4994, G2184, G2190, G2191, G2192, G2193, G4534, G4544, G4998, G2183,
    G4620, G5074, G4540, G1507, G4550, G1510, G2185, G5004, G2187, G1506,
    G1509, G4626, G2186, G2195, G5080, G1508, G1511, G2188, G1512, G1518,
    G2189, G1517, G2194, G4623, G5077, G1519, G4627, G2196, G5081, G1520,
    G2197, G1521, G2198, G840, G879, G1524, G2201, G3649, G3652, G3657,
    G3658, G3636, G3639, G3642, G3645, G3653, G3654, G3655, G3656, G763,
    G764, G803, G804, G1657, G1659, G2328, G2330, G1662, G2333, G657, G689;
  assign G144 = G141;
  assign G298 = G293;
  assign G4114 = G135 & G4115;
  assign G2825 = ~G2824;
  assign G973 = G3173;
  assign G3547 = ~G3546;
  assign G3549 = ~G3548;
  assign G3551 = ~G3550;
  assign G3553 = ~G3552;
  assign G594 = ~G545;
  assign G599 = ~G348;
  assign G600 = ~G366;
  assign G601 = G552 & G562;
  assign G602 = ~G549;
  assign G603 = ~G545;
  assign G604 = ~G545;
  assign G611 = ~G338;
  assign G612 = ~G358;
  assign G633 = ~G373 | ~G1;
  assign G810 = G141 & G145;
  assign G814 = ~G3173;
  assign G816 = ~G4114;
  assign G844 = G2825 & G27;
  assign G846 = G386 & G556;
  assign G848 = ~G245;
  assign G849 = ~G552;
  assign G850 = ~G562;
  assign G851 = ~G559;
  assign G852 = G552 & G556 & G386 & G559;
  assign G1502 = ~G1497;
  assign G1528 = G1689;
  assign G1552 = G1690;
  assign G1609 = G1689;
  assign G1633 = G1690;
  assign G1697 = G137;
  assign G1698 = G137;
  assign G1701 = G141;
  assign G2179 = ~G2174;
  assign G2203 = G1691;
  assign G2226 = G1694;
  assign G2281 = G1691;
  assign G2304 = G1694;
  assign G2361 = G254;
  assign G2370 = G251;
  assign G2382 = G251;
  assign G2393 = G248;
  assign G2405 = G248;
  assign G2418 = G4088;
  assign G2442 = G4087;
  assign G2476 = G4089;
  assign G2500 = G4090;
  assign G2533 = G210;
  assign G2537 = G210;
  assign G2541 = G218;
  assign G2545 = G218;
  assign G2549 = G226;
  assign G2553 = G226;
  assign G2557 = G234;
  assign G2561 = G234;
  assign G2627 = G257;
  assign G2631 = G257;
  assign G2635 = G265;
  assign G2639 = G265;
  assign G2643 = G273;
  assign G2647 = G273;
  assign G2651 = G281;
  assign G2655 = G281;
  assign G2721 = G335;
  assign G2734 = G335;
  assign G2816 = G206;
  assign G2822 = G27 & G31;
  assign G2826 = G1;
  assign G2828 = G2358;
  assign G2882 = G293;
  assign G2886 = G302;
  assign G2890 = G308;
  assign G2894 = G308;
  assign G2898 = G316;
  assign G2902 = G316;
  assign G2948 = G324;
  assign G2952 = G324;
  assign G2956 = G341;
  assign G2960 = G341;
  assign G2964 = G351;
  assign G2968 = G351;
  assign G3024 = G257;
  assign G3028 = G257;
  assign G3032 = G265;
  assign G3036 = G265;
  assign G3040 = G273;
  assign G3044 = G273;
  assign G3048 = G281;
  assign G3052 = G281;
  assign G3092 = G332;
  assign G3105 = G332;
  assign G3175 = G549;
  assign G3176 = G31 & G27;
  assign G3181 = ~G2358;
  assign G3204 = G324;
  assign G3208 = G324;
  assign G3212 = G341;
  assign G3216 = G341;
  assign G3220 = G351;
  assign G3224 = G351;
  assign G3256 = G293;
  assign G3260 = G302;
  assign G3264 = G308;
  assign G3268 = G308;
  assign G3272 = G316;
  assign G3276 = G316;
  assign G3302 = G361;
  assign G3314 = G361;
  assign G3354 = G210;
  assign G3358 = G210;
  assign G3362 = G218;
  assign G3366 = G218;
  assign G3370 = G226;
  assign G3374 = G226;
  assign G3378 = G234;
  assign G3382 = G234;
  assign G3440 = ~G324;
  assign G3554 = G242;
  assign G3555 = G242;
  assign G3556 = G254;
  assign G3558 = G4088;
  assign G3582 = G4087;
  assign G3616 = G4092;
  assign G3628 = G4091;
  assign G3660 = G4089;
  assign G3684 = G4090;
  assign G3721 = ~G3717;
  assign G3728 = ~G3724;
  assign G3737 = G4091;
  assign G3757 = G4092;
  assign G3795 = G4091;
  assign G3815 = G4092;
  assign G3972 = G4091;
  assign G3991 = G4092;
  assign G4030 = G4091;
  assign G4049 = G4092;
  assign G4110 = G299;
  assign G4119 = G446;
  assign G4127 = G457;
  assign G4135 = G468;
  assign G4143 = G422;
  assign G4151 = G435;
  assign G4159 = G389;
  assign G4167 = G400;
  assign G4175 = G411;
  assign G4183 = G374;
  assign G4188 = G4;
  assign G4276 = G446;
  assign G4284 = G457;
  assign G4292 = G468;
  assign G4300 = G435;
  assign G4308 = G389;
  assign G4316 = G400;
  assign G4324 = G411;
  assign G4332 = G422;
  assign G4340 = G374;
  assign G4631 = G479;
  assign G4639 = G490;
  assign G4647 = G503;
  assign G4655 = G514;
  assign G4663 = G523;
  assign G4671 = G534;
  assign G4676 = G54;
  assign G4764 = G479;
  assign G4772 = G503;
  assign G4780 = G514;
  assign G4788 = G523;
  assign G4796 = G534;
  assign G4804 = G490;
  assign G5082 = G361;
  assign G5085 = G369;
  assign G5090 = G341;
  assign G5093 = G351;
  assign G5098 = G308;
  assign G5101 = G316;
  assign G5108 = G293;
  assign G5111 = G302;
  assign G5332 = G281;
  assign G5335 = G289;
  assign G5340 = G265;
  assign G5343 = G273;
  assign G5348 = G234;
  assign G5351 = G257;
  assign G5356 = G218;
  assign G5359 = G226;
  assign G5369 = G210;
  assign G634 = ~G633;
  assign G815 = G136 & G814;
  assign G845 = ~G844;
  assign G847 = ~G846;
  assign G926 = G1697;
  assign G923 = G1701;
  assign G921 = G2826;
  assign G2979 = G3553 & G514;
  assign G2999 = G3547 | G514;
  assign G892 = G3175;
  assign G887 = G4110;
  assign G606 = ~G3175;
  assign G1580 = G1552 & G170 & G1528;
  assign G1586 = G1552 & G173 & G1528;
  assign G1592 = G1552 & G167 & G1528;
  assign G1598 = G1552 & G164 & G1528;
  assign G1604 = G1552 & G161 & G1528;
  assign G656 = ~G2822 | ~G140;
  assign G1668 = G1633 & G185 & G1609;
  assign G1674 = G1633 & G158 & G1609;
  assign G1680 = G1633 & G152 & G1609;
  assign G1686 = G1633 & G146 & G1609;
  assign G2254 = G2226 & G170 & G2203;
  assign G2260 = G2226 & G173 & G2203;
  assign G2266 = G2226 & G167 & G2203;
  assign G2272 = G2226 & G164 & G2203;
  assign G2278 = G2226 & G161 & G2203;
  assign G2339 = G2304 & G185 & G2281;
  assign G2345 = G2304 & G158 & G2281;
  assign G2351 = G2304 & G152 & G2281;
  assign G2357 = G2304 & G146 & G2281;
  assign G711 = G3684 & G106 & G3660;
  assign G721 = G2442 & G61 & G2418;
  assign G726 = G3582 & G106 & G3558;
  assign G731 = G3582 & G49 & G3558;
  assign G736 = G3582 & G103 & G3558;
  assign G741 = G3582 & G40 & G3558;
  assign G746 = G3582 & G37 & G3558;
  assign G751 = G2442 & G20 & G2418;
  assign G756 = G2442 & G17 & G2418;
  assign G761 = G2442 & G70 & G2418;
  assign G766 = G2442 & G64 & G2418;
  assign G771 = G3684 & G49 & G3660;
  assign G776 = G3684 & G103 & G3660;
  assign G781 = G3684 & G40 & G3660;
  assign G786 = G3684 & G37 & G3660;
  assign G791 = G2500 & G20 & G2476;
  assign G796 = G2500 & G17 & G2476;
  assign G801 = G2500 & G70 & G2476;
  assign G806 = G2500 & G64 & G2476;
  assign G809 = ~G2822;
  assign G3734 = G3717 & G123 & G3728;
  assign G842 = G3795 & G3815;
  assign G858 = G2500 & G61 & G2476;
  assign G881 = G3737 & G3757;
  assign G4123 = ~G4119;
  assign G4131 = ~G4127;
  assign G4139 = ~G4135;
  assign G4147 = ~G4143;
  assign G4155 = ~G4151;
  assign G4163 = ~G4159;
  assign G4171 = ~G4167;
  assign G4179 = ~G4175;
  assign G4187 = ~G4183;
  assign G4194 = ~G4188;
  assign G4282 = ~G4276;
  assign G4290 = ~G4284;
  assign G4298 = ~G4292;
  assign G4306 = ~G4300;
  assign G4314 = ~G4308;
  assign G4322 = ~G4316;
  assign G4330 = ~G4324;
  assign G4338 = ~G4332;
  assign G4346 = ~G4340;
  assign G1526 = G1697;
  assign G1540 = ~G1528;
  assign G1564 = ~G1552;
  assign G1606 = G1697;
  assign G1621 = ~G1609;
  assign G1645 = ~G1633;
  assign G1661 = G1633 & G179 & G1609;
  assign G1688 = G2826;
  assign G4635 = ~G4631;
  assign G4643 = ~G4639;
  assign G4651 = ~G4647;
  assign G4659 = ~G4655;
  assign G4667 = ~G4663;
  assign G4675 = ~G4671;
  assign G4682 = ~G4676;
  assign G4770 = ~G4764;
  assign G4778 = ~G4772;
  assign G4786 = ~G4780;
  assign G4794 = ~G4788;
  assign G4802 = ~G4796;
  assign G4810 = ~G4804;
  assign G2202 = G1698;
  assign G2215 = ~G2203;
  assign G2238 = ~G2226;
  assign G2279 = G1698;
  assign G2293 = ~G2281;
  assign G2316 = ~G2304;
  assign G2332 = G2304 & G179 & G2281;
  assign G2430 = ~G2418;
  assign G2454 = ~G2442;
  assign G2488 = ~G2476;
  assign G2512 = ~G2500;
  assign G2536 = ~G2533;
  assign G2540 = ~G2537;
  assign G2544 = ~G2541;
  assign G2548 = ~G2545;
  assign G2552 = ~G2549;
  assign G2556 = ~G2553;
  assign G2560 = ~G2557;
  assign G2564 = ~G2561;
  assign G2566 = G2537 & G3553 & G457;
  assign G2572 = G2545 & G3553 & G468;
  assign G2578 = G2553 & G3553 & G422;
  assign G2584 = G2561 & G3553 & G435;
  assign G2590 = G3547 & G2533;
  assign G2595 = G3547 & G2541;
  assign G2600 = G3547 & G2549;
  assign G2605 = G3547 & G2557;
  assign G2630 = ~G2627;
  assign G2634 = ~G2631;
  assign G2638 = ~G2635;
  assign G2642 = ~G2639;
  assign G2646 = ~G2643;
  assign G2650 = ~G2647;
  assign G2654 = ~G2651;
  assign G2658 = ~G2655;
  assign G2660 = G2631 & G3553 & G389;
  assign G2666 = G2639 & G3553 & G400;
  assign G2672 = G2647 & G3553 & G411;
  assign G2678 = G2655 & G3553 & G374;
  assign G2684 = G3547 & G2627;
  assign G2689 = G3547 & G2635;
  assign G2694 = G3547 & G2643;
  assign G2699 = G3547 & G2651;
  assign G2728 = ~G2721;
  assign G2741 = ~G2734;
  assign G2748 = G292 & G2721;
  assign G2750 = G288 & G2721;
  assign G2752 = G280 & G2721;
  assign G2754 = G272 & G2721;
  assign G2756 = G264 & G2721;
  assign G2758 = G241 & G2734;
  assign G2760 = G233 & G2734;
  assign G2762 = G225 & G2734;
  assign G2764 = G217 & G2734;
  assign G2766 = G209 & G2734;
  assign G2827 = G1701;
  assign G2838 = ~G2828;
  assign G2847 = ~G2822;
  assign G2885 = ~G2882;
  assign G2889 = ~G2886;
  assign G2893 = ~G2890;
  assign G2897 = ~G2894;
  assign G2901 = ~G2898;
  assign G2905 = ~G2902;
  assign G2906 = G2393 & G2886;
  assign G2909 = G2894 & G2393 & G479;
  assign G2913 = G2902 & G2393 & G490;
  assign G2918 = G3554 & G2882;
  assign G2922 = G3554 & G2890;
  assign G2927 = G3554 & G2898;
  assign G2951 = ~G2948;
  assign G2955 = ~G2952;
  assign G2959 = ~G2956;
  assign G2963 = ~G2960;
  assign G2967 = ~G2964;
  assign G2971 = ~G2968;
  assign G2973 = G2952 & G3553 & G503;
  assign G2980 = ~G2979;
  assign G2982 = G2960 & G3553 & G523;
  assign G2988 = G2968 & G3553 & G534;
  assign G2994 = G3547 & G2948;
  assign G3001 = G3547 & G2956;
  assign G3006 = G3547 & G2964;
  assign G3027 = ~G3024;
  assign G3031 = ~G3028;
  assign G3035 = ~G3032;
  assign G3039 = ~G3036;
  assign G3043 = ~G3040;
  assign G3047 = ~G3044;
  assign G3051 = ~G3048;
  assign G3055 = ~G3052;
  assign G3056 = G3028 & G2393 & G389;
  assign G3060 = G3036 & G2393 & G400;
  assign G3064 = G3044 & G2393 & G411;
  assign G3068 = G3052 & G2393 & G374;
  assign G3073 = G3554 & G3024;
  assign G3078 = G3554 & G3032;
  assign G3083 = G3554 & G3040;
  assign G3088 = G3554 & G3048;
  assign G3099 = ~G3092;
  assign G3112 = ~G3105;
  assign G3119 = G372 & G3092;
  assign G3121 = G366 & G3092;
  assign G3123 = G358 & G3092;
  assign G3125 = G348 & G3092;
  assign G3126 = G338 & G3092;
  assign G3128 = G331 & G3105;
  assign G3130 = G323 & G3105;
  assign G3132 = G315 & G3105;
  assign G3134 = G307 & G3105;
  assign G3136 = G299 & G3105;
  assign G3187 = ~G3181;
  assign G3193 = G83 & G3181;
  assign G3196 = G86 & G3181;
  assign G3199 = G88 & G3181;
  assign G3202 = G88 & G3181;
  assign G3207 = ~G3204;
  assign G3211 = ~G3208;
  assign G3215 = ~G3212;
  assign G3219 = ~G3216;
  assign G3223 = ~G3220;
  assign G3227 = ~G3224;
  assign G3228 = G3208 & G2405 & G503;
  assign G3232 = G2405 & G514;
  assign G3234 = G3216 & G2405 & G523;
  assign G3238 = G3224 & G2405 & G534;
  assign G3243 = G3555 & G3204;
  assign G3247 = G3555 | G514;
  assign G3249 = G3555 & G3212;
  assign G3253 = G3555 & G3220;
  assign G3259 = ~G3256;
  assign G3263 = ~G3260;
  assign G3267 = ~G3264;
  assign G3271 = ~G3268;
  assign G3275 = ~G3272;
  assign G3279 = ~G3276;
  assign G3280 = G2405 & G3260;
  assign G3283 = G3268 & G2405 & G479;
  assign G3287 = G3276 & G2405 & G490;
  assign G3292 = G3555 & G3256;
  assign G3295 = G3555 & G3264;
  assign G3299 = G3555 & G3272;
  assign G3305 = ~G3302;
  assign G3306 = G2816;
  assign G3310 = G2816;
  assign G3317 = ~G3314;
  assign G3318 = G2816;
  assign G3322 = G2816;
  assign G3326 = G2405 & G3302;
  assign G3333 = G2405 & G3314;
  assign G3357 = ~G3354;
  assign G3361 = ~G3358;
  assign G3365 = ~G3362;
  assign G3369 = ~G3366;
  assign G3373 = ~G3370;
  assign G3377 = ~G3374;
  assign G3381 = ~G3378;
  assign G3385 = ~G3382;
  assign G3386 = G3358 & G2393 & G457;
  assign G3390 = G3366 & G2393 & G468;
  assign G3394 = G3374 & G2393 & G422;
  assign G3398 = G3382 & G2393 & G435;
  assign G3403 = G3554 & G3354;
  assign G3408 = G3554 & G3362;
  assign G3413 = G3554 & G3370;
  assign G3418 = G3554 & G3378;
  assign G5088 = ~G5082;
  assign G5089 = ~G5085;
  assign G5096 = ~G5090;
  assign G5097 = ~G5093;
  assign G3489 = G3440;
  assign G3493 = G3440;
  assign G3570 = ~G3558;
  assign G3594 = ~G3582;
  assign G3622 = ~G3616;
  assign G3632 = ~G3628;
  assign G3637 = G97 & G3616;
  assign G3640 = G94 & G3616;
  assign G3643 = G97 & G3616;
  assign G3646 = G94 & G3616;
  assign G3672 = ~G3660;
  assign G3696 = ~G3684;
  assign G3745 = ~G3737;
  assign G3765 = ~G3757;
  assign G3803 = ~G3795;
  assign G3823 = ~G3815;
  assign G5338 = ~G5332;
  assign G5339 = ~G5335;
  assign G5346 = ~G5340;
  assign G5347 = ~G5343;
  assign G5354 = ~G5348;
  assign G5355 = ~G5351;
  assign G3979 = ~G3972;
  assign G3998 = ~G3991;
  assign G4037 = ~G4030;
  assign G4056 = ~G4049;
  assign G4094 = G4110;
  assign G5104 = ~G5098;
  assign G5105 = ~G5101;
  assign G5114 = ~G5108;
  assign G5115 = ~G5111;
  assign G5362 = ~G5356;
  assign G5363 = ~G5359;
  assign G5366 = G2816;
  assign G5373 = ~G5369;
  assign G993 = G1688;
  assign G978 = G1688;
  assign G949 = G1688;
  assign G939 = G1688;
  assign G2568 = G2540 & G457 & G3551;
  assign G2574 = G2548 & G468 & G3551;
  assign G2580 = G2556 & G422 & G3551;
  assign G2586 = G2564 & G435 & G3551;
  assign G2592 = G3549 & G2536;
  assign G2597 = G3549 & G2544;
  assign G2602 = G3549 & G2552;
  assign G2607 = G3549 & G2560;
  assign G2662 = G2634 & G389 & G3551;
  assign G2668 = G2642 & G400 & G3551;
  assign G2674 = G2650 & G411 & G3551;
  assign G2680 = G2658 & G374 & G3551;
  assign G2686 = G3549 & G2630;
  assign G2691 = G3549 & G2638;
  assign G2696 = G3549 & G2646;
  assign G2701 = G3549 & G2654;
  assign G2907 = G2370 & G2889;
  assign G2910 = G2897 & G479 & G2370;
  assign G2914 = G2905 & G490 & G2370;
  assign G2920 = G3556 & G2885;
  assign G2924 = G3556 & G2893;
  assign G2929 = G3556 & G2901;
  assign G2975 = G2955 & G503 & G3551;
  assign G2984 = G2963 & G523 & G3551;
  assign G2990 = G2971 & G534 & G3551;
  assign G2996 = G3549 & G2951;
  assign G3003 = G3549 & G2959;
  assign G3008 = G3549 & G2967;
  assign G3015 = G2980 & G2999;
  assign G3057 = G3031 & G389 & G2370;
  assign G3061 = G3039 & G400 & G2370;
  assign G3065 = G3047 & G411 & G2370;
  assign G3069 = G3055 & G374 & G2370;
  assign G3075 = G3556 & G3027;
  assign G3080 = G3556 & G3035;
  assign G3085 = G3556 & G3043;
  assign G3090 = G3556 & G3051;
  assign G3229 = G3211 & G503 & G2382;
  assign G3233 = ~G3232;
  assign G3235 = G3219 & G523 & G2382;
  assign G3239 = G3227 & G534 & G2382;
  assign G3244 = G2361 & G3207;
  assign G3250 = G2361 & G3215;
  assign G3254 = G2361 & G3223;
  assign G3281 = G2382 & G3263;
  assign G3284 = G3271 & G479 & G2382;
  assign G3288 = G3279 & G490 & G2382;
  assign G3293 = G2361 & G3259;
  assign G3296 = G2361 & G3267;
  assign G3300 = G2361 & G3275;
  assign G3327 = G2382 & G3305;
  assign G3334 = G2382 & G3317;
  assign G3387 = G3361 & G457 & G2370;
  assign G3391 = G3369 & G468 & G2370;
  assign G3395 = G3377 & G422 & G2370;
  assign G3399 = G3385 & G435 & G2370;
  assign G3405 = G3556 & G3357;
  assign G3410 = G3556 & G3365;
  assign G3415 = G3556 & G3373;
  assign G3420 = G3556 & G3381;
  assign G3422 = ~G5085 | ~G5088;
  assign G3423 = ~G5082 | ~G5089;
  assign G3431 = ~G5093 | ~G5096;
  assign G3432 = ~G5090 | ~G5097;
  assign G3895 = ~G5335 | ~G5338;
  assign G3896 = ~G5332 | ~G5339;
  assign G3904 = ~G5343 | ~G5346;
  assign G3905 = ~G5340 | ~G5347;
  assign G3913 = ~G5351 | ~G5354;
  assign G3914 = ~G5348 | ~G5355;
  assign G889 = G4094;
  assign G5106 = ~G5101 | ~G5104;
  assign G5107 = ~G5098 | ~G5105;
  assign G5116 = ~G5111 | ~G5114;
  assign G5117 = ~G5108 | ~G5115;
  assign G5364 = ~G5359 | ~G5362;
  assign G5365 = ~G5356 | ~G5363;
  assign G593 = ~G4094;
  assign G2880 = G2838 & G2847;
  assign G2881 = G2828 & G2847;
  assign G1579 = G1552 & G200 & G1540;
  assign G1585 = G1552 & G203 & G1540;
  assign G1591 = G1552 & G197 & G1540;
  assign G1597 = G1552 & G194 & G1540;
  assign G1603 = G1552 & G191 & G1540;
  assign G1667 = G1633 & G182 & G1621;
  assign G1673 = G1633 & G188 & G1621;
  assign G1679 = G1633 & G155 & G1621;
  assign G1685 = G1633 & G149 & G1621;
  assign G2876 = G2838 & G2847;
  assign G2877 = G2828 & G2847;
  assign G2253 = G2226 & G200 & G2215;
  assign G2259 = G2226 & G203 & G2215;
  assign G2265 = G2226 & G197 & G2215;
  assign G2271 = G2226 & G194 & G2215;
  assign G2277 = G2226 & G191 & G2215;
  assign G2338 = G2304 & G182 & G2293;
  assign G2344 = G2304 & G188 & G2293;
  assign G2350 = G2304 & G155 & G2293;
  assign G2356 = G2304 & G149 & G2293;
  assign G2868 = G2838 & G2847;
  assign G2869 = G2828 & G2847;
  assign G710 = G3684 & G109 & G3672;
  assign G2872 = G2838 & G2847;
  assign G2873 = G2828 & G2847;
  assign G720 = G2442 & G11 & G2430;
  assign G725 = G3582 & G109 & G3570;
  assign G730 = G3582 & G46 & G3570;
  assign G735 = G3582 & G100 & G3570;
  assign G740 = G3582 & G91 & G3570;
  assign G745 = G3582 & G43 & G3570;
  assign G750 = G2442 & G76 & G2430;
  assign G755 = G2442 & G73 & G2430;
  assign G760 = G2442 & G67 & G2430;
  assign G765 = G2442 & G14 & G2430;
  assign G770 = G3684 & G46 & G3672;
  assign G775 = G3684 & G100 & G3672;
  assign G780 = G3684 & G91 & G3672;
  assign G785 = G3684 & G43 & G3672;
  assign G790 = G2500 & G76 & G2488;
  assign G795 = G2500 & G73 & G2488;
  assign G800 = G2500 & G67 & G2488;
  assign G805 = G2500 & G14 & G2488;
  assign G841 = G3815 & G120 & G3803;
  assign G857 = G2500 & G11 & G2488;
  assign G880 = G3757 & G118 & G3745;
  assign G1660 = G1633 & G176 & G1621;
  assign G2331 = G2304 & G176 & G2293;
  assign G2569 = G2566 | G2568;
  assign G2575 = G2572 | G2574;
  assign G2581 = G2578 | G2580;
  assign G2587 = G2584 | G2586;
  assign G2593 = G457 | G2590 | G2592;
  assign G2598 = G468 | G2595 | G2597;
  assign G2603 = G422 | G2600 | G2602;
  assign G2608 = G435 | G2605 | G2607;
  assign G2663 = G2660 | G2662;
  assign G2669 = G2666 | G2668;
  assign G2675 = G2672 | G2674;
  assign G2681 = G2678 | G2680;
  assign G2687 = G389 | G2684 | G2686;
  assign G2692 = G400 | G2689 | G2691;
  assign G2697 = G411 | G2694 | G2696;
  assign G2702 = G374 | G2699 | G2701;
  assign G2747 = G289 & G2728;
  assign G2749 = G281 & G2728;
  assign G2751 = G273 & G2728;
  assign G2753 = G265 & G2728;
  assign G2755 = G257 & G2728;
  assign G2757 = G234 & G2741;
  assign G2759 = G226 & G2741;
  assign G2761 = G218 & G2741;
  assign G2763 = G210 & G2741;
  assign G2765 = G206 & G2741;
  assign G2857 = ~G2847;
  assign G2908 = G2906 | G2907;
  assign G2911 = G2909 | G2910;
  assign G2915 = G2913 | G2914;
  assign G2925 = G479 | G2922 | G2924;
  assign G2930 = G490 | G2927 | G2929;
  assign G2933 = G2918 | G2920;
  assign G2976 = G2973 | G2975;
  assign G2985 = G2982 | G2984;
  assign G2991 = G2988 | G2990;
  assign G2997 = G503 | G2994 | G2996;
  assign G3004 = G523 | G3001 | G3003;
  assign G3009 = G534 | G3006 | G3008;
  assign G3058 = G3056 | G3057;
  assign G3062 = G3060 | G3061;
  assign G3066 = G3064 | G3065;
  assign G3070 = G3068 | G3069;
  assign G3076 = G389 | G3073 | G3075;
  assign G3081 = G400 | G3078 | G3080;
  assign G3086 = G411 | G3083 | G3085;
  assign G3091 = G374 | G3088 | G3090;
  assign G3118 = G369 & G3099;
  assign G3120 = G361 & G3099;
  assign G3122 = G351 & G3099;
  assign G3124 = G341 & G3099;
  assign G3127 = G324 & G3112;
  assign G3129 = G316 & G3112;
  assign G3131 = G308 & G3112;
  assign G3133 = G302 & G3112;
  assign G3135 = G293 & G3112;
  assign G3147 = G3099 | G3126;
  assign G3192 = G83 & G3187;
  assign G3195 = G87 & G3187;
  assign G3198 = G34 & G3187;
  assign G3201 = G34 & G3187;
  assign G3230 = G3228 | G3229;
  assign G3236 = G3234 | G3235;
  assign G3240 = G3238 | G3239;
  assign G3245 = G503 | G3243 | G3244;
  assign G3251 = G523 | G3249 | G3250;
  assign G3255 = G534 | G3253 | G3254;
  assign G3282 = G3280 | G3281;
  assign G3285 = G3283 | G3284;
  assign G3289 = G3287 | G3288;
  assign G3297 = G479 | G3295 | G3296;
  assign G3301 = G490 | G3299 | G3300;
  assign G3309 = ~G3306;
  assign G3313 = ~G3310;
  assign G3321 = ~G3318;
  assign G3325 = ~G3322;
  assign G3328 = G3326 | G3327;
  assign G3329 = G3310 & G2405 & G446;
  assign G3335 = G3333 | G3334;
  assign G3336 = G3322 & G2405 & G446;
  assign G3341 = G3555 & G3306;
  assign G3345 = G3555 & G3318;
  assign G3388 = G3386 | G3387;
  assign G3392 = G3390 | G3391;
  assign G3396 = G3394 | G3395;
  assign G3400 = G3398 | G3399;
  assign G3406 = G457 | G3403 | G3405;
  assign G3411 = G468 | G3408 | G3410;
  assign G3416 = G422 | G3413 | G3415;
  assign G3421 = G435 | G3418 | G3420;
  assign G3424 = ~G3422 | ~G3423;
  assign G3433 = ~G3431 | ~G3432;
  assign G3492 = ~G3489;
  assign G3496 = ~G3493;
  assign G3780 = G3757 & G117 & G3745;
  assign G3783 = G3757 & G126 & G3745;
  assign G3786 = G3757 & G127 & G3745;
  assign G3789 = G3757 & G128 & G3745;
  assign G3838 = G3815 & G131 & G3803;
  assign G3841 = G3815 & G129 & G3803;
  assign G3844 = G3815 & G119 & G3803;
  assign G3847 = G3815 & G130 & G3803;
  assign G3897 = ~G3895 | ~G3896;
  assign G3906 = ~G3904 | ~G3905;
  assign G3915 = ~G3913 | ~G3914;
  assign G4011 = G3991 & G122 & G3979;
  assign G4014 = G3991 & G113 & G3979;
  assign G4017 = G3991 & G53 & G3979;
  assign G4020 = G3991 & G114 & G3979;
  assign G4023 = G3991 & G115 & G3979;
  assign G4069 = G4049 & G52 & G4037;
  assign G4072 = G4049 & G112 & G4037;
  assign G4075 = G4049 & G116 & G4037;
  assign G4078 = G4049 & G121 & G4037;
  assign G4081 = G4049 & G123 & G4037;
  assign G5206 = ~G5116 | ~G5117;
  assign G5209 = ~G5106 | ~G5107;
  assign G5307 = G3233 & G3247;
  assign G5322 = G3292 | G3293;
  assign G5372 = ~G5366;
  assign G5375 = ~G5366 | ~G5373;
  assign G5399 = ~G5364 | ~G5365;
  assign G2813 = ~G3015;
  assign G3197 = G3195 | G3196;
  assign G3200 = G3198 | G3199;
  assign G3203 = G3201 | G3202;
  assign G3194 = G3192 | G3193;
  assign G2570 = ~G2569;
  assign G2576 = ~G2575;
  assign G2582 = ~G2581;
  assign G2588 = ~G2587;
  assign G2664 = ~G2663;
  assign G2670 = ~G2669;
  assign G2676 = ~G2675;
  assign G2682 = ~G2681;
  assign G2767 = G2749 | G2750;
  assign G2772 = G2751 | G2752;
  assign G2776 = G2753 | G2754;
  assign G2780 = G2755 | G2756;
  assign G2784 = G2757 | G2758;
  assign G2788 = G2759 | G2760;
  assign G2794 = G2761 | G2762;
  assign G2798 = G2763 | G2764;
  assign G2802 = G2765 | G2766;
  assign G2912 = ~G2911;
  assign G2916 = ~G2915;
  assign G2936 = ~G2908;
  assign G2977 = ~G2976;
  assign G2986 = ~G2985;
  assign G2992 = ~G2991;
  assign G3059 = ~G3058;
  assign G3063 = ~G3062;
  assign G3067 = ~G3066;
  assign G3071 = ~G3070;
  assign G3137 = G3120 | G3121;
  assign G3139 = G3122 | G3123;
  assign G3143 = G3124 | G3125;
  assign G3151 = G3127 | G3128;
  assign G3155 = G3129 | G3130;
  assign G3161 = G3131 | G3132;
  assign G3165 = G3133 | G3134;
  assign G3167 = G3135 | G3136;
  assign G3231 = ~G3230;
  assign G3237 = ~G3236;
  assign G3241 = ~G3240;
  assign G3286 = ~G3285;
  assign G3290 = ~G3289;
  assign G3330 = G3313 & G446 & G2382;
  assign G3337 = G3325 & G446 & G2382;
  assign G3342 = G2361 & G3309;
  assign G3346 = G2361 & G3321;
  assign G3348 = ~G3328;
  assign G3352 = ~G3335;
  assign G3389 = ~G3388;
  assign G3393 = ~G3392;
  assign G3397 = ~G3396;
  assign G3401 = ~G3400;
  assign G3845 = G3823 & G3015 & G3803;
  assign G5126 = G3118 | G3119;
  assign G5178 = G2747 | G2748;
  assign G5325 = ~G3282;
  assign G5374 = ~G5369 | ~G5372;
  assign G2810 = ~G2933;
  assign G635 = G3197 & G3176;
  assign G2878 = G2857 & G24 & G2838;
  assign G2879 = G2857 & G25 & G2828;
  assign G2874 = G2857 & G26 & G2838;
  assign G2875 = G2857 & G81 & G2828;
  assign G703 = G3200 & G3176;
  assign G2866 = G2857 & G79 & G2838;
  assign G2867 = G2857 & G23 & G2828;
  assign G2870 = G2857 & G82 & G2838;
  assign G2871 = G2857 & G80 & G2828;
  assign G716 = G3203 & G3176;
  assign G819 = G3194 & G3176;
  assign G1789 = G3147 & G514;
  assign G2036 = G514 & G3147;
  assign G2611 = G2570 & G2593;
  assign G2615 = G2576 & G2598;
  assign G2619 = G2582 & G2603;
  assign G2623 = G2588 & G2608;
  assign G2705 = G2664 & G2687;
  assign G2709 = G2670 & G2692;
  assign G2713 = G2676 & G2697;
  assign G2717 = G2682 & G2702;
  assign G2939 = G2912 & G2925;
  assign G2942 = G2916 & G2930;
  assign G2945 = G2933;
  assign G3012 = G2977 & G2997;
  assign G3018 = G2986 & G3004;
  assign G3021 = G2992 & G3009;
  assign G3331 = G3329 | G3330;
  assign G3338 = G3336 | G3337;
  assign G3343 = G446 | G3341 | G3342;
  assign G3347 = G446 | G3345 | G3346;
  assign G3428 = ~G3424;
  assign G3437 = ~G3433;
  assign G3514 = G3489 & G3433 & G3424;
  assign G3836 = G3823 & G3352 & G3803;
  assign G3852 = G3071 & G3091;
  assign G5311 = ~G5307;
  assign G3901 = ~G3897;
  assign G3910 = ~G3906;
  assign G3934 = G3915;
  assign G3938 = G3915;
  assign G4652 = G3147;
  assign G4783 = G3147;
  assign G5137 = G3147;
  assign G5212 = ~G5206;
  assign G5213 = ~G5209;
  assign G5260 = G3063 & G3081;
  assign G5263 = G3067 & G3086;
  assign G5268 = G3401 & G3421;
  assign G5271 = G3059 & G3076;
  assign G5276 = G3393 & G3411;
  assign G5279 = G3397 & G3416;
  assign G5289 = G3389 & G3406;
  assign G5296 = G3237 & G3251;
  assign G5299 = G3241 & G3255;
  assign G5304 = G3231 & G3245;
  assign G5312 = G3286 & G3297;
  assign G5315 = G3290 & G3301;
  assign G5328 = ~G5322;
  assign G5396 = ~G5374 | ~G5375;
  assign G5403 = ~G5399;
  assign G1286 = G446 & G2802;
  assign G2809 = ~G2936;
  assign G597 = ~G3348;
  assign G1031 = G2802 & G446;
  assign G636 = ~G635;
  assign G637 = G2881 | G2880 | G2878 | G2879;
  assign G671 = G2877 | G2876 | G2874 | G2875;
  assign G704 = ~G703;
  assign G705 = G2869 | G2868 | G2866 | G2867;
  assign G713 = G2873 | G2872 | G2870 | G2871;
  assign G717 = ~G716;
  assign G820 = ~G819;
  assign G1046 = G2798 & G457;
  assign G1064 = G2794 & G468;
  assign G1071 = G422 & G2788;
  assign G1097 = G2784 & G435;
  assign G1111 = G2780 & G389;
  assign G1128 = G2776 & G400;
  assign G1145 = G2772 & G411;
  assign G1160 = G2767 & G374;
  assign G1301 = G457 & G2798;
  assign G1318 = G468 & G2794;
  assign G1324 = G422 & G2788;
  assign G1341 = G435 & G2784;
  assign G1359 = G389 & G2780;
  assign G1382 = G400 & G2776;
  assign G1404 = G411 & G2772;
  assign G1412 = G374 & G2767;
  assign G1704 = ~G3167;
  assign G1712 = ~G3165;
  assign G1724 = G3165;
  assign G1742 = G3161 & G479;
  assign G1749 = G490 & G3155;
  assign G1775 = G3151 & G503;
  assign G1806 = G3143 & G523;
  assign G1823 = G3139 & G534;
  assign G1829 = ~G3137;
  assign G1837 = G3137;
  assign G1958 = ~G3167;
  assign G1966 = ~G3165;
  assign G1978 = G3165;
  assign G1995 = G479 & G3161;
  assign G2001 = G490 & G3155;
  assign G2018 = G503 & G3151;
  assign G2059 = G523 & G3143;
  assign G2081 = G534 & G3139;
  assign G2089 = G3137;
  assign G2106 = ~G3137;
  assign G3170 = G3167;
  assign G3332 = ~G3331;
  assign G3339 = ~G3338;
  assign G5132 = ~G5126;
  assign G5184 = ~G5178;
  assign G3853 = ~G3852;
  assign G3874 = ~G3348;
  assign G4076 = G4056 & G2936 & G4037;
  assign G4116 = G2802;
  assign G4124 = G2798;
  assign G4132 = G2794;
  assign G4140 = G2788;
  assign G4148 = G2784;
  assign G4156 = G2780;
  assign G4164 = G2776;
  assign G4172 = G2772;
  assign G4180 = G2767;
  assign G4228 = ~G422 & ~G2788;
  assign G4279 = G2802;
  assign G4287 = G2798;
  assign G4295 = G2794;
  assign G4303 = G2784;
  assign G4311 = G2780;
  assign G4319 = G2776;
  assign G4327 = G2772;
  assign G4335 = G2788;
  assign G4343 = G2767;
  assign G4348 = ~G422 & ~G2788;
  assign G4464 = ~G374 & ~G2767;
  assign G4628 = G3161;
  assign G4636 = G3155;
  assign G4644 = G3151;
  assign G4660 = G3143;
  assign G4668 = G3139;
  assign G4716 = ~G490 & ~G3155;
  assign G4767 = G3161;
  assign G4775 = G3151;
  assign G4791 = G3143;
  assign G4799 = G3139;
  assign G4807 = G3155;
  assign G4812 = ~G490 & ~G3155;
  assign G5118 = G3139;
  assign G5121 = G3143;
  assign G5129 = G3137;
  assign G5134 = G3151;
  assign G5142 = G3161;
  assign G5145 = G3155;
  assign G5152 = G3167;
  assign G5155 = G3165;
  assign G5162 = G2788;
  assign G5165 = G2784;
  assign G5170 = G2798;
  assign G5173 = G2794;
  assign G5181 = G2802;
  assign G5186 = G2772;
  assign G5189 = G2767;
  assign G5196 = G2780;
  assign G5199 = G2776;
  assign G5214 = ~G5209 | ~G5212;
  assign G5215 = ~G5206 | ~G5213;
  assign G5329 = ~G5325;
  assign G5330 = ~G5325 | ~G5328;
  assign G2807 = ~G2942;
  assign G2808 = ~G2939;
  assign G2811 = ~G3021;
  assign G2812 = ~G3018;
  assign G2814 = ~G3012;
  assign G2626 = ~G2623;
  assign G2622 = ~G2619;
  assign G2618 = ~G2615;
  assign G2614 = ~G2611;
  assign G2720 = ~G2717;
  assign G2716 = ~G2713;
  assign G2712 = ~G2709;
  assign G2708 = ~G2705;
  assign G639 = G637 & G2827;
  assign G673 = G671 & G2827;
  assign G707 = G705 & G2827;
  assign G715 = G713 & G2827;
  assign G3731 = G3721 & G2945 & G3728;
  assign G4658 = ~G4652;
  assign G1777 = ~G4652 | ~G4659;
  assign G2019 = ~G4783 | ~G4786;
  assign G4787 = ~G4783;
  assign G3350 = G3332 & G3343;
  assign G3353 = G3339 & G3347;
  assign G5141 = ~G5137;
  assign G3513 = G3492 & G3428 & G3433;
  assign G3516 = G3496 & G3424 & G3437;
  assign G3517 = G3493 & G3437 & G3428;
  assign G3778 = G3765 & G2717 & G3745;
  assign G3781 = G3765 & G2713 & G3745;
  assign G3784 = G3765 & G2709 & G3745;
  assign G3787 = G3765 & G2705 & G3745;
  assign G3839 = G3823 & G3021 & G3803;
  assign G3842 = G3823 & G3018 & G3803;
  assign G5266 = ~G5260;
  assign G5267 = ~G5263;
  assign G5274 = ~G5268;
  assign G5275 = ~G5271;
  assign G5302 = ~G5296;
  assign G5303 = ~G5299;
  assign G5310 = ~G5304;
  assign G3891 = ~G5304 | ~G5311;
  assign G3937 = ~G3934;
  assign G3941 = ~G3938;
  assign G3955 = G3934 & G3906 & G3897;
  assign G3958 = G3938 & G3910 & G3901;
  assign G4009 = G3998 & G2623 & G3979;
  assign G4012 = G3998 & G2619 & G3979;
  assign G4015 = G3998 & G2615 & G3979;
  assign G4018 = G3998 & G2611 & G3979;
  assign G4067 = G4056 & G3012 & G4037;
  assign G4070 = G4056 & G2942 & G4037;
  assign G4073 = G4056 & G2939 & G4037;
  assign G4079 = G4056 & G2945 & G4037;
  assign G5239 = ~G5214 | ~G5215;
  assign G5282 = ~G5276;
  assign G5283 = ~G5279;
  assign G5293 = ~G5289;
  assign G5318 = ~G5312;
  assign G5319 = ~G5315;
  assign G5331 = ~G5322 | ~G5329;
  assign G5402 = ~G5396;
  assign G5405 = ~G5396 | ~G5403;
  assign G595 = G2810 & G2809 & G2807 & G2808;
  assign G596 = G2814 & G2813 & G2811 & G2812;
  assign G607 = G2614 & G2618 & G2626 & G2622;
  assign G608 = G2708 & G2712 & G2720 & G2716;
  assign G1845 = G1704 & G1724;
  assign G1846 = G1742 & G1712 & G1704;
  assign G2115 = G1958 & G1978;
  assign G2116 = G1995 & G1966 & G1958;
  assign G4122 = ~G4116;
  assign G1022 = ~G4116 | ~G4123;
  assign G4130 = ~G4124;
  assign G1033 = ~G4124 | ~G4131;
  assign G4138 = ~G4132;
  assign G1051 = ~G4132 | ~G4139;
  assign G4146 = ~G4140;
  assign G1079 = ~G4140 | ~G4147;
  assign G4154 = ~G4148;
  assign G1088 = ~G4148 | ~G4155;
  assign G4162 = ~G4156;
  assign G1099 = ~G4156 | ~G4163;
  assign G4170 = ~G4164;
  assign G1115 = ~G4164 | ~G4171;
  assign G4178 = ~G4172;
  assign G1133 = ~G4172 | ~G4179;
  assign G4186 = ~G4180;
  assign G1151 = ~G4180 | ~G4187;
  assign G4234 = ~G4228;
  assign G1276 = ~G4279 | ~G4282;
  assign G4283 = ~G4279;
  assign G1287 = ~G4287 | ~G4290;
  assign G4291 = ~G4287;
  assign G1305 = ~G4295 | ~G4298;
  assign G4299 = ~G4295;
  assign G1330 = ~G4303 | ~G4306;
  assign G4307 = ~G4303;
  assign G1342 = ~G4311 | ~G4314;
  assign G4315 = ~G4311;
  assign G1363 = ~G4319 | ~G4322;
  assign G4323 = ~G4319;
  assign G1388 = ~G4327 | ~G4330;
  assign G4331 = ~G4327;
  assign G1420 = ~G4335 | ~G4338;
  assign G4339 = ~G4335;
  assign G1428 = ~G4343 | ~G4346;
  assign G4347 = ~G4343;
  assign G4634 = ~G4628;
  assign G1729 = ~G4628 | ~G4635;
  assign G4642 = ~G4636;
  assign G1757 = ~G4636 | ~G4643;
  assign G4650 = ~G4644;
  assign G1766 = ~G4644 | ~G4651;
  assign G1776 = ~G4655 | ~G4658;
  assign G4666 = ~G4660;
  assign G1793 = ~G4660 | ~G4667;
  assign G4674 = ~G4668;
  assign G1811 = ~G4668 | ~G4675;
  assign G1849 = G1712 & G1742;
  assign G1852 = G1712 & G1742;
  assign G1875 = G54 & G1829;
  assign G4722 = ~G4716;
  assign G1982 = ~G4767 | ~G4770;
  assign G4771 = ~G4767;
  assign G2007 = ~G4775 | ~G4778;
  assign G4779 = ~G4775;
  assign G2020 = ~G4780 | ~G4787;
  assign G2040 = ~G4791 | ~G4794;
  assign G4795 = ~G4791;
  assign G2065 = ~G4799 | ~G4802;
  assign G4803 = ~G4799;
  assign G2097 = ~G4807 | ~G4810;
  assign G4811 = ~G4807;
  assign G2119 = G1966 & G1995;
  assign G2122 = G1966 & G1995;
  assign G5124 = ~G5118;
  assign G5125 = ~G5121;
  assign G3452 = ~G5129 | ~G5132;
  assign G5133 = ~G5129;
  assign G5140 = ~G5134;
  assign G3462 = ~G5134 | ~G5141;
  assign G5168 = ~G5162;
  assign G5169 = ~G5165;
  assign G5176 = ~G5170;
  assign G5177 = ~G5173;
  assign G3484 = ~G5181 | ~G5184;
  assign G5185 = ~G5181;
  assign G3515 = ~G3513 & ~G3514;
  assign G3518 = ~G3516 & ~G3517;
  assign G3857 = ~G3853;
  assign G3860 = ~G5263 | ~G5266;
  assign G3861 = ~G5260 | ~G5267;
  assign G3869 = ~G5271 | ~G5274;
  assign G3870 = ~G5268 | ~G5275;
  assign G3878 = ~G3874;
  assign G3881 = ~G5299 | ~G5302;
  assign G3882 = ~G5296 | ~G5303;
  assign G3890 = ~G5307 | ~G5310;
  assign G3954 = G3937 & G3901 & G3906;
  assign G3957 = G3941 & G3897 & G3910;
  assign G4021 = G3998 & G3353 & G3979;
  assign G4099 = ~G3170;
  assign G4236 = G1071;
  assign G4354 = ~G4348;
  assign G4406 = G1324;
  assign G4470 = ~G4464;
  assign G4552 = G1412;
  assign G4679 = G1829;
  assign G4687 = G1704;
  assign G4695 = G1704;
  assign G4703 = G1712;
  assign G4711 = G1712;
  assign G4724 = G1749;
  assign G4818 = ~G4812;
  assign G4855 = G1958;
  assign G4865 = G1966;
  assign G4870 = G2001;
  assign G4913 = G1958;
  assign G4923 = G1966;
  assign G4951 = G2106;
  assign G5006 = G2089;
  assign G5039 = G2106;
  assign G5148 = ~G5142;
  assign G5149 = ~G5145;
  assign G5158 = ~G5152;
  assign G5159 = ~G5155;
  assign G5192 = ~G5186;
  assign G5193 = ~G5189;
  assign G5202 = ~G5196;
  assign G5203 = ~G5199;
  assign G5284 = ~G5279 | ~G5282;
  assign G5285 = ~G5276 | ~G5283;
  assign G5320 = ~G5315 | ~G5318;
  assign G5321 = ~G5312 | ~G5319;
  assign G5386 = ~G5330 | ~G5331;
  assign G5404 = ~G5399 | ~G5402;
  assign G598 = G597 & G595 & G596;
  assign G609 = ~G3350;
  assign G1021 = ~G4119 | ~G4122;
  assign G1032 = ~G4127 | ~G4130;
  assign G1050 = ~G4135 | ~G4138;
  assign G1078 = ~G4143 | ~G4146;
  assign G1087 = ~G4151 | ~G4154;
  assign G1098 = ~G4159 | ~G4162;
  assign G1114 = ~G4167 | ~G4170;
  assign G1132 = ~G4175 | ~G4178;
  assign G1150 = ~G4183 | ~G4186;
  assign G1277 = ~G4276 | ~G4283;
  assign G1288 = ~G4284 | ~G4291;
  assign G1306 = ~G4292 | ~G4299;
  assign G1331 = ~G4300 | ~G4307;
  assign G1343 = ~G4308 | ~G4315;
  assign G1364 = ~G4316 | ~G4323;
  assign G1389 = ~G4324 | ~G4331;
  assign G1421 = ~G4332 | ~G4339;
  assign G1429 = ~G4340 | ~G4347;
  assign G1728 = ~G4631 | ~G4634;
  assign G1756 = ~G4639 | ~G4642;
  assign G1765 = ~G4647 | ~G4650;
  assign G1778 = ~G1776 | ~G1777;
  assign G1792 = ~G4663 | ~G4666;
  assign G1810 = ~G4671 | ~G4674;
  assign G1983 = ~G4764 | ~G4771;
  assign G2008 = ~G4772 | ~G4779;
  assign G2021 = ~G2019 | ~G2020;
  assign G2041 = ~G4788 | ~G4795;
  assign G2066 = ~G4796 | ~G4803;
  assign G2098 = ~G4804 | ~G4811;
  assign G3443 = ~G5121 | ~G5124;
  assign G3444 = ~G5118 | ~G5125;
  assign G3453 = ~G5126 | ~G5133;
  assign G3461 = ~G5137 | ~G5140;
  assign G3466 = ~G5165 | ~G5168;
  assign G3467 = ~G5162 | ~G5169;
  assign G3475 = ~G5173 | ~G5176;
  assign G3476 = ~G5170 | ~G5177;
  assign G3485 = ~G5178 | ~G5185;
  assign G5243 = ~G5239;
  assign G3862 = ~G3860 | ~G3861;
  assign G3871 = ~G3869 | ~G3870;
  assign G3883 = ~G3881 | ~G3882;
  assign G3892 = ~G3890 | ~G3891;
  assign G3956 = ~G3954 & ~G3955;
  assign G3959 = ~G3957 & ~G3958;
  assign G4756 = G1837 | G1875;
  assign G5150 = ~G5145 | ~G5148;
  assign G5151 = ~G5142 | ~G5149;
  assign G5160 = ~G5155 | ~G5158;
  assign G5161 = ~G5152 | ~G5159;
  assign G5194 = ~G5189 | ~G5192;
  assign G5195 = ~G5186 | ~G5193;
  assign G5204 = ~G5199 | ~G5202;
  assign G5205 = ~G5196 | ~G5203;
  assign G5236 = ~G3518 | ~G3515;
  assign G5286 = G3350;
  assign G5379 = ~G5284 | ~G5285;
  assign G5389 = ~G5320 | ~G5321;
  assign G5425 = ~G5404 | ~G5405;
  assign G610 = G609 & G607 & G608;
  assign G1023 = ~G1021 | ~G1022;
  assign G1034 = ~G1032 | ~G1033;
  assign G1052 = ~G1050 | ~G1051;
  assign G1080 = ~G1078 | ~G1079;
  assign G1089 = ~G1087 | ~G1088;
  assign G1100 = ~G1098 | ~G1099;
  assign G1116 = ~G1114 | ~G1115;
  assign G1134 = ~G1132 | ~G1133;
  assign G1152 = ~G1150 | ~G1151;
  assign G4242 = ~G4236;
  assign G1278 = ~G1276 | ~G1277;
  assign G1289 = ~G1287 | ~G1288;
  assign G1307 = ~G1305 | ~G1306;
  assign G1332 = ~G1330 | ~G1331;
  assign G1344 = ~G1342 | ~G1343;
  assign G1365 = ~G1363 | ~G1364;
  assign G1390 = ~G1388 | ~G1389;
  assign G1422 = ~G1420 | ~G1421;
  assign G1430 = ~G1428 | ~G1429;
  assign G1730 = ~G1728 | ~G1729;
  assign G1758 = ~G1756 | ~G1757;
  assign G1767 = ~G1765 | ~G1766;
  assign G1794 = ~G1792 | ~G1793;
  assign G1812 = ~G1810 | ~G1811;
  assign G1876 = ~G4679 | ~G4682;
  assign G4683 = ~G4679;
  assign G4691 = ~G4687;
  assign G4699 = ~G4695;
  assign G4707 = ~G4703;
  assign G4715 = ~G4711;
  assign G4730 = ~G4724;
  assign G1984 = ~G1982 | ~G1983;
  assign G2009 = ~G2007 | ~G2008;
  assign G2042 = ~G2040 | ~G2041;
  assign G2067 = ~G2065 | ~G2066;
  assign G2099 = ~G2097 | ~G2098;
  assign G4869 = ~G4865;
  assign G4927 = ~G4923;
  assign G3445 = ~G3443 | ~G3444;
  assign G3454 = ~G3452 | ~G3453;
  assign G3463 = ~G3461 | ~G3462;
  assign G3468 = ~G3466 | ~G3467;
  assign G3477 = ~G3475 | ~G3476;
  assign G3486 = ~G3484 | ~G3485;
  assign G4103 = G4099 & G3170;
  assign G4412 = ~G4406;
  assign G4558 = ~G4552;
  assign G4859 = ~G4855;
  assign G4876 = ~G4870;
  assign G4917 = ~G4913;
  assign G4955 = ~G4951;
  assign G5012 = ~G5006;
  assign G5043 = ~G5039;
  assign G5216 = ~G5160 | ~G5161;
  assign G5219 = ~G5150 | ~G5151;
  assign G5226 = ~G5204 | ~G5205;
  assign G5229 = ~G5194 | ~G5195;
  assign G5392 = ~G5386;
  assign G5422 = ~G3959 | ~G3956;
  assign G1866 = G1778 & G1806;
  assign G1877 = ~G4676 | ~G4683;
  assign G4762 = ~G4756;
  assign G2142 = G2021 & G2059;
  assign G2146 = G2021 & G2059;
  assign G5242 = ~G5236;
  assign G3532 = ~G5236 | ~G5243;
  assign G3866 = ~G3862;
  assign G3887 = ~G3883;
  assign G3918 = G3871;
  assign G3922 = G3871;
  assign G3926 = G3892;
  assign G3930 = G3892;
  assign G5429 = ~G5425;
  assign G4104 = G4099 | G4103;
  assign G4743 = G1778;
  assign G4991 = G2021;
  assign G5001 = G2021;
  assign G5292 = ~G5286;
  assign G5295 = ~G5286 | ~G5293;
  assign G5383 = ~G5379;
  assign G5393 = ~G5389;
  assign G5394 = ~G5389 | ~G5392;
  assign G1439 = G1278 & G1301;
  assign G1440 = G1318 & G1289 & G1278;
  assign G1441 = G1289 & G1324 & G1307 & G1278;
  assign G1847 = G1712 & G1749 & G1730 & G1704;
  assign G1168 = G1023 & G1046;
  assign G1169 = G1064 & G1034 & G1023;
  assign G1170 = G1034 & G1071 & G1052 & G1023;
  assign G2117 = G1966 & G2001 & G1984 & G1958;
  assign G1086 = ~G1080;
  assign G1166 = G1023 & G1052 & G1034 & G1080;
  assign G1171 = G1034 & G1064;
  assign G1172 = G1034 & G1052 & G1071;
  assign G1173 = G1034 & G1080 & G1052;
  assign G1174 = G1034 & G1064;
  assign G1175 = G1034 & G1071 & G1052;
  assign G1176 = G1052 & G1071;
  assign G1177 = G1080 & G1052;
  assign G1178 = G1052 & G1071;
  assign G1179 = G1134 & G1089 & G1116 & G1100 & G1152;
  assign G1181 = G1089 & G1111;
  assign G1182 = G1128 & G1100 & G1089;
  assign G1183 = G1100 & G1145 & G1116 & G1089;
  assign G1184 = G1100 & G1160 & G1089 & G1134 & G1116;
  assign G1188 = G1100 & G1128;
  assign G1189 = G1100 & G1116 & G1145;
  assign G1190 = G1100 & G1160 & G1134 & G1116;
  assign G1191 = G1100 & G1134 & G1116 & G4 & G1152;
  assign G1192 = G1145 & G1116;
  assign G1193 = G1160 & G1134 & G1116;
  assign G1194 = G1134 & G1116 & G4 & G1152;
  assign G1195 = G1134 & G1160;
  assign G1196 = G1134 & G4 & G1152;
  assign G1197 = G4 & G1152;
  assign G1437 = G1278 & G1289 & G1422 & G1307;
  assign G1442 = G1289 & G1318;
  assign G1443 = G1289 & G1307 & G1324;
  assign G1444 = G1289 & G1422 & G1307;
  assign G1445 = G1289 & G1318;
  assign G1446 = G1289 & G1307 & G1324;
  assign G1447 = G1307 & G1324;
  assign G1451 = G1332 & G1344 & G1365 & G1430 & G1390;
  assign G1454 = G1332 & G1359;
  assign G1455 = G1382 & G1344 & G1332;
  assign G1456 = G1344 & G1404 & G1365 & G1332;
  assign G1457 = G1344 & G1412 & G1332 & G1390 & G1365;
  assign G1465 = G1344 & G1382;
  assign G1466 = G1344 & G1365 & G1404;
  assign G1467 = G1344 & G1412 & G1390 & G1365;
  assign G1468 = G1390 & G1344 & G1430 & G1365;
  assign G1469 = G1344 & G1382;
  assign G1470 = G1344 & G1365 & G1404;
  assign G1471 = G1344 & G1412 & G1390 & G1365;
  assign G1472 = G1365 & G1404;
  assign G1473 = G1412 & G1390 & G1365;
  assign G1474 = G1390 & G1430 & G1365;
  assign G1475 = G1365 & G1404;
  assign G1476 = G1412 & G1390 & G1365;
  assign G1477 = G1390 & G1412;
  assign G1481 = G1422 & G1307;
  assign G1482 = G1430 & G1390;
  assign G1764 = ~G1758;
  assign G1843 = G1704 & G1730 & G1712 & G1758;
  assign G1850 = G1712 & G1730 & G1749;
  assign G1851 = G1712 & G1758 & G1730;
  assign G1853 = G1712 & G1749 & G1730;
  assign G1854 = G1730 & G1749;
  assign G1855 = G1758 & G1730;
  assign G1856 = G1730 & G1749;
  assign G1857 = G1812 & G1767 & G1794 & G1778 & G1829;
  assign G1859 = G1767 & G1789;
  assign G1860 = G1806 & G1778 & G1767;
  assign G1861 = G1778 & G1823 & G1794 & G1767;
  assign G1862 = G1778 & G1837 & G1767 & G1812 & G1794;
  assign G1867 = G1778 & G1794 & G1823;
  assign G1868 = G1778 & G1837 & G1812 & G1794;
  assign G1869 = G1778 & G1812 & G1794 & G54 & G1829;
  assign G1870 = G1823 & G1794;
  assign G1871 = G1837 & G1812 & G1794;
  assign G1872 = G1812 & G1794 & G54 & G1829;
  assign G1873 = G1812 & G1837;
  assign G1874 = G1812 & G54 & G1829;
  assign G1878 = ~G1876 | ~G1877;
  assign G2113 = G1958 & G1966 & G2099 & G1984;
  assign G2120 = G1966 & G1984 & G2001;
  assign G2121 = G1966 & G2099 & G1984;
  assign G2123 = G1966 & G1984 & G2001;
  assign G2124 = G1984 & G2001;
  assign G2128 = G2009 & G2021 & G2042 & G2106 & G2067;
  assign G2131 = G2009 & G2036;
  assign G2132 = G2059 & G2021 & G2009;
  assign G2133 = G2021 & G2081 & G2042 & G2009;
  assign G2134 = G2021 & G2089 & G2009 & G2067 & G2042;
  assign G2143 = G2021 & G2042 & G2081;
  assign G2144 = G2021 & G2089 & G2067 & G2042;
  assign G2145 = G2067 & G2021 & G2106 & G2042;
  assign G2147 = G2021 & G2042 & G2081;
  assign G2148 = G2021 & G2089 & G2067 & G2042;
  assign G2149 = G2042 & G2081;
  assign G2150 = G2089 & G2067 & G2042;
  assign G2151 = G2067 & G2106 & G2042;
  assign G2152 = G2042 & G2081;
  assign G2153 = G2089 & G2067 & G2042;
  assign G2154 = G2067 & G2089;
  assign G2158 = G2099 & G1984;
  assign G2159 = G2106 & G2067;
  assign G3449 = ~G3445;
  assign G3458 = ~G3454;
  assign G3472 = ~G3468;
  assign G3481 = ~G3477;
  assign G3497 = G3463;
  assign G3501 = G3463;
  assign G3505 = G3486;
  assign G3509 = G3486;
  assign G3531 = ~G5239 | ~G5242;
  assign G5428 = ~G5422;
  assign G3967 = ~G5422 | ~G5429;
  assign G4191 = G1152;
  assign G4199 = G1023;
  assign G4207 = G1023;
  assign G4215 = G1034;
  assign G4223 = G1034;
  assign G4231 = G1052;
  assign G4239 = G1052;
  assign G4247 = G1089;
  assign G4255 = G1100;
  assign G4263 = G1116;
  assign G4271 = G1134;
  assign G4371 = G1422;
  assign G4381 = G1307;
  assign G4391 = G1278;
  assign G4401 = G1289;
  assign G4429 = G1422;
  assign G4439 = G1307;
  assign G4449 = G1278;
  assign G4459 = G1289;
  assign G4497 = G1430;
  assign G4507 = G1390;
  assign G4517 = G1332;
  assign G4527 = G1365;
  assign G4537 = G1344;
  assign G4547 = G1344;
  assign G4585 = G1430;
  assign G4595 = G1390;
  assign G4605 = G1332;
  assign G4615 = G1365;
  assign G4719 = G1730;
  assign G4727 = G1730;
  assign G4735 = G1767;
  assign G4751 = G1794;
  assign G4759 = G1812;
  assign G4835 = G2099;
  assign G4845 = G1984;
  assign G4893 = G2099;
  assign G4903 = G1984;
  assign G4961 = G2067;
  assign G4971 = G2009;
  assign G4981 = G2042;
  assign G5049 = G2067;
  assign G5059 = G2009;
  assign G5069 = G2042;
  assign G5222 = ~G5216;
  assign G5223 = ~G5219;
  assign G5232 = ~G5226;
  assign G5233 = ~G5229;
  assign G5294 = ~G5289 | ~G5292;
  assign G5395 = ~G5386 | ~G5393;
  assign G589 = G1441 | G1440 | G1286 | G1439;
  assign G616 = G1847 | G1846 | G3167 | G1845;
  assign G619 = G1170 | G1169 | G1031 | G1168;
  assign G627 = G2117 | G2116 | G3167 | G2115;
  assign G1185 = G1184 | G1183 | G1182 | G1097 | G1181;
  assign G1448 = G1318 | G1447;
  assign G1458 = G1457 | G1456 | G1455 | G1341 | G1454;
  assign G1478 = G1404 | G1477;
  assign G1863 = G1862 | G1861 | G1860 | G1775 | G1859;
  assign G4747 = ~G4743;
  assign G2125 = G1995 | G2124;
  assign G2135 = G2134 | G2133 | G2132 | G2018 | G2131;
  assign G2155 = G2081 | G2154;
  assign G4995 = ~G4991;
  assign G5005 = ~G5001;
  assign G3533 = ~G3531 | ~G3532;
  assign G3921 = ~G3918;
  assign G3925 = ~G3922;
  assign G3929 = ~G3926;
  assign G3933 = ~G3930;
  assign G3943 = G3918 & G3862 & G3853;
  assign G3946 = G3922 & G3866 & G3857;
  assign G3949 = G3926 & G3883 & G3874;
  assign G3952 = G3930 & G3887 & G3878;
  assign G3966 = ~G5425 | ~G5428;
  assign G4107 = ~G4104 | ~G132;
  assign G4196 = G1173 | G1172 | G1046 | G1171;
  assign G4204 = ~G1175 & ~G1046 & ~G1174;
  assign G4212 = G1177 | G1064 | G1176;
  assign G4220 = ~G1064 & ~G1178;
  assign G4244 = G1191 | G1190 | G1189 | G1111 | G1188;
  assign G4252 = G1194 | G1193 | G1128 | G1192;
  assign G4260 = G1196 | G1145 | G1195;
  assign G4268 = G1160 | G1197;
  assign G4361 = G1444 | G1443 | G1301 | G1442;
  assign G4419 = ~G1446 & ~G1301 & ~G1445;
  assign G4467 = G1474 | G1473 | G1382 | G1472;
  assign G4487 = G1468 | G1467 | G1466 | G1359 | G1465;
  assign G4555 = ~G1476 & ~G1382 & ~G1475;
  assign G4575 = ~G1471 & ~G1470 & ~G1359 & ~G1469;
  assign G4684 = G1851 | G1850 | G1724 | G1849;
  assign G4692 = ~G1853 & ~G1724 & ~G1852;
  assign G4700 = G1855 | G1742 | G1854;
  assign G4708 = ~G1742 & ~G1856;
  assign G4732 = G1869 | G1868 | G1867 | G1789 | G1866;
  assign G4740 = G1872 | G1871 | G1806 | G1870;
  assign G4748 = G1874 | G1823 | G1873;
  assign G4825 = G2121 | G2120 | G1978 | G2119;
  assign G4883 = ~G2123 & ~G1978 & ~G2122;
  assign G4928 = G2151 | G2150 | G2059 | G2149;
  assign G4941 = G2145 | G2144 | G2143 | G2036 | G2142;
  assign G5009 = ~G2153 & ~G2059 & ~G2152;
  assign G5029 = ~G2148 & ~G2147 & ~G2036 & ~G2146;
  assign G5224 = ~G5219 | ~G5222;
  assign G5225 = ~G5216 | ~G5223;
  assign G5234 = ~G5229 | ~G5232;
  assign G5235 = ~G5226 | ~G5233;
  assign G5376 = ~G5294 | ~G5295;
  assign G5417 = ~G5394 | ~G5395;
  assign G576 = ~G1878;
  assign G588 = G1437 & G1451;
  assign G615 = G1843 & G1857;
  assign G626 = G2113 & G2128;
  assign G632 = G1166 & G1179;
  assign G1198 = ~G4191 | ~G4194;
  assign G4195 = ~G4191;
  assign G4203 = ~G4199;
  assign G4211 = ~G4207;
  assign G4219 = ~G4215;
  assign G4227 = ~G4223;
  assign G1217 = ~G4231 | ~G4234;
  assign G4235 = ~G4231;
  assign G1221 = ~G4239 | ~G4242;
  assign G4243 = ~G4239;
  assign G1224 = G1179 & G4;
  assign G4251 = ~G4247;
  assign G4259 = ~G4255;
  assign G4267 = ~G4263;
  assign G4275 = ~G4271;
  assign G1453 = ~G1451;
  assign G4405 = ~G4401;
  assign G4463 = ~G4459;
  assign G4541 = ~G4537;
  assign G4551 = ~G4547;
  assign G1895 = ~G4719 | ~G4722;
  assign G4723 = ~G4719;
  assign G1899 = ~G4727 | ~G4730;
  assign G4731 = ~G4727;
  assign G1902 = G1857 & G54;
  assign G4739 = ~G4735;
  assign G4755 = ~G4751;
  assign G1929 = ~G4759 | ~G4762;
  assign G4763 = ~G4759;
  assign G2130 = ~G2128;
  assign G3500 = ~G3497;
  assign G3504 = ~G3501;
  assign G3508 = ~G3505;
  assign G3512 = ~G3509;
  assign G3520 = G3497 & G3454 & G3445;
  assign G3523 = G3501 & G3458 & G3449;
  assign G3526 = G3505 & G3477 & G3468;
  assign G3529 = G3509 & G3481 & G3472;
  assign G1002 = G3533;
  assign G3837 = G3823 & G1878 & G3795;
  assign G3942 = G3921 & G3857 & G3862;
  assign G3945 = G3925 & G3853 & G3866;
  assign G3948 = G3929 & G3878 & G3883;
  assign G3951 = G3933 & G3874 & G3887;
  assign G3968 = ~G3966 | ~G3967;
  assign G4375 = ~G4371;
  assign G4385 = ~G4381;
  assign G4395 = ~G4391;
  assign G4433 = ~G4429;
  assign G4443 = ~G4439;
  assign G4453 = ~G4449;
  assign G4501 = ~G4497;
  assign G4511 = ~G4507;
  assign G4521 = ~G4517;
  assign G4531 = ~G4527;
  assign G4619 = ~G4615;
  assign G4589 = ~G4585;
  assign G4599 = ~G4595;
  assign G4609 = ~G4605;
  assign G4839 = ~G4835;
  assign G4849 = ~G4845;
  assign G4897 = ~G4893;
  assign G4907 = ~G4903;
  assign G4965 = ~G4961;
  assign G4975 = ~G4971;
  assign G4985 = ~G4981;
  assign G5073 = ~G5069;
  assign G5053 = ~G5049;
  assign G5063 = ~G5059;
  assign G5247 = ~G5224 | ~G5225;
  assign G5255 = ~G5234 | ~G5235;
  assign G590 = G1437 & G1458;
  assign G617 = G1863 & G1843;
  assign G620 = G1185 & G1166;
  assign G628 = G2113 & G2135;
  assign G3535 = ~G3533;
  assign G1199 = ~G4188 | ~G4195;
  assign G4202 = ~G4196;
  assign G1204 = ~G4196 | ~G4203;
  assign G4210 = ~G4204;
  assign G1207 = ~G4204 | ~G4211;
  assign G4218 = ~G4212;
  assign G1211 = ~G4212 | ~G4219;
  assign G4226 = ~G4220;
  assign G1214 = ~G4220 | ~G4227;
  assign G1218 = ~G4228 | ~G4235;
  assign G1222 = ~G4236 | ~G4243;
  assign G1225 = G1185 | G1224;
  assign G4250 = ~G4244;
  assign G1237 = ~G4244 | ~G4251;
  assign G4258 = ~G4252;
  assign G1242 = ~G4252 | ~G4259;
  assign G4266 = ~G4260;
  assign G1247 = ~G4260 | ~G4267;
  assign G4274 = ~G4268;
  assign G1252 = ~G4268 | ~G4275;
  assign G1462 = ~G1458;
  assign G4690 = ~G4684;
  assign G1882 = ~G4684 | ~G4691;
  assign G4698 = ~G4692;
  assign G1885 = ~G4692 | ~G4699;
  assign G4706 = ~G4700;
  assign G1889 = ~G4700 | ~G4707;
  assign G4714 = ~G4708;
  assign G1892 = ~G4708 | ~G4715;
  assign G1896 = ~G4716 | ~G4723;
  assign G1900 = ~G4724 | ~G4731;
  assign G1903 = G1863 | G1902;
  assign G4738 = ~G4732;
  assign G1915 = ~G4732 | ~G4739;
  assign G4746 = ~G4740;
  assign G1920 = ~G4740 | ~G4747;
  assign G4754 = ~G4748;
  assign G1925 = ~G4748 | ~G4755;
  assign G1930 = ~G4756 | ~G4763;
  assign G2139 = ~G2135;
  assign G3519 = G3500 & G3449 & G3454;
  assign G3522 = G3504 & G3445 & G3458;
  assign G3525 = G3508 & G3472 & G3477;
  assign G3528 = G3512 & G3468 & G3481;
  assign G3848 = G3838 | G3836 | G3837;
  assign G3944 = ~G3942 & ~G3943;
  assign G3947 = ~G3945 & ~G3946;
  assign G3950 = ~G3948 & ~G3949;
  assign G3953 = ~G3951 & ~G3952;
  assign G5421 = ~G5417;
  assign G1004 = G3968;
  assign G4111 = G4104 & G4107;
  assign G4112 = G4107 & G132;
  assign G4351 = G1448 | G1481;
  assign G4365 = ~G4361;
  assign G4409 = ~G1448;
  assign G4423 = ~G4419;
  assign G4471 = ~G4467;
  assign G4472 = ~G4467 | ~G4470;
  assign G4477 = G1478 | G1482;
  assign G4491 = ~G4487;
  assign G4559 = ~G4555;
  assign G4560 = ~G4555 | ~G4558;
  assign G4565 = ~G1478;
  assign G4579 = ~G4575;
  assign G4815 = G2125 | G2158;
  assign G4829 = ~G4825;
  assign G4873 = ~G2125;
  assign G4887 = ~G4883;
  assign G4931 = G2155 | G2159;
  assign G4934 = ~G4928;
  assign G4945 = ~G4941;
  assign G5013 = ~G5009;
  assign G5014 = ~G5009 | ~G5012;
  assign G5019 = ~G2155;
  assign G5033 = ~G5029;
  assign G5382 = ~G5376;
  assign G5385 = ~G5376 | ~G5383;
  assign G591 = G589 | G590;
  assign G618 = G616 | G617;
  assign G621 = G619 | G620;
  assign G629 = G627 | G628;
  assign G3970 = ~G3968;
  assign G1200 = ~G1198 | ~G1199;
  assign G1203 = ~G4199 | ~G4202;
  assign G1206 = ~G4207 | ~G4210;
  assign G1210 = ~G4215 | ~G4218;
  assign G1213 = ~G4223 | ~G4226;
  assign G1219 = ~G1217 | ~G1218;
  assign G1223 = ~G1221 | ~G1222;
  assign G1236 = ~G4247 | ~G4250;
  assign G1241 = ~G4255 | ~G4258;
  assign G1246 = ~G4263 | ~G4266;
  assign G1251 = ~G4271 | ~G4274;
  assign G1881 = ~G4687 | ~G4690;
  assign G1884 = ~G4695 | ~G4698;
  assign G1888 = ~G4703 | ~G4706;
  assign G1891 = ~G4711 | ~G4714;
  assign G1897 = ~G1895 | ~G1896;
  assign G1901 = ~G1899 | ~G1900;
  assign G1914 = ~G4735 | ~G4738;
  assign G1919 = ~G4743 | ~G4746;
  assign G1924 = ~G4751 | ~G4754;
  assign G1931 = ~G1929 | ~G1930;
  assign G3521 = ~G3519 & ~G3520;
  assign G3524 = ~G3522 & ~G3523;
  assign G3527 = ~G3525 & ~G3526;
  assign G3530 = ~G3528 & ~G3529;
  assign G5251 = ~G5247;
  assign G5259 = ~G5255;
  assign G4113 = G4111 | G4112;
  assign G4473 = ~G4464 | ~G4471;
  assign G4561 = ~G4552 | ~G4559;
  assign G5015 = ~G5006 | ~G5013;
  assign G5384 = ~G5379 | ~G5382;
  assign G5406 = ~G3947 | ~G3944;
  assign G5414 = ~G3953 | ~G3950;
  assign G1664 = G1645 & G3848 & G1621;
  assign G2335 = G2316 & G3848 & G2293;
  assign G718 = G2454 & G3848 & G2430;
  assign G822 = ~G3848;
  assign G855 = G2512 & G3848 & G2488;
  assign G1205 = ~G1203 | ~G1204;
  assign G1208 = ~G1206 | ~G1207;
  assign G1212 = ~G1210 | ~G1211;
  assign G1215 = ~G1213 | ~G1214;
  assign G1220 = ~G1219;
  assign G1231 = ~G1225;
  assign G1238 = ~G1236 | ~G1237;
  assign G1243 = ~G1241 | ~G1242;
  assign G1248 = ~G1246 | ~G1247;
  assign G1253 = ~G1251 | ~G1252;
  assign G1272 = G1225 & G1086;
  assign G1483 = G1462 & G1453;
  assign G1883 = ~G1881 | ~G1882;
  assign G1886 = ~G1884 | ~G1885;
  assign G1890 = ~G1888 | ~G1889;
  assign G1893 = ~G1891 | ~G1892;
  assign G1898 = ~G1897;
  assign G1909 = ~G1903;
  assign G1916 = ~G1914 | ~G1915;
  assign G1921 = ~G1919 | ~G1920;
  assign G1926 = ~G1924 | ~G1925;
  assign G1953 = G1903 & G1764;
  assign G2160 = G2139 & G2130;
  assign G4355 = ~G4351;
  assign G4356 = ~G4351 | ~G4354;
  assign G4413 = ~G4409;
  assign G4414 = ~G4409 | ~G4412;
  assign G4474 = ~G4472 | ~G4473;
  assign G4481 = ~G4477;
  assign G4562 = ~G4560 | ~G4561;
  assign G4569 = ~G4565;
  assign G4819 = ~G4815;
  assign G4820 = ~G4815 | ~G4818;
  assign G4877 = ~G4873;
  assign G4878 = ~G4873 | ~G4876;
  assign G4935 = ~G4931;
  assign G4936 = ~G4931 | ~G4934;
  assign G5016 = ~G5014 | ~G5015;
  assign G5023 = ~G5019;
  assign G5244 = ~G3524 | ~G3521;
  assign G5252 = ~G3530 | ~G3527;
  assign G5409 = ~G5384 | ~G5385;
  assign G566 = ~G1200;
  assign G577 = ~G1931;
  assign G3733 = G3721 & G4113 & G3724;
  assign G1209 = ~G1208;
  assign G1216 = ~G1215;
  assign G1257 = G1225 & G1205;
  assign G1262 = G1225 & G1212;
  assign G1267 = G1225 & G1220;
  assign G1887 = ~G1886;
  assign G1894 = ~G1893;
  assign G1935 = G1903 & G1883;
  assign G1943 = G1903 & G1890;
  assign G1948 = G1903 & G1898;
  assign G3779 = G3765 & G1200 & G3737;
  assign G3840 = G3823 & G1931 & G3795;
  assign G5412 = ~G5406;
  assign G5420 = ~G5414;
  assign G3964 = ~G5414 | ~G5421;
  assign G4357 = ~G4348 | ~G4355;
  assign G4415 = ~G4406 | ~G4413;
  assign G4821 = ~G4812 | ~G4819;
  assign G4879 = ~G4870 | ~G4877;
  assign G4937 = ~G4928 | ~G4935;
  assign G567 = ~G1253;
  assign G568 = ~G1248;
  assign G569 = ~G1243;
  assign G570 = ~G1238;
  assign G578 = ~G1926;
  assign G579 = ~G1921;
  assign G580 = ~G1916;
  assign G1256 = G1209 & G1231;
  assign G1261 = G1216 & G1231;
  assign G1266 = G1223 & G1231;
  assign G1271 = G1080 & G1231;
  assign G1486 = ~G1483;
  assign G1934 = G1887 & G1909;
  assign G1942 = G1894 & G1909;
  assign G1947 = G1901 & G1909;
  assign G1952 = G1758 & G1909;
  assign G2163 = ~G2160;
  assign G5250 = ~G5244;
  assign G3537 = ~G5244 | ~G5251;
  assign G5258 = ~G5252;
  assign G3542 = ~G5252 | ~G5259;
  assign G3782 = G3765 & G1253 & G3737;
  assign G3785 = G3765 & G1248 & G3737;
  assign G3788 = G3765 & G1243 & G3737;
  assign G3790 = G3780 | G3778 | G3779;
  assign G3843 = G3823 & G1926 & G3795;
  assign G3846 = G3823 & G1921 & G3795;
  assign G3849 = G3841 | G3839 | G3840;
  assign G3960 = ~G5409 | ~G5412;
  assign G5413 = ~G5409;
  assign G3963 = ~G5417 | ~G5420;
  assign G4010 = G3998 & G1238 & G3972;
  assign G4068 = G4056 & G1916 & G4030;
  assign G4358 = ~G4356 | ~G4357;
  assign G4416 = ~G4414 | ~G4415;
  assign G4480 = ~G4474;
  assign G4483 = ~G4474 | ~G4481;
  assign G4568 = ~G4562;
  assign G4571 = ~G4562 | ~G4569;
  assign G4822 = ~G4820 | ~G4821;
  assign G4880 = ~G4878 | ~G4879;
  assign G4938 = ~G4936 | ~G4937;
  assign G5022 = ~G5016;
  assign G5025 = ~G5016 | ~G5023;
  assign G1258 = G1256 | G1257;
  assign G1263 = G1261 | G1262;
  assign G1268 = G1266 | G1267;
  assign G1273 = G1271 | G1272;
  assign G1936 = G1934 | G1935;
  assign G1944 = G1942 | G1943;
  assign G1949 = G1947 | G1948;
  assign G1954 = G1952 | G1953;
  assign G3536 = ~G5247 | ~G5250;
  assign G3541 = ~G5255 | ~G5258;
  assign G3791 = G3783 | G3781 | G3782;
  assign G3792 = G3786 | G3784 | G3785;
  assign G3793 = G3789 | G3787 | G3788;
  assign G3850 = G3844 | G3842 | G3843;
  assign G3851 = G3847 | G3845 | G3846;
  assign G3961 = ~G5406 | ~G5413;
  assign G3965 = ~G3963 | ~G3964;
  assign G4024 = G4011 | G4009 | G4010;
  assign G4082 = G4069 | G4067 | G4068;
  assign G4482 = ~G4477 | ~G4480;
  assign G4570 = ~G4565 | ~G4568;
  assign G5024 = ~G5019 | ~G5022;
  assign G1666 = G1645 & G3790 & G1609;
  assign G1670 = G1645 & G3849 & G1621;
  assign G2337 = G2316 & G3790 & G2281;
  assign G2341 = G2316 & G3849 & G2293;
  assign G719 = G2454 & G3790 & G2418;
  assign G758 = G2454 & G3849 & G2430;
  assign G798 = G2512 & G3849 & G2488;
  assign G838 = ~G3849;
  assign G856 = G2512 & G3790 & G2476;
  assign G861 = ~G3790;
  assign G3538 = ~G3536 | ~G3537;
  assign G3543 = ~G3541 | ~G3542;
  assign G3962 = ~G3960 | ~G3961;
  assign G4364 = ~G4358;
  assign G4367 = ~G4358 | ~G4365;
  assign G4422 = ~G4416;
  assign G4425 = ~G4416 | ~G4423;
  assign G4484 = ~G4482 | ~G4483;
  assign G4572 = ~G4570 | ~G4571;
  assign G4828 = ~G4822;
  assign G4831 = ~G4822 | ~G4829;
  assign G4886 = ~G4880;
  assign G4889 = ~G4880 | ~G4887;
  assign G4944 = ~G4938;
  assign G4947 = ~G4938 | ~G4945;
  assign G5026 = ~G5024 | ~G5025;
  assign G571 = ~G1273;
  assign G572 = ~G1268;
  assign G573 = ~G1263;
  assign G574 = ~G1258;
  assign G581 = ~G1954;
  assign G582 = ~G1949;
  assign G583 = ~G1944;
  assign G584 = ~G1936;
  assign G623 = ~G1936;
  assign G1576 = G1564 & G4082 & G1540;
  assign G1578 = G1564 & G4024 & G1528;
  assign G659 = G1668 | G1667 | G1664 | G1666;
  assign G1672 = G1645 & G3791 & G1609;
  assign G1676 = G1645 & G3850 & G1621;
  assign G1678 = G1645 & G3792 & G1609;
  assign G1682 = G1645 & G3851 & G1621;
  assign G1684 = G1645 & G3793 & G1609;
  assign G2250 = G2238 & G4082 & G2215;
  assign G2252 = G2238 & G4024 & G2203;
  assign G691 = G2339 | G2338 | G2335 | G2337;
  assign G2343 = G2316 & G3791 & G2281;
  assign G2347 = G2316 & G3850 & G2293;
  assign G2349 = G2316 & G3792 & G2281;
  assign G2353 = G2316 & G3851 & G2293;
  assign G2355 = G2316 & G3793 & G2281;
  assign G722 = G721 | G720 | G718 | G719;
  assign G743 = G3594 & G4082 & G3570;
  assign G744 = G3594 & G4024 & G3558;
  assign G748 = G2454 & G3851 & G2430;
  assign G749 = G2454 & G3793 & G2418;
  assign G753 = G2454 & G3850 & G2430;
  assign G754 = G2454 & G3792 & G2418;
  assign G759 = G2454 & G3791 & G2418;
  assign G783 = G3696 & G4082 & G3672;
  assign G784 = G3696 & G4024 & G3660;
  assign G788 = G2512 & G3851 & G2488;
  assign G789 = G2512 & G3793 & G2476;
  assign G793 = G2512 & G3850 & G2488;
  assign G794 = G2512 & G3792 & G2476;
  assign G799 = G2512 & G3791 & G2476;
  assign G3735 = G3717 & G1936 & G3724;
  assign G832 = ~G4082;
  assign G834 = ~G3851;
  assign G836 = ~G3850;
  assign G3835 = ~G3965;
  assign G859 = G858 | G857 | G855 | G856;
  assign G871 = ~G4024;
  assign G873 = ~G3793;
  assign G875 = ~G3792;
  assign G877 = ~G3791;
  assign G998 = G3538;
  assign G1000 = G3543;
  assign G3651 = G3965 & G3632;
  assign G4013 = G3998 & G1273 & G3972;
  assign G4016 = G3998 & G1268 & G3972;
  assign G4019 = G3998 & G1263 & G3972;
  assign G4022 = G3998 & G1258 & G3972;
  assign G4071 = G4056 & G1954 & G4030;
  assign G4074 = G4056 & G1949 & G4030;
  assign G4077 = G4056 & G1944 & G4030;
  assign G4080 = G4056 & G1936 & G4030;
  assign G4096 = ~G4113 | ~G1936;
  assign G4366 = ~G4361 | ~G4364;
  assign G4424 = ~G4419 | ~G4422;
  assign G4830 = ~G4825 | ~G4828;
  assign G4888 = ~G4883 | ~G4886;
  assign G4946 = ~G4941 | ~G4944;
  assign G575 = G574 & G573 & G572 & G571 & G570 & G569 & G568 & G566 & G567;
  assign G585 = G584 & G583 & G582 & G581 & G580 & G579 & G578 & G576 & G577;
  assign G640 = G1580 | G1579 | G1576 | G1578;
  assign G661 = G659 & G1606;
  assign G662 = G1674 | G1673 | G1670 | G1672;
  assign G665 = G1680 | G1679 | G1676 | G1678;
  assign G668 = G1686 | G1685 | G1682 | G1684;
  assign G674 = G2254 | G2253 | G2250 | G2252;
  assign G693 = G691 & G2279;
  assign G694 = G2345 | G2344 | G2341 | G2343;
  assign G697 = G2351 | G2350 | G2347 | G2349;
  assign G700 = G2357 | G2356 | G2353 | G2355;
  assign G747 = G746 | G745 | G743 | G744;
  assign G752 = G751 | G750 | G748 | G749;
  assign G757 = G756 | G755 | G753 | G754;
  assign G762 = G761 | G760 | G758 | G759;
  assign G787 = G786 | G785 | G783 | G784;
  assign G792 = G791 | G790 | G788 | G789;
  assign G797 = G796 | G795 | G793 | G794;
  assign G802 = G801 | G800 | G798 | G799;
  assign G817 = G3735 | G3734 | G3731 | G3733;
  assign G839 = G3823 & G3835 & G3803;
  assign G3540 = ~G3538;
  assign G3545 = ~G3543;
  assign G3777 = ~G3962;
  assign G3648 = G3962 & G3632;
  assign G4025 = G4014 | G4012 | G4013;
  assign G4026 = G4017 | G4015 | G4016;
  assign G4027 = G4020 | G4018 | G4019;
  assign G4028 = G4023 | G4021 | G4022;
  assign G4083 = G4072 | G4070 | G4071;
  assign G4084 = G4075 | G4073 | G4074;
  assign G4085 = G4078 | G4076 | G4077;
  assign G4086 = G4081 | G4079 | G4080;
  assign G4368 = ~G4366 | ~G4367;
  assign G4426 = ~G4424 | ~G4425;
  assign G4490 = ~G4484;
  assign G4493 = ~G4484 | ~G4491;
  assign G4578 = ~G4572;
  assign G4581 = ~G4572 | ~G4579;
  assign G4832 = ~G4830 | ~G4831;
  assign G4890 = ~G4888 | ~G4889;
  assign G4948 = ~G4946 | ~G4947;
  assign G5032 = ~G5026;
  assign G5035 = ~G5026 | ~G5033;
  assign G642 = G640 & G1526;
  assign G664 = G662 & G1606;
  assign G667 = G665 & G1606;
  assign G670 = G668 & G1606;
  assign G676 = G674 & G2202;
  assign G696 = G694 & G2279;
  assign G699 = G697 & G2279;
  assign G702 = G700 & G2279;
  assign G811 = G4113 & G4096;
  assign G812 = G4096 & G1936;
  assign G818 = G816 & G817;
  assign G853 = G3970 & G3535 & G3545 & G562 & G3540;
  assign G878 = G3765 & G3777 & G3745;
  assign G4492 = ~G4487 | ~G4490;
  assign G4580 = ~G4575 | ~G4578;
  assign G5034 = ~G5029 | ~G5032;
  assign G1582 = G1564 & G4083 & G1540;
  assign G1584 = G1564 & G4025 & G1528;
  assign G1588 = G1564 & G4084 & G1540;
  assign G1590 = G1564 & G4026 & G1528;
  assign G1594 = G1564 & G4085 & G1540;
  assign G1596 = G1564 & G4027 & G1528;
  assign G1600 = G1564 & G4086 & G1540;
  assign G1602 = G1564 & G4028 & G1528;
  assign G2256 = G2238 & G4083 & G2215;
  assign G2258 = G2238 & G4025 & G2203;
  assign G2262 = G2238 & G4084 & G2215;
  assign G2264 = G2238 & G4026 & G2203;
  assign G2268 = G2238 & G4085 & G2215;
  assign G2270 = G2238 & G4027 & G2203;
  assign G2274 = G2238 & G4086 & G2215;
  assign G2276 = G2238 & G4028 & G2203;
  assign G708 = G3696 & G4086 & G3672;
  assign G709 = G3696 & G4028 & G3660;
  assign G723 = G3594 & G4086 & G3570;
  assign G724 = G3594 & G4028 & G3558;
  assign G728 = G3594 & G4085 & G3570;
  assign G729 = G3594 & G4027 & G3558;
  assign G733 = G3594 & G4084 & G3570;
  assign G734 = G3594 & G4026 & G3558;
  assign G738 = G3594 & G4083 & G3570;
  assign G739 = G3594 & G4025 & G3558;
  assign G768 = G3696 & G4085 & G3672;
  assign G769 = G3696 & G4027 & G3660;
  assign G773 = G3696 & G4084 & G3672;
  assign G774 = G3696 & G4026 & G3660;
  assign G778 = G3696 & G4083 & G3672;
  assign G779 = G3696 & G4025 & G3660;
  assign G813 = G811 | G812;
  assign G824 = ~G4086;
  assign G826 = ~G4085;
  assign G828 = ~G4084;
  assign G830 = ~G4083;
  assign G854 = G245 & G852 & G853;
  assign G863 = ~G4028;
  assign G865 = ~G4027;
  assign G867 = ~G4026;
  assign G869 = ~G4025;
  assign G4374 = ~G4368;
  assign G4377 = ~G4368 | ~G4375;
  assign G4432 = ~G4426;
  assign G4435 = ~G4426 | ~G4433;
  assign G4494 = ~G4492 | ~G4493;
  assign G4582 = ~G4580 | ~G4581;
  assign G4838 = ~G4832;
  assign G4841 = ~G4832 | ~G4839;
  assign G4896 = ~G4890;
  assign G4899 = ~G4890 | ~G4897;
  assign G4954 = ~G4948;
  assign G4957 = ~G4948 | ~G4955;
  assign G5036 = ~G5034 | ~G5035;
  assign G643 = G1586 | G1585 | G1582 | G1584;
  assign G646 = G1592 | G1591 | G1588 | G1590;
  assign G649 = G1598 | G1597 | G1594 | G1596;
  assign G652 = G1604 | G1603 | G1600 | G1602;
  assign G677 = G2260 | G2259 | G2256 | G2258;
  assign G680 = G2266 | G2265 | G2262 | G2264;
  assign G683 = G2272 | G2271 | G2268 | G2270;
  assign G686 = G2278 | G2277 | G2274 | G2276;
  assign G712 = G711 | G710 | G708 | G709;
  assign G727 = G726 | G725 | G723 | G724;
  assign G732 = G731 | G730 | G728 | G729;
  assign G737 = G736 | G735 | G733 | G734;
  assign G742 = G741 | G740 | G738 | G739;
  assign G772 = G771 | G770 | G768 | G769;
  assign G777 = G776 | G775 | G773 | G774;
  assign G782 = G781 | G780 | G778 | G779;
  assign G4376 = ~G4371 | ~G4374;
  assign G4434 = ~G4429 | ~G4432;
  assign G4840 = ~G4835 | ~G4838;
  assign G4898 = ~G4893 | ~G4896;
  assign G4956 = ~G4951 | ~G4954;
  assign G645 = G643 & G1526;
  assign G648 = G646 & G1526;
  assign G651 = G649 & G1526;
  assign G654 = G652 & G1526;
  assign G679 = G677 & G2202;
  assign G682 = G680 & G2202;
  assign G685 = G683 & G2202;
  assign G688 = G686 & G2202;
  assign G4378 = ~G4376 | ~G4377;
  assign G4436 = ~G4434 | ~G4435;
  assign G4500 = ~G4494;
  assign G4503 = ~G4494 | ~G4501;
  assign G4588 = ~G4582;
  assign G4591 = ~G4582 | ~G4589;
  assign G4842 = ~G4840 | ~G4841;
  assign G4900 = ~G4898 | ~G4899;
  assign G4958 = ~G4956 | ~G4957;
  assign G5042 = ~G5036;
  assign G5045 = ~G5036 | ~G5043;
  assign G4502 = ~G4497 | ~G4500;
  assign G4590 = ~G4585 | ~G4588;
  assign G5044 = ~G5039 | ~G5042;
  assign G4384 = ~G4378;
  assign G4387 = ~G4378 | ~G4385;
  assign G4442 = ~G4436;
  assign G4445 = ~G4436 | ~G4443;
  assign G4504 = ~G4502 | ~G4503;
  assign G4592 = ~G4590 | ~G4591;
  assign G4848 = ~G4842;
  assign G4851 = ~G4842 | ~G4849;
  assign G4906 = ~G4900;
  assign G4909 = ~G4900 | ~G4907;
  assign G4964 = ~G4958;
  assign G4967 = ~G4958 | ~G4965;
  assign G5046 = ~G5044 | ~G5045;
  assign G4386 = ~G4381 | ~G4384;
  assign G4444 = ~G4439 | ~G4442;
  assign G4850 = ~G4845 | ~G4848;
  assign G4908 = ~G4903 | ~G4906;
  assign G4966 = ~G4961 | ~G4964;
  assign G4388 = ~G4386 | ~G4387;
  assign G4446 = ~G4444 | ~G4445;
  assign G4510 = ~G4504;
  assign G4513 = ~G4504 | ~G4511;
  assign G4598 = ~G4592;
  assign G4601 = ~G4592 | ~G4599;
  assign G4852 = ~G4850 | ~G4851;
  assign G4910 = ~G4908 | ~G4909;
  assign G4968 = ~G4966 | ~G4967;
  assign G5052 = ~G5046;
  assign G5055 = ~G5046 | ~G5053;
  assign G4512 = ~G4507 | ~G4510;
  assign G4600 = ~G4595 | ~G4598;
  assign G5054 = ~G5049 | ~G5052;
  assign G4394 = ~G4388;
  assign G4397 = ~G4388 | ~G4395;
  assign G4452 = ~G4446;
  assign G4455 = ~G4446 | ~G4453;
  assign G4514 = ~G4512 | ~G4513;
  assign G4602 = ~G4600 | ~G4601;
  assign G4858 = ~G4852;
  assign G4861 = ~G4852 | ~G4859;
  assign G4916 = ~G4910;
  assign G4919 = ~G4910 | ~G4917;
  assign G4974 = ~G4968;
  assign G4977 = ~G4968 | ~G4975;
  assign G5056 = ~G5054 | ~G5055;
  assign G4396 = ~G4391 | ~G4394;
  assign G4454 = ~G4449 | ~G4452;
  assign G4860 = ~G4855 | ~G4858;
  assign G4918 = ~G4913 | ~G4916;
  assign G4976 = ~G4971 | ~G4974;
  assign G4398 = ~G4396 | ~G4397;
  assign G4456 = ~G4454 | ~G4455;
  assign G4520 = ~G4514;
  assign G4523 = ~G4514 | ~G4521;
  assign G4608 = ~G4602;
  assign G4611 = ~G4602 | ~G4609;
  assign G4862 = ~G4860 | ~G4861;
  assign G4920 = ~G4918 | ~G4919;
  assign G4978 = ~G4976 | ~G4977;
  assign G5062 = ~G5056;
  assign G5065 = ~G5056 | ~G5063;
  assign G4522 = ~G4517 | ~G4520;
  assign G4610 = ~G4605 | ~G4608;
  assign G5064 = ~G5059 | ~G5062;
  assign G4404 = ~G4398;
  assign G1488 = ~G4398 | ~G4405;
  assign G4462 = ~G4456;
  assign G1493 = ~G4456 | ~G4463;
  assign G4868 = ~G4862;
  assign G2165 = ~G4862 | ~G4869;
  assign G4926 = ~G4920;
  assign G2170 = ~G4920 | ~G4927;
  assign G4524 = ~G4522 | ~G4523;
  assign G4612 = ~G4610 | ~G4611;
  assign G4984 = ~G4978;
  assign G4987 = ~G4978 | ~G4985;
  assign G5066 = ~G5064 | ~G5065;
  assign G1487 = ~G4401 | ~G4404;
  assign G1492 = ~G4459 | ~G4462;
  assign G2164 = ~G4865 | ~G4868;
  assign G2169 = ~G4923 | ~G4926;
  assign G4986 = ~G4981 | ~G4984;
  assign G1489 = ~G1487 | ~G1488;
  assign G1494 = ~G1492 | ~G1493;
  assign G2166 = ~G2164 | ~G2165;
  assign G2171 = ~G2169 | ~G2170;
  assign G4530 = ~G4524;
  assign G4533 = ~G4524 | ~G4531;
  assign G4618 = ~G4612;
  assign G4543 = ~G4612 | ~G4619;
  assign G4988 = ~G4986 | ~G4987;
  assign G5072 = ~G5066;
  assign G4997 = ~G5066 | ~G5073;
  assign G4532 = ~G4527 | ~G4530;
  assign G4542 = ~G4615 | ~G4618;
  assign G4996 = ~G5069 | ~G5072;
  assign G1513 = G1502 & G1494 & G1462;
  assign G1514 = G1502 & G1489 & G1458;
  assign G1515 = G1497 & G1494 & G1483;
  assign G1516 = G1497 & G1489 & G1486;
  assign G4994 = ~G4988;
  assign G2184 = ~G4988 | ~G4995;
  assign G2190 = G2179 & G2171 & G2139;
  assign G2191 = G2179 & G2166 & G2135;
  assign G2192 = G2174 & G2171 & G2160;
  assign G2193 = G2174 & G2166 & G2163;
  assign G4534 = ~G4532 | ~G4533;
  assign G4544 = ~G4542 | ~G4543;
  assign G4998 = ~G4996 | ~G4997;
  assign G2183 = ~G4991 | ~G4994;
  assign G4620 = G1516 | G1515 | G1513 | G1514;
  assign G5074 = G2193 | G2192 | G2190 | G2191;
  assign G4540 = ~G4534;
  assign G1507 = ~G4534 | ~G4541;
  assign G4550 = ~G4544;
  assign G1510 = ~G4544 | ~G4551;
  assign G2185 = ~G2183 | ~G2184;
  assign G5004 = ~G4998;
  assign G2187 = ~G4998 | ~G5005;
  assign G1506 = ~G4537 | ~G4540;
  assign G1509 = ~G4547 | ~G4550;
  assign G4626 = ~G4620;
  assign G2186 = ~G5001 | ~G5004;
  assign G2195 = G2174 & G2185;
  assign G5080 = ~G5074;
  assign G1508 = ~G1506 | ~G1507;
  assign G1511 = ~G1509 | ~G1510;
  assign G2188 = ~G2186 | ~G2187;
  assign G1512 = ~G1511;
  assign G1518 = G1497 & G1508;
  assign G2189 = ~G2188;
  assign G1517 = G1512 & G1502;
  assign G2194 = G2189 & G2179;
  assign G4623 = G1517 | G1518;
  assign G5077 = G2194 | G2195;
  assign G1519 = ~G4623 | ~G4626;
  assign G4627 = ~G4623;
  assign G2196 = ~G5077 | ~G5080;
  assign G5081 = ~G5077;
  assign G1520 = ~G4620 | ~G4627;
  assign G2197 = ~G5074 | ~G5081;
  assign G1521 = ~G1519 | ~G1520;
  assign G2198 = ~G2196 | ~G2197;
  assign G840 = G3823 & G2198 & G3795;
  assign G879 = G3765 & G1521 & G3737;
  assign G1524 = ~G1521;
  assign G2201 = ~G2198;
  assign G843 = G842 | G841 | G839 | G840;
  assign G882 = G881 | G880 | G878 | G879;
  assign G3649 = G1524 & G3628;
  assign G3652 = G2201 & G3628;
  assign G3657 = G3648 | G3649;
  assign G3658 = G3651 | G3652;
  assign G3636 = G3657 & G3622;
  assign G3639 = G3658 & G3622;
  assign G3642 = G3657 & G3622;
  assign G3645 = G3658 & G3622;
  assign G3653 = G3636 | G3637;
  assign G3654 = G3639 | G3640;
  assign G3655 = G3642 | G3643;
  assign G3656 = G3645 | G3646;
  assign G763 = G2454 & G3656 & G2430;
  assign G764 = G2454 & G3655 & G2418;
  assign G803 = G2512 & G3656 & G2488;
  assign G804 = G2512 & G3655 & G2476;
  assign G1657 = G1645 & G3654 & G1621;
  assign G1659 = G1645 & G3653 & G1609;
  assign G2328 = G2316 & G3654 & G2293;
  assign G2330 = G2316 & G3653 & G2281;
  assign G1662 = G1661 | G1660 | G1657 | G1659;
  assign G2333 = G2332 | G2331 | G2328 | G2330;
  assign G767 = G766 | G765 | G763 | G764;
  assign G807 = G806 | G805 | G803 | G804;
  assign G657 = G1662 & G1606;
  assign G689 = G2333 & G2279;
  assign G658 = ~G657;
  assign G690 = ~G689;
endmodule


