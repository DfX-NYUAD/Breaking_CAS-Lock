// Benchmark "b18_C_lock" written by ABC on Thu May 13 23:53:21 2021

module b18_C_lock ( 
    keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
    keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
    keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
    keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
    keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
    keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
    keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
    keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
    keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
    keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
    keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
    keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
    keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
    keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
    keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
    keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
    keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
    keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
    keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
    keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
    keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
    keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
    keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
    keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
    keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
    keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
    keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
    keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
    keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
    keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
    keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
    keyinput_156, keyinput_157, keyinput_158, keyinput_159, SEL, DIN_30_,
    DIN_29_, DIN_28_, DIN_27_, DIN_26_, DIN_25_, DIN_24_, DIN_23_, DIN_22_,
    DIN_21_, DIN_20_, DIN_19_, DIN_18_, DIN_17_, DIN_16_, DIN_15_, DIN_14_,
    DIN_13_, DIN_12_, DIN_11_, DIN_10_, DIN_9_, DIN_8_, DIN_7_, DIN_6_,
    DIN_5_, DIN_4_, DIN_3_, DIN_2_, DIN_1_, DIN_0_,
    P2_P1_ADS_N_REG_SCAN_IN, P1_BUF1_REG_14__SCAN_IN,
    P1_BUF1_REG_30__SCAN_IN, P1_READY11_REG_SCAN_IN,
    P4_DATAO_REG_0__SCAN_IN, P4_DATAO_REG_1__SCAN_IN,
    P4_DATAO_REG_2__SCAN_IN, P4_DATAO_REG_3__SCAN_IN,
    P4_DATAO_REG_4__SCAN_IN, P4_DATAO_REG_5__SCAN_IN,
    P4_DATAO_REG_6__SCAN_IN, P4_DATAO_REG_7__SCAN_IN,
    P4_DATAO_REG_8__SCAN_IN, P4_DATAO_REG_9__SCAN_IN,
    P4_DATAO_REG_10__SCAN_IN, P4_DATAO_REG_11__SCAN_IN,
    P4_DATAO_REG_12__SCAN_IN, P4_DATAO_REG_13__SCAN_IN,
    P4_DATAO_REG_14__SCAN_IN, P4_DATAO_REG_15__SCAN_IN,
    P4_DATAO_REG_16__SCAN_IN, P4_DATAO_REG_17__SCAN_IN,
    P4_DATAO_REG_18__SCAN_IN, P4_DATAO_REG_19__SCAN_IN,
    P4_DATAO_REG_20__SCAN_IN, P4_DATAO_REG_21__SCAN_IN,
    P4_DATAO_REG_22__SCAN_IN, P4_DATAO_REG_23__SCAN_IN,
    P4_DATAO_REG_24__SCAN_IN, P4_DATAO_REG_25__SCAN_IN,
    P4_DATAO_REG_26__SCAN_IN, P4_DATAO_REG_27__SCAN_IN,
    P4_DATAO_REG_28__SCAN_IN, P4_DATAO_REG_29__SCAN_IN,
    P4_DATAO_REG_30__SCAN_IN, P1_P1_ADDRESS_REG_29__SCAN_IN,
    P1_P1_ADDRESS_REG_28__SCAN_IN, P1_P1_ADDRESS_REG_27__SCAN_IN,
    P1_P1_ADDRESS_REG_26__SCAN_IN, P1_P1_ADDRESS_REG_25__SCAN_IN,
    P1_P1_ADDRESS_REG_24__SCAN_IN, P1_P1_ADDRESS_REG_23__SCAN_IN,
    P1_P1_ADDRESS_REG_22__SCAN_IN, P1_P1_ADDRESS_REG_21__SCAN_IN,
    P1_P1_ADDRESS_REG_20__SCAN_IN, P1_P1_ADDRESS_REG_19__SCAN_IN,
    P1_P1_ADDRESS_REG_18__SCAN_IN, P1_P1_ADDRESS_REG_17__SCAN_IN,
    P1_P1_ADDRESS_REG_16__SCAN_IN, P1_P1_ADDRESS_REG_15__SCAN_IN,
    P1_P1_ADDRESS_REG_14__SCAN_IN, P1_P1_ADDRESS_REG_13__SCAN_IN,
    P1_P1_ADDRESS_REG_12__SCAN_IN, P1_P1_ADDRESS_REG_11__SCAN_IN,
    P1_P1_ADDRESS_REG_10__SCAN_IN, P1_P1_ADDRESS_REG_9__SCAN_IN,
    P1_P1_ADDRESS_REG_8__SCAN_IN, P1_P1_ADDRESS_REG_7__SCAN_IN,
    P1_P1_ADDRESS_REG_6__SCAN_IN, P1_P1_ADDRESS_REG_5__SCAN_IN,
    P1_P1_ADDRESS_REG_4__SCAN_IN, P1_P1_ADDRESS_REG_3__SCAN_IN,
    P1_P1_ADDRESS_REG_2__SCAN_IN, P1_P1_ADDRESS_REG_1__SCAN_IN,
    P1_P1_ADDRESS_REG_0__SCAN_IN, P1_P1_STATE2_REG_2__SCAN_IN,
    P1_P1_STATE2_REG_1__SCAN_IN, P1_P1_STATE2_REG_0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_P1_INSTQUEUE_REG_15__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_P1_INSTQUEUE_REG_15__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_P1_INSTQUEUE_REG_15__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_P1_INSTQUEUE_REG_15__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_P1_INSTQUEUE_REG_14__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_P1_INSTQUEUE_REG_14__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_P1_INSTQUEUE_REG_14__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_P1_INSTQUEUE_REG_14__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_P1_INSTQUEUE_REG_13__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_P1_INSTQUEUE_REG_13__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_P1_INSTQUEUE_REG_13__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_P1_INSTQUEUE_REG_13__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_P1_INSTQUEUE_REG_12__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_P1_INSTQUEUE_REG_12__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_P1_INSTQUEUE_REG_12__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_P1_INSTQUEUE_REG_12__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_P1_INSTQUEUE_REG_11__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_P1_INSTQUEUE_REG_11__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_P1_INSTQUEUE_REG_11__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_P1_INSTQUEUE_REG_11__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_P1_INSTQUEUE_REG_10__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_P1_INSTQUEUE_REG_10__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_P1_INSTQUEUE_REG_10__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_P1_INSTQUEUE_REG_10__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_P1_INSTQUEUE_REG_9__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_P1_INSTQUEUE_REG_9__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_P1_INSTQUEUE_REG_9__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_P1_INSTQUEUE_REG_9__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_P1_INSTQUEUE_REG_8__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_P1_INSTQUEUE_REG_8__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_P1_INSTQUEUE_REG_8__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_P1_INSTQUEUE_REG_8__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_P1_INSTQUEUE_REG_7__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_P1_INSTQUEUE_REG_7__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_P1_INSTQUEUE_REG_7__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_P1_INSTQUEUE_REG_7__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_P1_INSTQUEUE_REG_6__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_P1_INSTQUEUE_REG_6__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_P1_INSTQUEUE_REG_6__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_P1_INSTQUEUE_REG_6__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_P1_INSTQUEUE_REG_5__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_P1_INSTQUEUE_REG_5__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_P1_INSTQUEUE_REG_5__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_P1_INSTQUEUE_REG_5__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_P1_INSTQUEUE_REG_4__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_P1_INSTQUEUE_REG_4__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_P1_INSTQUEUE_REG_4__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_4__1__SCAN_IN, P1_P1_INSTQUEUE_REG_4__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_P1_INSTQUEUE_REG_3__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_P1_INSTQUEUE_REG_3__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_P1_INSTQUEUE_REG_3__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_P1_INSTQUEUE_REG_3__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_P1_INSTQUEUE_REG_2__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_P1_INSTQUEUE_REG_2__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_P1_INSTQUEUE_REG_2__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_P1_INSTQUEUE_REG_2__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_P1_INSTQUEUE_REG_1__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_P1_INSTQUEUE_REG_1__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_P1_INSTQUEUE_REG_1__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_P1_INSTQUEUE_REG_1__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_P1_INSTQUEUE_REG_0__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_P1_INSTQUEUE_REG_0__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_P1_INSTQUEUE_REG_0__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_P1_INSTQUEUE_REG_0__0__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_P1_EAX_REG_0__SCAN_IN,
    P1_P1_EAX_REG_1__SCAN_IN, P1_P1_EAX_REG_2__SCAN_IN,
    P1_P1_EAX_REG_3__SCAN_IN, P1_P1_EAX_REG_4__SCAN_IN,
    P1_P1_EAX_REG_5__SCAN_IN, P1_P1_EAX_REG_6__SCAN_IN,
    P1_P1_EAX_REG_7__SCAN_IN, P1_P1_EAX_REG_8__SCAN_IN,
    P1_P1_EAX_REG_9__SCAN_IN, P1_P1_EAX_REG_10__SCAN_IN,
    P1_P1_EAX_REG_11__SCAN_IN, P1_P1_EAX_REG_12__SCAN_IN,
    P1_P1_EAX_REG_13__SCAN_IN, P1_P1_EAX_REG_14__SCAN_IN,
    P1_P1_EAX_REG_15__SCAN_IN, P1_P1_EAX_REG_16__SCAN_IN,
    P1_P1_EAX_REG_17__SCAN_IN, P1_P1_EAX_REG_18__SCAN_IN,
    P1_P1_EAX_REG_19__SCAN_IN, P1_P1_EAX_REG_20__SCAN_IN,
    P1_P1_EAX_REG_21__SCAN_IN, P1_P1_EAX_REG_22__SCAN_IN,
    P1_P1_EAX_REG_23__SCAN_IN, P1_P1_EAX_REG_24__SCAN_IN,
    P1_P1_EAX_REG_25__SCAN_IN, P1_P1_EAX_REG_26__SCAN_IN,
    P1_P1_EAX_REG_27__SCAN_IN, P1_P1_EAX_REG_28__SCAN_IN,
    P1_P1_EAX_REG_29__SCAN_IN, P1_P1_EAX_REG_30__SCAN_IN,
    P1_P1_U2721  );
  input  keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4,
    keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9,
    keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14,
    keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19,
    keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24,
    keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29,
    keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34,
    keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39,
    keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44,
    keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49,
    keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54,
    keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59,
    keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64,
    keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69,
    keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74,
    keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79,
    keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84,
    keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89,
    keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94,
    keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99,
    keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104,
    keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109,
    keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114,
    keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119,
    keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124,
    keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129,
    keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134,
    keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139,
    keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144,
    keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149,
    keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154,
    keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159,
    SEL, DIN_30_, DIN_29_, DIN_28_, DIN_27_, DIN_26_, DIN_25_, DIN_24_,
    DIN_23_, DIN_22_, DIN_21_, DIN_20_, DIN_19_, DIN_18_, DIN_17_, DIN_16_,
    DIN_15_, DIN_14_, DIN_13_, DIN_12_, DIN_11_, DIN_10_, DIN_9_, DIN_8_,
    DIN_7_, DIN_6_, DIN_5_, DIN_4_, DIN_3_, DIN_2_, DIN_1_, DIN_0_,
    P2_P1_ADS_N_REG_SCAN_IN, P1_BUF1_REG_14__SCAN_IN,
    P1_BUF1_REG_30__SCAN_IN, P1_READY11_REG_SCAN_IN,
    P4_DATAO_REG_0__SCAN_IN, P4_DATAO_REG_1__SCAN_IN,
    P4_DATAO_REG_2__SCAN_IN, P4_DATAO_REG_3__SCAN_IN,
    P4_DATAO_REG_4__SCAN_IN, P4_DATAO_REG_5__SCAN_IN,
    P4_DATAO_REG_6__SCAN_IN, P4_DATAO_REG_7__SCAN_IN,
    P4_DATAO_REG_8__SCAN_IN, P4_DATAO_REG_9__SCAN_IN,
    P4_DATAO_REG_10__SCAN_IN, P4_DATAO_REG_11__SCAN_IN,
    P4_DATAO_REG_12__SCAN_IN, P4_DATAO_REG_13__SCAN_IN,
    P4_DATAO_REG_14__SCAN_IN, P4_DATAO_REG_15__SCAN_IN,
    P4_DATAO_REG_16__SCAN_IN, P4_DATAO_REG_17__SCAN_IN,
    P4_DATAO_REG_18__SCAN_IN, P4_DATAO_REG_19__SCAN_IN,
    P4_DATAO_REG_20__SCAN_IN, P4_DATAO_REG_21__SCAN_IN,
    P4_DATAO_REG_22__SCAN_IN, P4_DATAO_REG_23__SCAN_IN,
    P4_DATAO_REG_24__SCAN_IN, P4_DATAO_REG_25__SCAN_IN,
    P4_DATAO_REG_26__SCAN_IN, P4_DATAO_REG_27__SCAN_IN,
    P4_DATAO_REG_28__SCAN_IN, P4_DATAO_REG_29__SCAN_IN,
    P4_DATAO_REG_30__SCAN_IN, P1_P1_ADDRESS_REG_29__SCAN_IN,
    P1_P1_ADDRESS_REG_28__SCAN_IN, P1_P1_ADDRESS_REG_27__SCAN_IN,
    P1_P1_ADDRESS_REG_26__SCAN_IN, P1_P1_ADDRESS_REG_25__SCAN_IN,
    P1_P1_ADDRESS_REG_24__SCAN_IN, P1_P1_ADDRESS_REG_23__SCAN_IN,
    P1_P1_ADDRESS_REG_22__SCAN_IN, P1_P1_ADDRESS_REG_21__SCAN_IN,
    P1_P1_ADDRESS_REG_20__SCAN_IN, P1_P1_ADDRESS_REG_19__SCAN_IN,
    P1_P1_ADDRESS_REG_18__SCAN_IN, P1_P1_ADDRESS_REG_17__SCAN_IN,
    P1_P1_ADDRESS_REG_16__SCAN_IN, P1_P1_ADDRESS_REG_15__SCAN_IN,
    P1_P1_ADDRESS_REG_14__SCAN_IN, P1_P1_ADDRESS_REG_13__SCAN_IN,
    P1_P1_ADDRESS_REG_12__SCAN_IN, P1_P1_ADDRESS_REG_11__SCAN_IN,
    P1_P1_ADDRESS_REG_10__SCAN_IN, P1_P1_ADDRESS_REG_9__SCAN_IN,
    P1_P1_ADDRESS_REG_8__SCAN_IN, P1_P1_ADDRESS_REG_7__SCAN_IN,
    P1_P1_ADDRESS_REG_6__SCAN_IN, P1_P1_ADDRESS_REG_5__SCAN_IN,
    P1_P1_ADDRESS_REG_4__SCAN_IN, P1_P1_ADDRESS_REG_3__SCAN_IN,
    P1_P1_ADDRESS_REG_2__SCAN_IN, P1_P1_ADDRESS_REG_1__SCAN_IN,
    P1_P1_ADDRESS_REG_0__SCAN_IN, P1_P1_STATE2_REG_2__SCAN_IN,
    P1_P1_STATE2_REG_1__SCAN_IN, P1_P1_STATE2_REG_0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_P1_INSTQUEUE_REG_15__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_P1_INSTQUEUE_REG_15__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_P1_INSTQUEUE_REG_15__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_P1_INSTQUEUE_REG_15__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_P1_INSTQUEUE_REG_14__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_P1_INSTQUEUE_REG_14__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_P1_INSTQUEUE_REG_14__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_P1_INSTQUEUE_REG_14__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_P1_INSTQUEUE_REG_13__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_P1_INSTQUEUE_REG_13__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_P1_INSTQUEUE_REG_13__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_P1_INSTQUEUE_REG_13__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_P1_INSTQUEUE_REG_12__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_P1_INSTQUEUE_REG_12__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_P1_INSTQUEUE_REG_12__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_P1_INSTQUEUE_REG_12__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_P1_INSTQUEUE_REG_11__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_P1_INSTQUEUE_REG_11__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_P1_INSTQUEUE_REG_11__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_P1_INSTQUEUE_REG_11__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_P1_INSTQUEUE_REG_10__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_P1_INSTQUEUE_REG_10__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_P1_INSTQUEUE_REG_10__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_P1_INSTQUEUE_REG_10__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_P1_INSTQUEUE_REG_9__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_P1_INSTQUEUE_REG_9__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_P1_INSTQUEUE_REG_9__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_P1_INSTQUEUE_REG_9__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_P1_INSTQUEUE_REG_8__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_P1_INSTQUEUE_REG_8__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_P1_INSTQUEUE_REG_8__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_P1_INSTQUEUE_REG_8__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_P1_INSTQUEUE_REG_7__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_P1_INSTQUEUE_REG_7__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_P1_INSTQUEUE_REG_7__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_P1_INSTQUEUE_REG_7__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_P1_INSTQUEUE_REG_6__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_P1_INSTQUEUE_REG_6__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_P1_INSTQUEUE_REG_6__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_P1_INSTQUEUE_REG_6__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_P1_INSTQUEUE_REG_5__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_P1_INSTQUEUE_REG_5__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_P1_INSTQUEUE_REG_5__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_P1_INSTQUEUE_REG_5__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_P1_INSTQUEUE_REG_4__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_P1_INSTQUEUE_REG_4__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_P1_INSTQUEUE_REG_4__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_4__1__SCAN_IN, P1_P1_INSTQUEUE_REG_4__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_P1_INSTQUEUE_REG_3__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_P1_INSTQUEUE_REG_3__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_P1_INSTQUEUE_REG_3__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_P1_INSTQUEUE_REG_3__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_P1_INSTQUEUE_REG_2__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_P1_INSTQUEUE_REG_2__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_P1_INSTQUEUE_REG_2__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_P1_INSTQUEUE_REG_2__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_P1_INSTQUEUE_REG_1__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_P1_INSTQUEUE_REG_1__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_P1_INSTQUEUE_REG_1__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_P1_INSTQUEUE_REG_1__0__SCAN_IN,
    P1_P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_P1_INSTQUEUE_REG_0__6__SCAN_IN,
    P1_P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_P1_INSTQUEUE_REG_0__4__SCAN_IN,
    P1_P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_P1_INSTQUEUE_REG_0__2__SCAN_IN,
    P1_P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_P1_INSTQUEUE_REG_0__0__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    P1_P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_P1_EAX_REG_0__SCAN_IN,
    P1_P1_EAX_REG_1__SCAN_IN, P1_P1_EAX_REG_2__SCAN_IN,
    P1_P1_EAX_REG_3__SCAN_IN, P1_P1_EAX_REG_4__SCAN_IN,
    P1_P1_EAX_REG_5__SCAN_IN, P1_P1_EAX_REG_6__SCAN_IN,
    P1_P1_EAX_REG_7__SCAN_IN, P1_P1_EAX_REG_8__SCAN_IN,
    P1_P1_EAX_REG_9__SCAN_IN, P1_P1_EAX_REG_10__SCAN_IN,
    P1_P1_EAX_REG_11__SCAN_IN, P1_P1_EAX_REG_12__SCAN_IN,
    P1_P1_EAX_REG_13__SCAN_IN, P1_P1_EAX_REG_14__SCAN_IN,
    P1_P1_EAX_REG_15__SCAN_IN, P1_P1_EAX_REG_16__SCAN_IN,
    P1_P1_EAX_REG_17__SCAN_IN, P1_P1_EAX_REG_18__SCAN_IN,
    P1_P1_EAX_REG_19__SCAN_IN, P1_P1_EAX_REG_20__SCAN_IN,
    P1_P1_EAX_REG_21__SCAN_IN, P1_P1_EAX_REG_22__SCAN_IN,
    P1_P1_EAX_REG_23__SCAN_IN, P1_P1_EAX_REG_24__SCAN_IN,
    P1_P1_EAX_REG_25__SCAN_IN, P1_P1_EAX_REG_26__SCAN_IN,
    P1_P1_EAX_REG_27__SCAN_IN, P1_P1_EAX_REG_28__SCAN_IN,
    P1_P1_EAX_REG_29__SCAN_IN, P1_P1_EAX_REG_30__SCAN_IN;
  output P1_P1_U2721;
  wire n60029, n67389, n74249, n74250, n74411, n74402, n76063, n60391,
    n71659, n59826, n64666, n64646, n60099, n60746, n64475, n64530, n67227,
    n71298, n61148, n64350, n97978, n64163, n60274, n64744, n67854, n64444,
    n63124, n63069, n70069, n63200, n64095, n60986, n71512, n59789, n61370,
    n64562, n63897, n63999, n59828, n63434, n63632, n61570, n71397, n62965,
    n60408, n59835, n59829, n64574, n59830, n74835, n59911, n63724, n59991,
    n76045, n60623, n60899, n71664, n67268, n67807, n70003, n71404, n63329,
    n63327, n64214, n59923, n60214, n59790, n64008, n63613, n64645, n60503,
    n59791, n60007, n61366, n64635, n63852, n60101, n68769, n60502, n64231,
    n59796, n64787, n70143, n71294, n71187, n59798, n71265, n60844, n70035,
    n63441, n63162, n59799, n60192, n70067, n68788, n63374, n59800, n60094,
    n71365, n64237, n61260, n63458, n71608, n63134, n68854, n68961, n63000,
    n63186, n60133, n60276, n64688, n60389, n60078, n60839, n59805, n64599,
    n60388, n60024, n75900, n64578, n61495, n64579, n59806, n60134, n64263,
    n71669, n60481, n61145, n59813, n59814, n67886, n60117, n61435, n59815,
    n59816, n64504, n63918, n63614, n64543, n60882, n67361, n63331, n64190,
    n64110, n71230, n71372, n61483, n64701, n63863, n61474, n63619, n64022,
    n64614, n59827, n70158, n68945, n62915, n63129, n64497, n62937, n61255,
    n59831, n71696, n63581, n71410, n71402, n63941, n63620, n63478, n63935,
    n59832, n67939, n61410, n70174, n71199, n60937, n63882, n59836, n63504,
    n59837, n67275, n64031, n68802, n60263, n64683, n70160, n63387, n68955,
    n63670, n64362, n59841, n59842, n64136, n71374, n59863, n61443, n67255,
    n67853, n67860, n59846, n63287, n63284, n67751, n64566, n59850, n60077,
    n74790, n74336, n70047, n71575, n74348, n75984, n75987, n74277, n60455,
    n63436, n64297, n60486, n65183, n59854, n71487, n67799, n60093, n61147,
    n64049, n64240, n64238, n64457, n59857, n59858, n63886, n60032, n60880,
    n59859, n59860, n59861, n71213, n61361, n59862, n68806, n59864, n60832,
    n71619, n67296, n59865, n59866, n59867, n59868, n59869, n59870, n68927,
    n60478, n64717, n64409, n63270, n74416, n64758, n76064, n61389, n76182,
    n74846, n74361, n74396, n59892, n59893, n59896, n59961, n59897, n59912,
    n59901, n63483, n63202, n59902, n59903, n59904, n67364, n63282, n59995,
    n64038, n64643, n64748, n67360, n61149, n67776, n60034, n59997, n74739,
    n64157, n64144, n64523, n63656, n63898, n59905, n59906, n59907, n59908,
    n59909, n59910, n74830, n75995, n59994, n70178, n70074, n70028, n74774,
    n61161, n60087, n68875, n60444, n71198, n64307, n60025, n60022, n63912,
    n67331, n64011, n60279, n60185, n64208, n71248, n60863, n64770, n64387,
    n63847, n64452, n74119, n59913, n59914, n63317, n60096, n71589, n71577,
    n64568, n67359, n70148, n64573, n67827, n64281, n68894, n68895, n64659,
    n67358, n63976, n59915, n64652, n74431, n67842, n68882, n70191, n63849,
    n74409, n75949, n68766, n67916, n71597, n71588, n60452, n74220, n60626,
    n71697, n71683, n74749, n71692, n71175, n69996, n74446, n67920, n71390,
    n67197, n74248, n68956, n61319, n60283, n60281, n68782, n64115, n64795,
    n64472, n64463, n60090, n67236, n60103, n60089, n60915, n64460, n61442,
    n60136, n64549, n63924, n70107, n60037, n60233, n70022, n64209, n60928,
    n68891, n63488, n67321, n63837, n67849, n61159, n63226, n64282, n60225,
    n60451, n63390, n60506, n63351, n63337, n60492, n67278, n60264, n60417,
    n63247, n63246, n64817, n60465, n67781, n59976, n64577, n60497, n64065,
    n71483, n59980, n74798, n74730, n59984, n59930, n76054, n76037, n74315,
    n59935, n59936, n59937, n59938, n60500, n76051, n64694, n64697, n64369,
    n59940, n74747, n76213, n61577, n71684, n61491, n60467, n60414, n74754,
    n71691, n71694, n71183, n71172, n71176, n60188, n71478, n69992, n71678,
    n74769, n69991, n60231, n61444, n67940, n71180, n60131, n71403, n67927,
    n61261, n59942, n68765, n74785, n67933, n67937, n68998, n68996, n75941,
    n68997, n67935, n74246, n68993, n74222, n67929, n68980, n68995, n67928,
    n67936, n68974, n67380, n68976, n67382, n61131, n60469, n74254, n74253,
    n67193, n71657, n75933, n60395, n67375, n67367, n74430, n68771, n74437,
    n64332, n70190, n60462, n67371, n76793, n64800, n64508, n64663, n74945,
    n67899, n60209, n64329, n74960, n64661, n68949, n64487, n67219, n73153,
    n64125, n60050, n67216, n67215, n71492, n72804, n67748, n64325, n63939,
    n64116, n64130, n64481, n63792, n70145, n64321, n61322, n61323, n70254,
    n64127, n64336, n64122, n71496, n68789, n60458, n64343, n63933, n75991,
    n67223, n60123, n71210, n64517, n74920, n64112, n64132, n64790, n71358,
    n64533, n63809, n63934, n63585, n70011, n68822, n63584, n64477, n60102,
    n60235, n60191, n63802, n63589, n64531, n60040, n63477, n64133, n74903,
    n61452, n63799, n61455, n61090, n67228, n64775, n60513, n63570, n63928,
    n74902, n71221, n64105, n63952, n60097, n60091, n71349, n76137, n61367,
    n63946, n64166, n60086, n64165, n64182, n71343, n60083, n63303, n60400,
    n60403, n71603, n64761, n63834, n63831, n60402, n60459, n63587, n64180,
    n64759, n60232, n74269, n64633, n63685, n70119, n61002, n71327, n60033,
    n60271, n63829, n60270, n60212, n74885, n70124, n63681, n68926, n63554,
    n71237, n63552, n64100, n63666, n63993, n63591, n60629, n60058, n64626,
    n64450, n60927, n68918, n60213, n68917, n68919, n74880, n63470, n63465,
    n64088, n60376, n64312, n64235, n70097, n71313, n60183, n60016, n70112,
    n63219, n74797, n64446, n60018, n63460, n61019, n60382, n63669, n63968,
    n60224, n60043, n63454, n60017, n60210, n64301, n63216, n71559, n60277,
    n74865, n60044, n63222, n61141, n63449, n60211, n60045, n63448, n63450,
    n64679, n71289, n63139, n74863, n61372, n60404, n63445, n63358, n63117,
    n74332, n67855, n71546, n63439, n63438, n63111, n60218, n60226, n61357,
    n70087, n63651, n60895, n71295, n64288, n60446, n63368, n67309, n70077,
    n64063, n59954, n63106, n63355, n63433, n63223, n61130, n63365, n60216,
    n63495, n63431, n67845, n63019, n68837, n60182, n64608, n63386, n70080,
    n59955, n64010, n63055, n67837, n68877, n68873, n60115, n60509, n71507,
    n74834, n63858, n60636, n61359, n63635, n60840, n60638, n60510, n64054,
    n70066, n60637, n63642, n64407, n70068, n63862, n67289, n71274, n70062,
    n63424, n63631, n63338, n63347, n67830, n62913, n62970, n67284, n67283,
    n61249, n67831, n67822, n60924, n63277, n62966, n62984, n67261, n67282,
    n63093, n60175, n62918, n62964, n62911, n70052, n63268, n64273, n62979,
    n62981, n63255, n61362, n60457, n67824, n63521, n63343, n60877, n67256,
    n74799, n60201, n67801, n67808, n60200, n64699, n62994, n71520, n63340,
    n63160, n63167, n63263, n62917, n60202, n63624, n62995, n64587, n60454,
    n60949, n62893, n62924, n63076, n61320, n62920, n63039, n97991, n60448,
    n67812, n60039, n60577, n60464, n63157, n64581, n64712, n60084, n61496,
    n60082, n60051, n60450, n60631, n60265, n63841, n60490, n64632, n64196,
    n97185, n71197, n98007, n70176, n70096, n67752, n63152, n60221, n97988,
    n71212, n97987, n98011, n59967, n97999, n68928, n59969, n98008, n98002,
    n71203, n97982, n67880, n60630, n70043, n59970, n60449, n67780, n59972,
    n74360, n64249, n64710, n67272, n60262, n60498, n63860, n59974, n76000,
    n74367, n60184, n60047, n76067, n64376, n60483, n65136, n64390, n65129,
    n97866, n64808, n61527, n98052, n64827, n61526, n61500, n67287, n74806,
    n64709, n60723, n63874, n76012, n74881, n60375, n71521, n68848, n64706,
    n64832, n100056, n71192, n59986, n64824, n59988, n64375, n60517,
    n61062, n60179, n60634, n60501, n68904, n63412, n64250, n62986, n67777,
    n59992, n71171, n64572, n74763, n60721, n100090, n100136, n63855,
    n100087, n99991, n65089, n100072, n61063, n60715, n62928, n60178,
    n60493, n60904, n71188, n64607, n59993, n60079, n67756, n59996, n67332,
    n67329, n64742, n59998, n64613, n64612, n59999, n71394, n70023, n67898,
    n71205, n68965, n67312, n64669, n64527, n60006, n68774, n63406, n60411,
    n60505, n60008, n64424, n63596, n60009, n60507, n64414, n64247, n64252,
    n64251, n64244, n60013, n64032, n60642, n60484, n60015, n61150, n70098,
    n60019, n67266, n60020, n75002, n64721, n60021, n74761, n74759, n60023,
    n60026, n71479, n60487, n60027, n60028, n60627, n60624, n60639, n68779,
    n64089, n68768, n74831, n60035, n74288, n74314, n60038, n61569, n60508,
    n63349, n60516, n60892, n64314, n64522, n64348, n68952, n60041, n60722,
    n64512, n60042, n63910, n64662, n60046, n71240, n63097, n60048, n63121,
    n60049, n60261, n67365, n63798, n60644, n63092, n70071, n60056, n60336,
    n68939, n64565, n60132, n67800, n60399, n67743, n60057, n60220, n61089,
    n61318, n60255, n61095, n61487, n64354, n64451, n60409, n61479, n71200,
    n61390, n63845, n68773, n70192, n60080, n67735, n71364, n76218, n64593,
    n60065, n64590, n61411, n67744, n63415, n63601, n67762, n68938, n60073,
    n67760, n70016, n74733, n67319, n60076, n61164, n64682, n68798, n64650,
    n67738, n60081, n64768, n60085, n60098, n67888, n64774, n60088, n64783,
    n68957, n67907, n60092, n64640, n68968, n71387, n61143, n63951, n63807,
    n63691, n63797, n60095, n63636, n67891, n64335, n60100, n64347, n64532,
    n63345, n60114, n63644, n60116, n67377, n64342, n60252, n64384, n64389,
    n64629, n60135, n64772, n60230, n67324, n67328, n64364, n71481, n67875,
    n64401, n64400, n60173, n60174, n67881, n67883, n60176, n63618, n63625,
    n60177, n60936, n60180, n64068, n60181, n68921, n64513, n64514, n60189,
    n60186, n71412, n60187, n74206, n60190, n70020, n61365, n63257, n63258,
    n64367, n70102, n70095, n60198, n60199, n60208, n64211, n60215, n61383,
    n60217, n60219, n60222, n64796, n60223, n67205, n63972, n60763, n60227,
    n60228, n63627, n60229, n71672, n63833, n60234, n61135, n63836, n63647,
    n60249, n64405, n60657, n61489, n60253, n71190, n71405, n60258, n60259,
    n67902, n67897, n60260, n64242, n68954, n60266, n60267, n60268, n64548,
    n60269, n60272, n64631, n60273, n64455, n60278, n60275, n63633, n60282,
    n60280, n71648, n71650, n71655, n60328, n71363, n74434, n60334, n68821,
    n60335, n67238, n67224, n64792, n60337, n60519, n63077, n62879, n71251,
    n62883, n64440, n64449, n71500, n60995, n60377, n64283, n60379, n71268,
    n60378, n64275, n60380, n71310, n60381, n74436, n71384, n60383, n70049,
    n60384, n60385, n60386, n60387, n70122, n71473, n71392, n74452, n64678,
    n67333, n64627, n60390, n60393, n60392, n60394, n60396, n60401, n60405,
    n63630, n63423, n60410, n60413, n76210, n60415, n60859, n60889, n74210,
    n60441, n60442, n60443, n60445, n60447, n67784, n68851, n64417, n74735,
    n60453, n77917, n60456, n62919, n63487, n63112, n63791, n63562, n63772,
    n64333, n60461, n60463, n60466, n60628, n60471, n60470, n64391, n60480,
    n60479, n60482, n74782, n60485, n61446, n75899, n67327, n67865, n60488,
    n60489, n70128, n60491, n70125, n60494, n60496, n74804, n74812, n60499,
    n67915, n68767, n64647, n60504, n61572, n63350, n64134, n60511, n60512,
    n60514, n60515, n60518, n71182, n60534, n71676, n74216, n60625, n71234,
    n68846, n60632, n60633, n60635, n71202, n75007, n60641, n75005, n60640,
    n74226, n74770, n60643, n76206, n60647, n60648, n67755, n60650, n67353,
    n67347, n60651, n70001, n60652, n70002, n71389, n70196, n60656, n63316,
    n68841, n64412, n64408, n64406, n60672, n60673, n60716, n67325, n60718,
    n64232, n60950, n60720, n67866, n63353, n64019, n63156, n74822, n71381,
    n61412, n61137, n63592, n70173, n68899, n64270, n60908, n64303, n74760,
    n63672, n68947, n74466, n61075, n64745, n64365, n61061, n64260, n67295,
    n64075, n61387, n61393, n61394, n67847, n64557, n67320, n61038, n74295,
    n67343, n63144, n60856, n74326, n64183, n74346, n64537, n63363, n63292,
    n64177, n71616, n61009, n61007, n70186, n61344, n71647, n71646, n63676,
    n69997, n61350, n64337, n64496, n64318, n76211, n61436, n64033, n60893,
    n64386, n61259, n64693, n67791, n67273, n60948, n61247, n67292, n63864,
    n60900, n63407, n63878, n63323, n63321, n64051, n60858, n67310, n64359,
    n64426, n67833, n61386, n71269, n61023, n71545, n62942, n67339, n61243,
    n61165, n71526, n71561, n60988, n60989, n60990, n61470, n64753, n64755,
    n63432, n63429, n70135, n61385, n60841, n61018, n64204, n61485, n61490,
    n64200, n63279, n74824, n61449, n61450, n74328, n62888, n63180, n61454,
    n71600, n74368, n63657, n63437, n63447, n61017, n74255, n61021, n63662,
    n63832, n63373, n60875, n60854, n60994, n71633, n74260, n61020, n74948,
    n61463, n61465, n68948, n60945, n61477, n68958, n74445, n68982, n64484,
    n61126, n61127, n64128, n61124, n63588, n63473, n63474, n61346, n61347,
    n61345, n76076, n64109, n74738, n71186, n68992, n64328, n64117, n61445,
    n60881, n64576, n64361, n63888, n63877, n64592, n64395, n64396, n60947,
    n61484, n61250, n67250, n61360, n63148, n63150, n67841, n60940, n64677,
    n64081, n64059, n64052, n63623, n71533, n68843, n61262, n67848, n64432,
    n64224, n63980, n63417, n63163, n63158, n62997, n60852, n70082, n60939,
    n67330, n64437, n64304, n67862, n68915, n61263, n71288, n60991, n74330,
    n61022, n64628, n64447, n63981, n63905, n61369, n63276, n74284, n74300,
    n71315, n62922, n67233, n67350, n64756, n64754, n63649, n63174, n60847,
    n70149, n60998, n74343, n63603, n64546, n60968, n64206, n61001, n61003,
    n68787, n63923, n63357, n63014, n63006, n60996, n71361, n61458, n74376,
    n67890, n64156, n74939, n70187, n62909, n64671, n61480, n64316, n63956,
    n61133, n61343, n63022, n71660, n71658, n74976, n74395, n71388, n63026,
    n64511, n60853, n74447, n64506, n61138, n74221, n61476, n61373, n63574,
    n74219, n61241, n76038, n67913, n61256, n61348, n61439, n76061, n63575,
    n63706, n64837, n64835, n76046, n76043, n61437, n63931, n75033, n97746,
    n67923, n60873, n68989, n78645, n99992, n96865, n76802, n71174, n99201,
    n97648, n62435, n76224, n98061, n97645, n60728, n75006, n60862, n60729,
    n60730, n60731, n61012, n60734, n60736, n74820, n74882, n60740, n61251,
    n60747, n60878, n64056, n61004, n60750, n60752, n60759, n60761, n63885,
    n60762, n61162, n60764, n75994, n64266, n60926, n61395, n60768, n60769,
    n60773, n60774, n60776, n60778, n63296, n97204, n60788, n60790, n60791,
    n60792, n60796, n60799, n60802, n61246, n64536, n61160, n64456, n61146,
    n61460, n60803, n60805, n60806, n60808, n60810, n60811, n60812, n60814,
    n60933, n60816, n60819, n61364, n61142, n67884, n61132, n68803, n64397,
    n61163, n61144, n63638, n61078, n60834, n64147, n60835, n60836, n63066,
    n68804, n68801, n60838, n64731, n61462, n71572, n74261, n60842, n74793,
    n61151, n64596, n71264, n70144, n70105, n60846, n63165, n63281, n60848,
    n61349, n60851, n60855, n63143, n60857, n61079, n61492, n64352, n67225,
    n63828, n68878, n61094, n61082, n60876, n60860, n60861, n64431, n68970,
    n60865, n71325, n74391, n63970, n60871, n68797, n60872, n70195, n63199,
    n63827, n63810, n60874, n63950, n63140, n64588, n71681, n71635, n75000,
    n68815, n64402, n60879, n68824, n67761, n64044, n64776, n68884, n60938,
    n68819, n68813, n64366, n74208, n64801, n64415, n60890, n68775, n67911,
    n64024, n64028, n60925, n64269, n64296, n60894, n64292, n64425, n64295,
    n64428, n61104, n64586, n64618, n64445, n64624, n64767, n67207, n71391,
    n64239, n64018, n63917, n69998, n61125, n68978, n60929, n60931, n60932,
    n60934, n61475, n64442, n60935, n64057, n67867, n70118, n67306, n68836,
    n60943, n60946, n60941, n60942, n60944, n67241, n67354, n60984, n60985,
    n71516, n71256, n60987, n60992, n60993, n74407, n60997, n74832, n60999,
    n61000, n74265, n61008, n61005, n61006, n61014, n61016, n61010, n61011,
    n61013, n61015, n74380, n71524, n71547, n71506, n74456, n71401, n61036,
    n67771, n61039, n64603, n61065, n64752, n64743, n61080, n61081, n70193,
    n61371, n61093, n67213, n67212, n61441, n64198, n64636, n68791, n68790,
    n67889, n61128, n61129, n67921, n68984, n61134, n64797, n61136, n63594,
    n63677, n61139, n67859, n61140, n61245, n63334, n64459, n67829, n61152,
    n61158, n64005, n63903, n64399, n61166, n74217, n74209, n74743, n61242,
    n61244, n64735, n61248, n64357, n61252, n61253, n61254, n64026, n61258,
    n71287, n71582, n71675, n61440, n68888, n70108, n68893, n64720, n64695,
    n71371, n64616, n64737, n61321, n61324, n63668, n63313, n61358, n64556,
    n64558, n61363, n63404, n68972, n61368, n63915, n64289, n68777, n61384,
    n61388, n61391, n61392, n71474, n67753, n67244, n67368, n64657, n61438,
    n63803, n64478, n61447, n63899, n74787, n75001, n61448, n74915, n74932,
    n61451, n61456, n61453, n61461, n61457, n61459, n74404, n61464, n61471,
    n74841, n61472, n64766, n61473, n64630, n61478, n68964, n64791, n67220,
    n61481, n61482, n74448, n71668, n61486, n61488, n61493, n61494, n64093,
    n64580, n63902, n74240, n67240, n63611, n64718, n64225, n64218, n67362,
    n63896, n61511, n61519, n61522, n71345, n68776, n61528, n61534, n61535,
    n68816, n64015, n61549, n61551, n64528, n61553, n97723, n61554, n61555,
    n76028, n62954, n61571, n61573, n63796, n61574, n61575, n64261, n68856,
    n64380, n64255, n64589, n63607, n68852, n64074, n71279, n67840, n68880,
    n71293, n64061, n64221, n63402, n74353, n64443, n67872, n68935, n63653,
    n67878, n63907, n70170, n63444, n68944, n63663, n71501, n68781, n64473,
    n64173, n63466, n76081, n63671, n63023, n63468, n63308, n63221, n74245,
    n74982, n63382, n63808, n76056, n68778, n64642, n74788, n74771, n63929,
    n64491, n71398, n74780, n68979, n74930, n71181, n67379, n64651, n75055,
    n97761, n97225, n63775, n71469, n99178, n100130, n70255, n62410,
    n99199, n97747, n74470, n71419, n71693, n75022, n99221, n99213,
    n100048, n97895, n70278, n96896, n99179, n97620, n97930, n100479,
    n96895, n97928, n99180, n100164, n62434, n96899, n97556, n97636,
    n97929, n97971, n100044, n62412, n62408, n62407, n62409, n62411,
    n62428, n62414, n62413, n62418, n62416, n62415, n62417, n62426, n62420,
    n62419, n62424, n62422, n62421, n62423, n62425, n62427, n62433, n62430,
    n62429, n62431, n62432, n74276, n62926, n62880, n64259, n62881, n62921,
    n62882, n62884, n62885, n62897, n62886, n62887, n62892, n62890, n62889,
    n62914, n62891, n62907, n62895, n62894, n62896, n63029, n62898, n63040,
    n62901, n62899, n62900, n63031, n62903, n62902, n62905, n63028, n63027,
    n62904, n62906, n62908, n62910, n63024, n62912, n62939, n62916, n62923,
    n62957, n62944, n62925, n62932, n62927, n62948, n62989, n62930, n62929,
    n62931, n62945, n62956, n62960, n62961, n62967, n62933, n62934, n62935,
    n62938, n63057, n62936, n62941, n62940, n62976, n63005, n62974, n63064,
    n62943, n62947, n62946, n62949, n62952, n62950, n62951, n62953, n62996,
    n62998, n62955, n62982, n62980, n62959, n62958, n63181, n62963, n62962,
    n62969, n62968, n62973, n62971, n62972, n63179, n63188, n63178, n63062,
    n62978, n62975, n62977, n63224, n62985, n62983, n63175, n63166, n62987,
    n62988, n62993, n62992, n62990, n62991, n63164, n62999, n63142, n63001,
    n63002, n63003, n63004, n63020, n63395, n63011, n63008, n63007, n63018,
    n63182, n63190, n63010, n63009, n63016, n63012, n63013, n63015, n63017,
    n63021, n63227, n63197, n63204, n63025, n63053, n63049, n63030, n63045,
    n63032, n63080, n63034, n63033, n63035, n63037, n63036, n63038, n63074,
    n63043, n63041, n63042, n63044, n63090, n63089, n63047, n63046, n63048,
    n63099, n63098, n63051, n63050, n63052, n63104, n63103, n63054, n63058,
    n63059, n63071, n63072, n63061, n63060, n63063, n63067, n63065, n63070,
    n63203, n63068, n63482, n63073, n63075, n63087, n63078, n63079, n63083,
    n63082, n63511, n63081, n63502, n63085, n63084, n63086, n63516, n63517,
    n63088, n63091, n63096, n63094, n63095, n63497, n63496, n63101, n63100,
    n63490, n63491, n63102, n63108, n63107, n63489, n63105, n63110, n63109,
    n63486, n63114, n63113, n63481, n63115, n63116, n63122, n63119, n63118,
    n63120, n63123, n63548, n63549, n63553, n63125, n63127, n63128, n63126,
    n63130, n63212, n63136, n63131, n63838, n63132, n63843, n63133, n63135,
    n63137, n63138, n63141, n63271, n63145, n63274, n63172, n63146, n63147,
    n63149, n63151, n63241, n63244, n63243, n63153, n63154, n63252, n63266,
    n63155, n63161, n63159, n63251, n63265, n63261, n63170, n63169, n63168,
    n63260, n63273, n63171, n63285, n63173, n63289, n63177, n63288, n63176,
    n63233, n63184, n63189, n63183, n63185, n63195, n63187, n63193, n63191,
    n63192, n63194, n63232, n63231, n63196, n63230, n63198, n63201, n63209,
    n63207, n63205, n63206, n63208, n63217, n63215, n63211, n63214, n63210,
    n63479, n63213, n63218, n63307, n63220, n63306, n63225, n63228, n63235,
    n63234, n63361, n63238, n63236, n63237, n63239, n63240, n63328, n63242,
    n63245, n63333, n63339, n63341, n63248, n63249, n63250, n63253, n63262,
    n63254, n63256, n63346, n63348, n63259, n63264, n63267, n63269, n63272,
    n63275, n63278, n63280, n63312, n63310, n63299, n63283, n63286, n63295,
    n63293, n63291, n63290, n63294, n63356, n63362, n63366, n63297, n63298,
    n63360, n63300, n63372, n63305, n63301, n63379, n63563, n63302, n63572,
    n63304, n63378, n63309, n63472, n63311, n63315, n63314, n63320, n63318,
    n63319, n63414, n63325, n63322, n63326, n63324, n63330, n63332, n63336,
    n63335, n63427, n63426, n63342, n63393, n63344, n63389, n63352, n63440,
    n63442, n63354, n63359, n63369, n63364, n63367, n63370, n63451, n63371,
    n63459, n63462, n63376, n63461, n63375, n63679, n63469, n63377, n63571,
    n63385, n63565, n63383, n63381, n63380, n63384, n63388, n63392, n63391,
    n63652, n63394, n63397, n63396, n63401, n63399, n63398, n63400, n63403,
    n63405, n63641, n63430, n63408, n63616, n63410, n63867, n63409, n63411,
    n63413, n63600, n63416, n63615, n63422, n63418, n63419, n63420, n63421,
    n63634, n63425, n63428, n63597, n63435, n63908, n63443, n63658, n63446,
    n63455, n63453, n63452, n63667, n63456, n63457, n63464, n63463, n63467,
    n63590, n63682, n63471, n63475, n63476, n63582, n63693, n63480, n63560,
    n63558, n63700, n63485, n63484, n63544, n63541, n63540, n63709, n63537,
    n63493, n63492, n63494, n63531, n63527, n63498, n63501, n63499, n63500,
    n63503, n63510, n63505, n63506, n63717, n72811, n63723, n63716, n63509,
    n63507, n63508, n63512, n63513, n63732, n63731, n63515, n63514, n63523,
    n63522, n63715, n63519, n63518, n63520, n63714, n63525, n63524, n63526,
    n63742, n63741, n63529, n63528, n63532, n63713, n63712, n63530, n63535,
    n63533, n63534, n63536, n63755, n63754, n63539, n63538, n63710, n63543,
    n63542, n63545, n63708, n63707, n63547, n63546, n63555, n63551, n63550,
    n63702, n63703, n63557, n63556, n63559, n63561, n63568, n63567, n63699,
    n63564, n63566, n63698, n63569, n63579, n63573, n63577, n63576, n63578,
    n63697, n63696, n63580, n63694, n63583, n63692, n63593, n63595, n63599,
    n63906, n63598, n63602, n63605, n76062, n63604, n63606, n63608, n64036,
    n63871, n63873, n63609, n63883, n63610, n63612, n63621, n63617, n63890,
    n63893, n63622, n63626, n63628, n63629, n63891, n63848, n63637, n63996,
    n63835, n63639, n63640, n63643, n63645, n63646, n63648, n63650, n63655,
    n63654, n63974, n63904, n63914, n63916, n63661, n63660, n63659, n63664,
    n63830, n63665, n63673, n63826, n63674, n63675, n63678, n63688, n63680,
    n63686, n63684, n63683, n63687, n63943, n63800, n63689, n63945, n63690,
    n63932, n63790, n63695, n63787, n63785, n97644, n63782, n63781, n75021,
    n63778, n63777, n74469, n63701, n63773, n71699, n63705, n63704, n63769,
    n63768, n71420, n63765, n63764, n70199, n63711, n63761, n63760, n69006,
    n63749, n63750, n67465, n63748, n63738, n63737, n78651, n63718, n63719,
    n63730, n76798, n63720, n73159, n63722, n63721, n73158, n63728, n63726,
    n63725, n63727, n76797, n63729, n63734, n63733, n74125, n74124, n63736,
    n63735, n78650, n63740, n63739, n63744, n63743, n65162, n65161, n63746,
    n63745, n67466, n63747, n63753, n63751, n63752, n63757, n63756, n67984,
    n67985, n63759, n63758, n69007, n63763, n63762, n70200, n63767, n63766,
    n63771, n63770, n71700, n63776, n63774, n63780, n63779, n63784, n63783,
    n97643, n63789, n63786, n63788, n63938, n63960, n63793, n63794, n63795,
    n63805, n63801, n63804, n63806, n63942, n63811, n63944, n63948, n63812,
    n63825, n63814, n63813, n63816, n63815, n63823, n63817, n63821, n63818,
    n63819, n63820, n63822, n63824, n64142, n63998, n63840, n63839, n63842,
    n63844, n63846, n63982, n63850, n63851, n64007, n63853, n63854, n63856,
    n63857, n63859, n63861, n63865, n64041, n63866, n63869, n63868, n64037,
    n64267, n64016, n63870, n63872, n63876, n63875, n63880, n63879, n63881,
    n63889, n63884, n63887, n64066, n63894, n63892, n63895, n64220, n64006,
    n63900, n63901, n64090, n63909, n63911, n64092, n64091, n64094, n63913,
    n64099, n63920, n63919, n63922, n63921, n63925, n64168, n64104, n63957,
    n63926, n63947, n63927, n64108, n63930, n64120, n64119, n63937, n63936,
    n64118, n72805, n63940, n64124, n63949, n63953, n64154, n63954, n63955,
    n63964, n63958, n63959, n63962, n64146, n63965, n63961, n63963, n63967,
    n64137, n63966, n63969, n63971, n63973, n63975, n63977, n63979, n64201,
    n63986, n63994, n63985, n63983, n63984, n63988, n63987, n63991, n63989,
    n63990, n63992, n63995, n64002, n63997, n64000, n64001, n64003, n64004,
    n64087, n64309, n64073, n64009, n64014, n64012, n64013, n64236, n64062,
    n64017, n64271, n64027, n64029, n64020, n64021, n64023, n64025, n64030,
    n64262, n64034, n64035, n64045, n64040, n64039, n64042, n64043, n64241,
    n64046, n64047, n64048, n64050, n64286, n64284, n64060, n64053, n64055,
    n64058, n64083, n64072, n64064, n64070, n64067, n64069, n64071, n64080,
    n64078, n64076, n64077, n64079, n64082, n64222, n64310, n64084, n64085,
    n64086, n64313, n64199, n64097, n64096, n64185, n64098, n64187, n64102,
    n64186, n64101, n64171, n64103, n64106, n64107, n64139, n64150, n64164,
    n64131, n64114, n64111, n64113, n64319, n64123, n64323, n64121, n73154,
    n64126, n64129, n64135, n64141, n64138, n64140, n64153, n64143, n64145,
    n64149, n64148, n64151, n64152, n64162, n64155, n64160, n64158, n64159,
    n64161, n64175, n64170, n64167, n64174, n64169, n64172, n64179, n64176,
    n64178, n64525, n64181, n64184, n64188, n64189, n64192, n64191, n64195,
    n64193, n64194, n64197, n64207, n64203, n64202, n64205, n64213, n64210,
    n64212, n64216, n64215, n64353, n64217, n64435, n64230, n64219, n64229,
    n64223, n64306, n64436, n64227, n64226, n64228, n64233, n64234, n64305,
    n64419, n64243, n64403, n64567, n64246, n64392, n64245, n64248, n64253,
    n64254, n64256, n64257, n64258, n64583, n64381, n64264, n64265, n64268,
    n64272, n64276, n64274, n64277, n64410, n64278, n64418, n64280, n64279,
    n64422, n64285, n64287, n64427, n64291, n64302, n64290, n64293, n64300,
    n64294, n64298, n64299, n64308, n64311, n64355, n64349, n64315, n64339,
    n64334, n64338, n64317, n64492, n64327, n64320, n64322, n64324, n64326,
    n64490, n64489, n64330, n64331, n64495, n64340, n64341, n64470, n64526,
    n64346, n64777, n64344, n64345, n64461, n64539, n64351, n64356, n64358,
    n64622, n64617, n64551, n64360, n64434, n64363, n64584, n64368, n64372,
    n64370, n64371, n64374, n64373, n64379, n64377, n64378, n64382, n64383,
    n64385, n64388, n64393, n64394, n64398, n64600, n64404, n64601, n64413,
    n64411, n64416, n64561, n64420, n64421, n64423, n64429, n64555, n64430,
    n64620, n64433, n64438, n64439, n64441, n64448, n64453, n64454, n64458,
    n64469, n64462, n64466, n64464, n64465, n64467, n64468, n64471, n64474,
    n64476, n64479, n64509, n64515, n64480, n64644, n64482, n64483, n64486,
    n64499, n64485, n64488, n64655, n64653, n64494, n64493, n74120, n64498,
    n64505, n67369, n64502, n64500, n64501, n64503, n64507, n64510, n64518,
    n64516, n64519, n67214, n64520, n64521, n64524, n64534, n64529, n64667,
    n64535, n64538, n64541, n64540, n64542, n64547, n64545, n64544, n64673,
    n64769, n64621, n64550, n64553, n64552, n64554, n64559, n64739, n64560,
    n64563, n64564, n64569, n64570, n64571, n67274, n64575, n64582, n64585,
    n64698, n67291, n67293, n64725, n64591, n64594, n64595, n64598, n64597,
    n64729, n64602, n64730, n64605, n64604, n64733, n64606, n64684, n64685,
    n64609, n64610, n64611, n64615, n64738, n64619, n64625, n64623, n64634,
    n64757, n67229, n64637, n64638, n64674, n64639, n64670, n64641, n64648,
    n64649, n64654, n64656, n64658, n67387, n64660, n67195, n64665, n64664,
    n64803, n64668, n64672, n67741, n64794, n64675, n64676, n64680, n64681,
    n64736, n67323, n64686, n64687, n67318, n64692, n64689, n64690, n64691,
    n67251, n64723, n64696, n64700, n64703, n64702, n64705, n64704, n64707,
    n64708, n64711, n67276, n67279, n64714, n64713, n64716, n67262, n64715,
    n64719, n67257, n64722, n67299, n67248, n64724, n64727, n64726, n64728,
    n67247, n67313, n64734, n64732, n64741, n64740, n67335, n67334, n67338,
    n67341, n64746, n64747, n67342, n64749, n64751, n64750, n67243, n67239,
    n67242, n67348, n64763, n64760, n64762, n67351, n64764, n67346, n64765,
    n64773, n64771, n67226, n64778, n64784, n64781, n64779, n64780, n64782,
    n64788, n64786, n64789, n67221, n64793, n64798, n67208, n64799, n67203,
    n67374, n64802, n67198, n64804, n67192, n67194, n64805, n67384, n76044,
    n67390, n67381, n100184, n100434, n96193, n97203, n64810, n97743,
    n64809, n64814, n64812, n97998, n64811, n64813, n64823, n64816, n97754,
    n64815, n64821, n100108, n100123, n64819, n64818, n64820, n64822,
    n64845, n64826, n64825, n64831, n97303, n64829, n64828, n64830, n64843,
    n64834, n64836, n75052, n64833, n64841, n64839, n64838, n64840, n64842,
    n64844, n64847, n64846, n64851, n64849, n64848, n64850, n64859, n64853,
    n64852, n64857, n64855, n64854, n64856, n64858, n64875, n64861, n64860,
    n64865, n64863, n64862, n64864, n64873, n64867, n64866, n64871, n64869,
    n64868, n64870, n64872, n64874, n64877, n64876, n64881, n64879, n64878,
    n64880, n64889, n64883, n64882, n64887, n64885, n64884, n64886, n64888,
    n64905, n64891, n64890, n64895, n64893, n64892, n64894, n64903, n64897,
    n64896, n64901, n64899, n64898, n64900, n64902, n64904, n64907, n64906,
    n64911, n64909, n64908, n64910, n64935, n64913, n64912, n64915, n64914,
    n64917, n64916, n64933, n64919, n64918, n64923, n64921, n64920, n64922,
    n64931, n64925, n64924, n64929, n64927, n64926, n64928, n64930, n64932,
    n64934, n65062, n64936, n64967, n64938, n64937, n64942, n64940, n97979,
    n64939, n64941, n64950, n64944, n64943, n64948, n64946, n64945, n64947,
    n64949, n64966, n64952, n64951, n64956, n64954, n64953, n64955, n64964,
    n64958, n64957, n64962, n64960, n64959, n64961, n64963, n64965, n96898,
    n64999, n64969, n64968, n64973, n64971, n64970, n64972, n64981, n64975,
    n64974, n64979, n64977, n64976, n64978, n64980, n64997, n64983, n64982,
    n64987, n64985, n64984, n64986, n64995, n64989, n64988, n64993, n64991,
    n64990, n64992, n64994, n64996, n65071, n64998, n65066, n65001, n65000,
    n65005, n65003, n65002, n65004, n65013, n65007, n65006, n65011, n65009,
    n65008, n65010, n65012, n65029, n65015, n65014, n65019, n65017, n65016,
    n65018, n65027, n65021, n65020, n65025, n65023, n65022, n65024, n65026,
    n65028, n98214, n99186, n65031, n65030, n65035, n65033, n65032, n65034,
    n65043, n65037, n65036, n65041, n65039, n65038, n65040, n65042, n65059,
    n65045, n65044, n65049, n65047, n65046, n65048, n65057, n65051, n65050,
    n65055, n65053, n65052, n65054, n65056, n65058, n65060, n65061, n65120,
    n65126, n99191, n65064, n65063, n65065, n65079, n100065, n97651,
    n98071, n100471, n99197, n65085, n65067, n65068, n65069, n65070,
    n65077, n65122, n65074, n65072, n65073, n65075, n65076, n65078, n96897,
    n99214, n65080, n100066, n100481, n96146, n65081, n65083, n65082,
    n96131, n100107, n65088, n65084, n99194, n65086, n96132, n96893,
    n65087, n98211, n65111, n100023, n65092, n65103, n65090, n65091,
    n65093, n65094, n65113, n65100, n100141, n65096, n65095, n65098,
    n65105, n65097, n65102, n65099, n65106, n65101, n65116, n96143, n65112,
    n65104, n65110, n65107, n65109, n65108, n65118, n65124, n100076,
    n96141, n65115, n65114, n65117, n65119, n100046, n65121, n99188,
    n99216, n96892, n65123, n100085, n65125, n71418, n97564, n98034,
    n98037, n97591, n97630, n97604, n98337, n98326, n98291, n65168, n97846,
    n65170, n65169, n97808, n97730, n65171, n97708, n97698, n98362, n98357,
    n97655, n97621, n65173, n65172, n97605, n65174, n65175, n97595, n97555,
    n71742, n98024, n67201, n67196, n67199, n67200, n68985, n68983, n67202,
    n67914, n67918, n67204, n67366, n67206, n67210, n67209, n67211, n67217,
    n67218, n67222, n67747, n67234, n67231, n67230, n67232, n67235, n67237,
    n67750, n67246, n67245, n68799, n67345, n67249, n67253, n67252, n67254,
    n67844, n67307, n67259, n67258, n67260, n67263, n67264, n75996, n67270,
    n67265, n67267, n68849, n68857, n68858, n67269, n67814, n68845, n67271,
    n67805, n67813, n67823, n67832, n67277, n67280, n67281, n67836, n67304,
    n67286, n67285, n67288, n67290, n67302, n67294, n67298, n67297, n67300,
    n67301, n67303, n67305, n67308, n67316, n67311, n67314, n67315, n67852,
    n67317, n67322, n67861, n67773, n67864, n67326, n67759, n67770, n67337,
    n67336, n67340, n67344, n67349, n67357, n67352, n67355, n67356, n67363,
    n68959, n67373, n67370, n67372, n67376, n67378, n76055, n67930, n67383,
    n67385, n67386, n67388, n67391, n67397, n67396, n67401, n67399, n67398,
    n67400, n67409, n67403, n67402, n67407, n67405, n67404, n67406, n67408,
    n67425, n67411, n67410, n67415, n67413, n67412, n67414, n67423, n67417,
    n67416, n67421, n67419, n67418, n67420, n67422, n67424, n67943, n67427,
    n67426, n67431, n67429, n67428, n67430, n67439, n67433, n67432, n67437,
    n67435, n67434, n67436, n67438, n67455, n67441, n67440, n67445, n67443,
    n67442, n67444, n67453, n67447, n67446, n67451, n67449, n67448, n67450,
    n67452, n67454, n67942, n67732, n67734, n68994, n67733, n67740, n67736,
    n67737, n67739, n67742, n67746, n67745, n67749, n68950, n68793, n67754,
    n67757, n68936, n67758, n67765, n67763, n67764, n67769, n67767, n67768,
    n67766, n68825, n68827, n67772, n67774, n67775, n67874, n76032, n67782,
    n67778, n67779, n67783, n67785, n67786, n67787, n67793, n67788, n67789,
    n67794, n67790, n67792, n67798, n67795, n67796, n67797, n68863, n67802,
    n67803, n68868, n67804, n67806, n67810, n67809, n67819, n67811, n67817,
    n67815, n67816, n67818, n68867, n67821, n67820, n68871, n68876, n67826,
    n67825, n67828, n67834, n67835, n67838, n68881, n67839, n67843, n67846,
    n68886, n68889, n67851, n67850, n67858, n67856, n67857, n68892, n67863,
    n70110, n70113, n68920, n67873, n67871, n67869, n67868, n67870, n68826,
    n68810, n68809, n68807, n67876, n67877, n67879, n67885, n67882, n67887,
    n67892, n67894, n67893, n68780, n68783, n67895, n67910, n67901, n67896,
    n67904, n67900, n67909, n67903, n67905, n67906, n67908, n67912, n68973,
    n68975, n67922, n67917, n67919, n67924, n67926, n67925, n67934, n67932,
    n67931, n67938, n69047, n67945, n67944, n67949, n67947, n67946, n67948,
    n67973, n67951, n67950, n67953, n67952, n67955, n67954, n67971, n67957,
    n67956, n67961, n67959, n67958, n67960, n67969, n67963, n67962, n67967,
    n67965, n67964, n67966, n67968, n67970, n67972, n69046, n68770, n68772,
    n68784, n70000, n70179, n70188, n68785, n68786, n68792, n68795, n68794,
    n68796, n70182, n70005, n70180, n68800, n68805, n68808, n68811, n68812,
    n68814, n68817, n68818, n70165, n70164, n68820, n68946, n68823, n70146,
    n68828, n68829, n68830, n68833, n68831, n68832, n68834, n68835, n76007,
    n68839, n68840, n70038, n68842, n68844, n68847, n70053, n70054, n70033,
    n68850, n68853, n70057, n70060, n68855, n68861, n68859, n68860, n68862,
    n70059, n68865, n68864, n68866, n68869, n68870, n68872, n70029, n68874,
    n70075, n70089, n68879, n68885, n68883, n70099, n68887, n68890, n68898,
    n68896, n68897, n68900, n68902, n68901, n68903, n68906, n68905, n68908,
    n68907, n68914, n68909, n68912, n68910, n68911, n68913, n68916, n68923,
    n68922, n70129, n70138, n68924, n68925, n68930, n68929, n68931, n68934,
    n70010, n70013, n68932, n68933, n68943, n68937, n68942, n68940, n68941,
    n70166, n70007, n70184, n68951, n68953, n68966, n68960, n68962, n68963,
    n68969, n68967, n68971, n68977, n68981, n69999, n68987, n68986, n68991,
    n68988, n68990, n68999, n75004, n69995, n69000, n98242, n69011, n69012,
    n71457, n69017, n69016, n69021, n69019, n69018, n69020, n69029, n69023,
    n69022, n69027, n69025, n69024, n69026, n69028, n69045, n69031, n69030,
    n69035, n69033, n69032, n69034, n69043, n69037, n69036, n69041, n69039,
    n69038, n69040, n69042, n69044, n70205, n70204, n74457, n71177, n71671,
    n71368, n71385, n71373, n71382, n70004, n70006, n70009, n70008, n70175,
    n70021, n70012, n70015, n70014, n70019, n70017, n70018, n71227, n70024,
    n70025, n71232, n71329, n70026, n70106, n70027, n70031, n70030, n70032,
    n71303, n70073, n70034, n71243, n70036, n71258, n70037, n70039, n70046,
    n70040, n70045, n75999, n70041, n70042, n71517, n70044, n71259, n70048,
    n71242, n70051, n70050, n71246, n70055, n70056, n70058, n71275, n70061,
    n70065, n71278, n71283, n70070, n71284, n70072, n71239, n70085, n70076,
    n70078, n70086, n70079, n70092, n70081, n70083, n70084, n71300, n71308,
    n70088, n70091, n70090, n70093, n70094, n71307, n70100, n70101, n70104,
    n70103, n70109, n70116, n70111, n70114, n70115, n70117, n70120, n71335,
    n70121, n70123, n71223, n70127, n70132, n71352, n71341, n70126, n71216,
    n70131, n70130, n70133, n70134, n70142, n70137, n70136, n70140, n70139,
    n70141, n71219, n70155, n70153, n70147, n70151, n70150, n70154, n70152,
    n71206, n70156, n70157, n70161, n70159, n70163, n70162, n70168, n70167,
    n70169, n70171, n70172, n71196, n71194, n71191, n71193, n71369, n70177,
    n70181, n70183, n70185, n70189, n71377, n71383, n70194, n71189, n71406,
    n70197, n71455, n70207, n70206, n70211, n70209, n70208, n70210, n70235,
    n70213, n70212, n70215, n70214, n70217, n70216, n70233, n70219, n70218,
    n70223, n70221, n70220, n70222, n70231, n70225, n70224, n70229, n70227,
    n70226, n70228, n70230, n70232, n70234, n71454, n71456, n74458, n74762,
    n71688, n71173, n71184, n71178, n71179, n76082, n74204, n71673, n71195,
    n71654, n74238, n71201, n71204, n71207, n71640, n71639, n71638, n71209,
    n71208, n71211, n71215, n71214, n71488, n71489, n71362, n71217, n71218,
    n71222, n71220, n71225, n71226, n71224, n71229, n71228, n71497, n71326,
    n71231, n71332, n71233, n71235, n71606, n71605, n71324, n71236, n71596,
    n71238, n71241, n71244, n71245, n71513, n71247, n71249, n71527, n71254,
    n71250, n71253, n71252, n71255, n71257, n71534, n71261, n71260, n71537,
    n71262, n71263, n71508, n71266, n71267, n71270, n71511, n71272, n71271,
    n71273, n71502, n71276, n71277, n71503, n71281, n71280, n71548, n71564,
    n71282, n71285, n71286, n71549, n71292, n71291, n71290, n71571, n71580,
    n71296, n71297, n71299, n71306, n71302, n71301, n71304, n71305, n71578,
    n71590, n71309, n71587, n71312, n71311, n71322, n71316, n71314, n71318,
    n71317, n71319, n71321, n71320, n71598, n71323, n71337, n71328, n71331,
    n71330, n71333, n71334, n71612, n71610, n71336, n71614, n71339, n71338,
    n71340, n71342, n71348, n71355, n71344, n71620, n71618, n71626, n71346,
    n71347, n71360, n71351, n71350, n71354, n71353, n71356, n71357, n71359,
    n71636, n71653, n71367, n71366, n71665, n71666, n71482, n71370, n71376,
    n71375, n71380, n71378, n71379, n71386, n71485, n71393, n71476, n71395,
    n71399, n71396, n71400, n71470, n71471, n71411, n71408, n71407, n71409,
    n74212, n71425, n71424, n71429, n71427, n71426, n71428, n71437, n71431,
    n71430, n71435, n71433, n71432, n71434, n71436, n71453, n71439, n71438,
    n71443, n71441, n71440, n71442, n71451, n71445, n71444, n71449, n71447,
    n71446, n71448, n71450, n71452, n71705, n71704, n71741, n71472, n74460,
    n71475, n71477, n74451, n71480, n71484, n71486, n71493, n71491, n71490,
    n71495, n71494, n71498, n71499, n74400, n74962, n71504, n71505, n71509,
    n71510, n74319, n71514, n71515, n74309, n74307, n74317, n71518, n71519,
    n74291, n74290, n71531, n71522, n74279, n71523, n74270, n74271, n71525,
    n74274, n71528, n71529, n71530, n71532, n74296, n71538, n71535, n71536,
    n71539, n74299, n71541, n71540, n71542, n74316, n74322, n71543, n71544,
    n74329, n71551, n71558, n71560, n71567, n71556, n71557, n74337, n71550,
    n71554, n71552, n71553, n71555, n74335, n71563, n71562, n71566, n71565,
    n71569, n71568, n71570, n74349, n71573, n74352, n71574, n71576, n74267,
    n71579, n71583, n71581, n74266, n71585, n71584, n71586, n71594, n71592,
    n71591, n71593, n74262, n71595, n71599, n74364, n74362, n71601, n74366,
    n71602, n71604, n74373, n71607, n74374, n71609, n71611, n71613, n74378,
    n74377, n71615, n71617, n74393, n71625, n71624, n71629, n71621, n71622,
    n71623, n71628, n71627, n71630, n71631, n74256, n71632, n71634, n71637,
    n71642, n71641, n71644, n71643, n71645, n74440, n74432, n71649, n71651,
    n74247, n71652, n71656, n74232, n71661, n71662, n71663, n75008, n71667,
    n74454, n74462, n71670, n74463, n74203, n71674, n71677, n71679, n71680,
    n74211, n74207, n71682, n71687, n74728, n71685, n71686, n71689, n71690,
    n74756, n71695, n74475, n71707, n71706, n71711, n71709, n71708, n71710,
    n71735, n71715, n71713, n71712, n71714, n71717, n71716, n71733, n71719,
    n71718, n71723, n71721, n71720, n71722, n71731, n71725, n71724, n71729,
    n71727, n71726, n71728, n71730, n71732, n71734, n74474, n71744, n71743,
    n74508, n75028, n74205, n74732, n74218, n74214, n74213, n74215, n74737,
    n74223, n74224, n74225, n74237, n74227, n74230, n74228, n74229, n74231,
    n74235, n74233, n74234, n74236, n74244, n74242, n74239, n74241, n74243,
    n74783, n74252, n74251, n74776, n74766, n74444, n74258, n74257, n74259,
    n74937, n74950, n74263, n74264, n74268, n74897, n74896, n74358, n74272,
    n74273, n74800, n74275, n74821, n74278, n74282, n74280, n74281, n74283,
    n74286, n74285, n74287, n74289, n74802, n74292, n74293, n74294, n74842,
    n74297, n74298, n74301, n74845, n74303, n74302, n74304, n74856, n74306,
    n74305, n74311, n74308, n74310, n74855, n74312, n74313, n74858, n74862,
    n74321, n74318, n74320, n74325, n74323, n74324, n74327, n74795, n74794,
    n74333, n74331, n74334, n74340, n74339, n74338, n74342, n74341, n74878,
    n74876, n74344, n74345, n74347, n74891, n74350, n74351, n74892, n74355,
    n74354, n74895, n74356, n74357, n74899, n74359, n74789, n74363, n74365,
    n74904, n74369, n74907, n74371, n74370, n74372, n74917, n74375, n74916,
    n74379, n74923, n74919, n74924, n74381, n74385, n74383, n74382, n74384,
    n74390, n74386, n74388, n74387, n74389, n74392, n74394, n74931, n74398,
    n74397, n74935, n74399, n74413, n74401, n74403, n74405, n74956, n74406,
    n74408, n74958, n74410, n74412, n74963, n74414, n74415, n74429, n74418,
    n74417, n74423, n74421, n74419, n74420, n74422, n74427, n74425, n74424,
    n74426, n74428, n74957, n75932, n74433, n74435, n74439, n74438, n74441,
    n74970, n75930, n74442, n74773, n74775, n74443, n74764, n74449, n74450,
    n74453, n74455, n74758, n74751, n74459, n74750, n74461, n74464, n74465,
    n75064, n74477, n74476, n74481, n74479, n74478, n74480, n74489, n74483,
    n74482, n74487, n74485, n74484, n74486, n74488, n74505, n74491, n74490,
    n74495, n74493, n74492, n74494, n74503, n74497, n74496, n74501, n74499,
    n74498, n74500, n74502, n74504, n75065, n97721, n74509, n74510, n75026,
    n74729, n75020, n74731, n74740, n74734, n74736, n74746, n74745, n74741,
    n76220, n74742, n74744, n74748, n76217, n74755, n74753, n74752, n74757,
    n75019, n76205, n75018, n74765, n74768, n74767, n75910, n75906, n75901,
    n74772, n75017, n74777, n74779, n74778, n75921, n75918, n76194, n74781,
    n74784, n74786, n76197, n74791, n74792, n76160, n76161, n76159, n74796,
    n76114, n76112, n74871, n74801, n76096, n74803, n76019, n74805, n74809,
    n74810, n74807, n74808, n74814, n74811, n74813, n74816, n74815, n75992,
    n74817, n74818, n75993, n74819, n76105, n76106, n74825, n74823, n74826,
    n76109, n74828, n74827, n74829, n76097, n76095, n76094, n76127, n74833,
    n76126, n74836, n74837, n76129, n74839, n74838, n74840, n76089, n74843,
    n74844, n76090, n74848, n74847, n76093, n74849, n74850, n74851, n76147,
    n74853, n74852, n74854, n74860, n74857, n74859, n76146, n74861, n76117,
    n74864, n76118, n74866, n74867, n76121, n74869, n74868, n74870, n74872,
    n76116, n74874, n74873, n74875, n74887, n74877, n74879, n74884, n74883,
    n76151, n74888, n74886, n76150, n74889, n74890, n76139, n76138, n74893,
    n74894, n76136, n76133, n74898, n76132, n74900, n74901, n76135, n76158,
    n74909, n74905, n74906, n74908, n75990, n74910, n74912, n74911, n74913,
    n75985, n74914, n74922, n74918, n75982, n75979, n74921, n74927, n74926,
    n74925, n74929, n74928, n75977, n75976, n75975, n75967, n74933, n74934,
    n75970, n75971, n75968, n74941, n74947, n74936, n74953, n74938, n74940,
    n74942, n75965, n74944, n74943, n75925, n75961, n75924, n74946, n74949,
    n74952, n74951, n74954, n74955, n75950, n75954, n74969, n74959, n74968,
    n74961, n74965, n74964, n74966, n74967, n75953, n75928, n75931, n74983,
    n74972, n74977, n74971, n74973, n74975, n74974, n74981, n74979, n74978,
    n74980, n74984, n75938, n76181, n74991, n74985, n74990, n74986, n74988,
    n74993, n74987, n74989, n74997, n74992, n74994, n74995, n74996, n74998,
    n74999, n76192, n75015, n75003, n75013, n75011, n75009, n75010, n75012,
    n75014, n75916, n75016, n75915, n76204, n75075, n75023, n75025, n75024,
    n97668, n98286, n75073, n75071, n75027, n76225, n98287, n75029, n75030,
    n75069, n75032, n75031, n75037, n75035, n75034, n75036, n75045, n75039,
    n75038, n75043, n75041, n75040, n75042, n75044, n75063, n75047, n75046,
    n75051, n75049, n75048, n75050, n75061, n75054, n75053, n75059, n75057,
    n75056, n75058, n75060, n75062, n75067, n75066, n96922, n75068, n75070,
    n75072, n75074, P1_P1_U2721_Lock, input_0, input_1, AND_1, input_2,
    OR_2, input_3, AND_3, input_4, OR_4, input_5, OR_5, input_6, OR_6,
    input_7, OR_7, input_8, AND_8, input_9, OR_9, input_10, AND_10,
    input_11, OR_11, input_12, OR_12, input_13, AND_13, input_14, OR_14,
    input_15, AND_15, input_16, AND_16, input_17, AND_17, input_18, AND_18,
    input_19, OR_19, input_20, AND_20, input_21, AND_21, input_22, AND_22,
    input_23, AND_23, input_24, AND_24, input_25, OR_25, input_26, OR_26,
    input_27, AND_27, input_28, AND_28, input_29, AND_29, input_30, AND_30,
    input_31, AND_31, input_32, OR_32, input_33, AND_33, input_34, AND_34,
    input_35, OR_35, input_36, OR_36, input_37, AND_37, input_38, AND_38,
    input_39, AND_39, input_40, AND_40, input_41, AND_41, input_42, AND_42,
    input_43, AND_43, input_44, AND_44, input_45, AND_45, input_46, AND_46,
    input_47, AND_47, input_48, OR_48, input_49, AND_49, input_50, AND_50,
    input_51, AND_51, input_52, AND_52, input_53, AND_53, input_54, OR_54,
    input_55, OR_55, input_56, OR_56, input_57, OR_57, input_58, AND_58,
    input_59, OR_59, input_60, OR_60, input_61, OR_61, input_62, OR_62,
    input_63, OR_63, input_64, AND_64, input_65, OR_65, input_66, AND_66,
    input_67, AND_67, input_68, OR_68, input_69, OR_69, input_70, OR_70,
    input_71, AND_71, input_72, OR_72, input_73, OR_73, input_74, AND_74,
    input_75, OR_75, input_76, AND_76, input_77, OR_77, input_78, OR_78,
    input_79, AND_79, input_80, input_81, AND_81, input_82, OR_82,
    input_83, AND_83, input_84, OR_84, input_85, OR_85, input_86, OR_86,
    input_87, OR_87, input_88, AND_88, input_89, OR_89, input_90, AND_90,
    input_91, OR_91, input_92, OR_92, input_93, AND_93, input_94, OR_94,
    input_95, AND_95, input_96, AND_96, input_97, AND_97, input_98, AND_98,
    input_99, OR_99, input_100, AND_100, input_101, AND_101, input_102,
    AND_102, input_103, AND_103, input_104, AND_104, input_105, OR_105,
    input_106, OR_106, input_107, AND_107, input_108, AND_108, input_109,
    AND_109, input_110, AND_110, input_111, AND_111, input_112, OR_112,
    input_113, AND_113, input_114, AND_114, input_115, OR_115, input_116,
    OR_116, input_117, AND_117, input_118, AND_118, input_119, AND_119,
    input_120, AND_120, input_121, AND_121, input_122, AND_122, input_123,
    AND_123, input_124, AND_124, input_125, AND_125, input_126, AND_126,
    input_127, AND_127, input_128, OR_128, input_129, AND_129, input_130,
    AND_130, input_131, AND_131, input_132, AND_132, input_133, AND_133,
    input_134, OR_134, input_135, OR_135, input_136, OR_136, input_137,
    OR_137, input_138, AND_138, input_139, OR_139, input_140, OR_140,
    input_141, OR_141, input_142, OR_142, input_143, OR_143, input_144,
    AND_144, input_145, OR_145, input_146, AND_146, input_147, AND_147,
    input_148, OR_148, input_149, OR_149, input_150, OR_150, input_151,
    AND_151, input_152, OR_152, input_153, OR_153, input_154, AND_154,
    input_155, OR_155, input_156, AND_156, input_157, OR_157, input_158,
    OR_158, input_159, AND_159, AND_159_INV, CASOP;
  assign n60029 = ~n59806 | ~n74220;
  assign n67389 = ~n60471 | ~n60469;
  assign n74249 = ~n74431 ^ n74430;
  assign n74250 = ~n71651 | ~n71650;
  assign n74411 = ~n74260 | ~n71634;
  assign n74402 = ~n71500 | ~n71499;
  assign n76063 = ~n76028 | ~DIN_24_;
  assign n60391 = ~n71191 ^ n59969;
  assign n71659 = ~n76044;
  assign n59826 = ~n76051;
  assign n64666 = ~n64648 | ~n64647;
  assign n64646 = ~n60503;
  assign n60099 = ~n64136 | ~n64135;
  assign n60746 = n64479 & n64474;
  assign n64475 = ~n64527;
  assign n64530 = ~n64348 | ~n64315;
  assign n67227 = ~n64776 | ~n64775;
  assign n71298 = n71294 | n71238;
  assign n61148 = ~n64182 | ~n64183;
  assign n64350 = n76028 & DIN_14_;
  assign n97978 = ~n60791;
  assign n64163 = n63925 & n64180;
  assign n60274 = ~n64453 | ~n64452;
  assign n64744 = ~n67333 | ~n64627;
  assign n67854 = ~n67847 | ~n67308;
  assign n64444 = ~n64437 | ~n64436;
  assign n63124 = ~n63069 ^ n63068;
  assign n63069 = ~n63200 ^ n63204;
  assign n70069 = ~n70062 | ~n68866;
  assign n63200 = ~n63227 | ~n63023;
  assign n64095 = ~n64090 | ~n64092;
  assign n60986 = ~n71512 ^ n71513;
  assign n71512 = ~n71537 | ~n71262;
  assign n59789 = ~n63977;
  assign n61370 = ~n63599 | ~n63598;
  assign n64562 = ~n74396 & ~n59984;
  assign n63897 = ~n63647 ^ n63999;
  assign n63999 = ~n61383 | ~n63646;
  assign n59828 = ~n62938;
  assign n63434 = ~n63353 ^ n63352;
  assign n63632 = ~n74835 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n61570 = n64030 | n64029;
  assign n71397 = ~P4_DATAO_REG_2__SCAN_IN;
  assign n62965 = n62960 | n62961;
  assign n60408 = n63418 & n61081;
  assign n59835 = ~n63610;
  assign n59829 = ~n59831 & ~n59830;
  assign n64574 = n74804 | n74882;
  assign n59830 = ~n64266;
  assign n74835 = ~n63855;
  assign n59911 = ~n74830;
  assign n63724 = ~n64367;
  assign n59991 = ~n74812;
  assign n76045 = ~P4_DATAO_REG_9__SCAN_IN;
  assign n60623 = ~n74210 | ~n74211;
  assign n60899 = ~n67345 ^ n61361;
  assign n71664 = ~n71481;
  assign n67268 = ~n74812 & ~n67266;
  assign n67807 = n67812 | n67269;
  assign n70003 = ~n70001 | ~n70000;
  assign n71404 = ~n74763 & ~n76055;
  assign n63329 = ~n63240 | ~n63323;
  assign n63327 = ~n63329 ^ n63328;
  assign n64214 = ~n64211 | ~n64193;
  assign n59923 = ~n63624;
  assign n60214 = ~n59790 & ~n59789;
  assign n59790 = n63973 & n61159;
  assign n64008 = ~n64075 ^ n63896;
  assign n63613 = ~n64051 & ~n74820;
  assign n64645 = ~n60505 | ~n60503;
  assign n60503 = ~n59791 ^ n64480;
  assign n59791 = ~n64481;
  assign n60007 = n63319 & n63414;
  assign n61366 = ~n68779 | ~n60810;
  assign n64635 = ~n64549 ^ n60399;
  assign n63852 = ~n60249 | ~n63835;
  assign n60101 = n68775 & n68774;
  assign n68769 = ~n64800 | ~n61441;
  assign n60502 = ~n68769 | ~n67203;
  assign n64231 = n61252 & n64083;
  assign n59796 = ~n64786;
  assign n64787 = ~n59796 | ~n64784;
  assign n70143 = ~n70127 ^ n71216;
  assign n71294 = ~n71240 ^ n71239;
  assign n71187 = ~n59798 | ~n71671;
  assign n59798 = ~n60230 | ~n60231;
  assign n71265 = ~n70057 | ~n70056;
  assign n60844 = n61258 | n70072;
  assign n70035 = ~n68844 | ~n68843;
  assign n63441 = ~n63434 ^ n63433;
  assign n63162 = ~n63157 ^ n63158;
  assign n59799 = ~n63249;
  assign n60192 = ~n63160 & ~n59799;
  assign n70067 = n70066 | n70065;
  assign n68788 = n68791 & n68793;
  assign n63374 = ~n59800 | ~n63228;
  assign n59800 = ~n63222 | ~n63221;
  assign n60094 = ~n60259 | ~n60258;
  assign n71365 = ~n71364 ^ n71653;
  assign n64237 = n64236 | n64015;
  assign n61260 = ~n71571 | ~n71292;
  assign n63458 = n63460 | n63372;
  assign n71608 = n71324 | n71323;
  assign n63134 = n63136 | n63843;
  assign n68854 = n68852 | n68853;
  assign n68961 = n68958 | n68957;
  assign n63000 = n62999 | n62998;
  assign n63186 = n63284 & n63004;
  assign n60133 = n64264 & n64380;
  assign n60276 = n60278 & n64678;
  assign n64688 = ~n59999 | ~n64609;
  assign n60389 = ~n60078 ^ n61411;
  assign n60078 = n64613 & n64688;
  assign n60839 = ~n64597 | ~n59805;
  assign n59805 = ~n64599;
  assign n64599 = ~n67296 ^ n61484;
  assign n60388 = ~n60024 | ~n71474;
  assign n60024 = ~n71391 ^ n71485;
  assign n75900 = ~n61446 | ~n61445;
  assign n64578 = ~n64579;
  assign n61495 = n64579 & n60184;
  assign n64579 = n64575 & n64576;
  assign n59806 = n74218 & n74217;
  assign n60134 = n64263 & n64264;
  assign n64263 = ~n60497 & ~n60500;
  assign n71669 = ~n74456 | ~n71480;
  assign n60481 = n60482 & n64253;
  assign n61145 = n61147 & n61146;
  assign n59813 = ~n67223;
  assign n59814 = ~n67224;
  assign n67886 = ~n59814 | ~n59813;
  assign n60117 = ~n64508 | ~n61435;
  assign n61435 = ~n64507 | ~n64506;
  assign n59815 = ~n61572;
  assign n59816 = ~n64484;
  assign n64504 = ~n59816 | ~n59815;
  assign n63918 = n63662 & n63663;
  assign n63614 = ~n60177 | ~n63616;
  assign n64543 = n61090 | n64460;
  assign n60882 = n71187 & n71186;
  assign n67361 = n67744 | n67741;
  assign n63331 = n63246 & n63245;
  assign n64190 = ~n64184 | ~n64185;
  assign n64110 = ~n63928 ^ n63927;
  assign n71230 = ~P4_DATAO_REG_11__SCAN_IN;
  assign n71372 = ~n71369 ^ n60383;
  assign n61483 = ~n71487 | ~n61575;
  assign n64701 = ~n64032;
  assign n63863 = n63890 | n74835;
  assign n61474 = n63865 & n63857;
  assign n63619 = n61473 & n63416;
  assign n64022 = ~n63876 | ~n63875;
  assign n64614 = ~n64613 | ~n64612;
  assign n59827 = ~n70165;
  assign n70158 = ~n59827 | ~n59826;
  assign n68945 = ~n70148 ^ n70146;
  assign n62915 = n62890 | n62889;
  assign n63129 = ~n63553 | ~n63125;
  assign n64497 = ~n64496 | ~n64495;
  assign n62937 = ~n62939 ^ n59828;
  assign n61255 = ~n63876 | ~n59829;
  assign n59831 = ~n63875;
  assign n71696 = n71695 | n71694;
  assign n63581 = n63697 | n63696;
  assign n71410 = ~n71402 | ~n71403;
  assign n71402 = ~n69999 | ~n69998;
  assign n63941 = n72804 | n72805;
  assign n63620 = ~n63619 | ~n63618;
  assign n63478 = n63130 & n63212;
  assign n63935 = ~n59832 | ~n63585;
  assign n59832 = ~n63694 | ~n63693;
  assign n67939 = ~n67938 & ~n67937;
  assign n61410 = n60388 & n71393;
  assign n70174 = ~n71198 ^ n71199;
  assign n71199 = ~n70156 ^ n71203;
  assign n60937 = ~n68903 | ~n60629;
  assign n63882 = ~n59836 | ~n59835;
  assign n59836 = ~n63611;
  assign n63504 = ~n64032;
  assign n59837 = ~n67273;
  assign n67275 = ~n59837 | ~n64709;
  assign n64031 = n64026 & n64025;
  assign n68802 = n67246 & n67245;
  assign n60263 = ~n64262 ^ n60483;
  assign n64683 = ~n60032 | ~n64615;
  assign n70160 = n70157 & n70166;
  assign n63387 = n63345 & n63644;
  assign n68955 = ~n60652 ^ n68948;
  assign n63670 = ~n63662 | ~n61438;
  assign n64362 = ~DIN_1_ | ~P4_DATAO_REG_19__SCAN_IN;
  assign n59841 = ~n64131;
  assign n59842 = ~n64132;
  assign n64136 = ~n59842 | ~n59841;
  assign n71374 = n71377 & n70190;
  assign n59863 = ~n68807;
  assign n61443 = n68998 & n68999;
  assign n67255 = n67248 | n67247;
  assign n67853 = ~n67854 ^ n67855;
  assign n67860 = ~n67853 ^ n67317;
  assign n59846 = n63621 & n63620;
  assign n63287 = ~n63174 ^ n63175;
  assign n63284 = n63287 | n63003;
  assign n67751 = n67238 & n67237;
  assign n64566 = ~n64384 | ~n64383;
  assign n59850 = ~n64688 | ~n64687;
  assign n60077 = ~n64688 | ~n64687;
  assign n74790 = ~n74265 | ~n74264;
  assign n74336 = ~n74332 | ~n71547;
  assign n70047 = ~n60385 & ~n70045;
  assign n71575 = ~n74348 ^ n61018;
  assign n74348 = ~n61019 | ~n71559;
  assign n75984 = ~n75987 ^ n75985;
  assign n75987 = ~n75991 | ~n74913;
  assign n74277 = ~n64701;
  assign n60455 = ~n76217 ^ n76218;
  assign n63436 = n63441 | n63440;
  assign n64297 = ~n64281 | ~n64422;
  assign n60486 = n60015 & n74226;
  assign n65183 = DIN_0_ | DIN_1_;
  assign n59854 = ~n71486 | ~n71485;
  assign n71487 = ~n71486 | ~n71485;
  assign n67799 = ~n67798 & ~n67797;
  assign n60093 = ~n64545 | ~n64544;
  assign n61147 = n64190 & n64189;
  assign n64049 = ~n64238 ^ n60924;
  assign n64240 = n64049 | n64048;
  assign n64238 = ~n60046 ^ n60380;
  assign n64457 = ~n61148 | ~n61147;
  assign n59857 = ~n61473 | ~n63602;
  assign n59858 = ~n61473 | ~n63602;
  assign n63886 = ~n61473 | ~n63602;
  assign n60032 = ~n64614 ^ n61411;
  assign n60880 = n68809 & n68808;
  assign n59859 = ~n70019 | ~n70018;
  assign n59860 = ~n70019 | ~n70018;
  assign n59861 = ~n70111;
  assign n71213 = ~n70019 | ~n70018;
  assign n61361 = ~n68801;
  assign n59862 = ~n64761 ^ n64759;
  assign n68806 = ~n59864 & ~n59863;
  assign n59864 = ~n68798 & ~n68799;
  assign n60832 = n64565 & n64424;
  assign n71619 = ~n71340 | ~n71614;
  assign n67296 = ~n67292;
  assign n59865 = n70021 & n70012;
  assign n59866 = ~n67776 | ~n67775;
  assign n59867 = ~n59854 | ~n61575;
  assign n59868 = ~n74210;
  assign n59869 = ~n59868;
  assign n59870 = SEL & DIN_2_;
  assign n68927 = ~n67776 | ~n67775;
  assign n60478 = ~n60480;
  assign n64717 = ~n67274;
  assign n64409 = ~n76062 & ~n59910;
  assign n63270 = ~n63351 ^ n63259;
  assign n74416 = ~P4_DATAO_REG_10__SCAN_IN;
  assign n64758 = ~n64761 ^ n64759;
  assign n76064 = ~P4_DATAO_REG_7__SCAN_IN;
  assign n61389 = ~n61390 ^ n74249;
  assign n76182 = ~n75949 ^ n75928;
  assign n74846 = ~n63005;
  assign n74361 = ~P4_DATAO_REG_17__SCAN_IN;
  assign n74396 = ~P4_DATAO_REG_13__SCAN_IN;
  assign n59892 = n64412 & n64411;
  assign n59893 = n62927 | n62882;
  assign n59896 = n64037 & n59870;
  assign n59961 = ~n64677;
  assign n59897 = n64355 ^ n64349;
  assign n59912 = ~n74830;
  assign n59901 = n67293 ^ n64725;
  assign n63483 = n63114 | n63113;
  assign n63202 = ~n63066 ^ n63067;
  assign n59902 = n60512 & n63963;
  assign n59903 = n64150 ^ n64173;
  assign n59904 = n64315 & n59974;
  assign n67364 = ~n67363 | ~n67362;
  assign n63282 = ~n63313 ^ n61349;
  assign n59995 = ~n67327 ^ n59996;
  assign n64038 = n63504 & P4_DATAO_REG_17__SCAN_IN;
  assign n64643 = ~n60034 ^ n61135;
  assign n64748 = ~n60135 | ~n64628;
  assign n67360 = ~n60098 ^ n67225;
  assign n61149 = ~n64669 ^ n64535;
  assign n67776 = ~n67772 | ~n67771;
  assign n60034 = ~n67205 ^ n59976;
  assign n59997 = ~n59998 ^ n60673;
  assign n74739 = n60023 & n74746;
  assign n64157 = ~n64144 | ~n64142;
  assign n64144 = n63827 | n63826;
  assign n64523 = ~n64179 | ~n64178;
  assign n63656 = ~n63898 ^ n63974;
  assign n63898 = ~n63655 | ~n63654;
  assign n59905 = ~n75995;
  assign n59906 = ~n75995;
  assign n59907 = ~n75995;
  assign n59908 = ~n75995;
  assign n59909 = ~n75995;
  assign n59910 = ~n74830;
  assign n74830 = SEL & DIN_4_;
  assign n75995 = ~n74830;
  assign n59994 = ~n59995 ^ n67770;
  assign n70178 = ~n71368 ^ n70004;
  assign n70074 = ~n70028 ^ n70029;
  assign n70028 = ~n60638 ^ n70069;
  assign n74774 = ~n75932 ^ n74976;
  assign n61161 = ~n64548 ^ n61162;
  assign n60087 = ~n67222 | ~n67221;
  assign n68875 = ~n60444 ^ n68876;
  assign n60444 = ~n67822 | ~n68871;
  assign n71198 = ~n60639 | ~n70171;
  assign n64307 = ~n64231;
  assign n60025 = ~n60024;
  assign n60022 = ~n60642 | ~n74770;
  assign n63912 = ~n63656 ^ n63899;
  assign n67331 = n59997 | n60672;
  assign n64011 = n60279 | n63632;
  assign n60279 = ~n63631 ^ n63891;
  assign n60185 = ~n64162 | ~n64161;
  assign n64208 = ~n64088 | ~n64313;
  assign n71248 = DIN_0_ & DIN_1_;
  assign n60863 = ~n64770 ^ n60082;
  assign n64770 = ~n60086 | ~n60083;
  assign n64387 = ~n60479 | ~n60481;
  assign n63847 = ~n63840 & ~n63839;
  assign n64452 = ~n64451 | ~n64450;
  assign n74119 = ~n64496 ^ n64495;
  assign n59913 = ~n63317;
  assign n59914 = ~n63317;
  assign n63317 = ~n64259;
  assign n60096 = ~n60222 | ~n60220;
  assign n71589 = ~n71577 ^ n71578;
  assign n71577 = ~n61260 ^ n71580;
  assign n64568 = ~n64379 | ~n64378;
  assign n67359 = ~n67751 ^ n67750;
  assign n70148 = ~n68823 | ~n68824;
  assign n64573 = n64032 & n60493;
  assign n67827 = ~n67282 | ~n67281;
  assign n64281 = n64280 | n64279;
  assign n68894 = ~n67858 | ~n67857;
  assign n68895 = ~n60038 | ~n68889;
  assign n64659 = ~n60117 ^ n64661;
  assign n67358 = ~n60176 ^ n67880;
  assign n63976 = n63897 | n63898;
  assign n59915 = ~n63504;
  assign n64652 = ~n64655 ^ n64653;
  assign n74431 = ~n74436 ^ n74437;
  assign n67842 = ~n68882 ^ n68881;
  assign n68882 = ~n60938 | ~n67838;
  assign n70191 = ~n70177 ^ n70178;
  assign n63849 = ~n63638 | ~n63637;
  assign n74409 = ~n74402 ^ n74400;
  assign n75949 = ~n75925 ^ n74946;
  assign n68766 = n67916 & n68776;
  assign n67916 = ~n60092 ^ n68958;
  assign n71597 = ~n71588 ^ n71587;
  assign n71588 = ~n71589 ^ n71590;
  assign n60452 = ~n74742 & ~n60453;
  assign n74220 = ~n60453 | ~n74737;
  assign n60626 = n61436 & n60494;
  assign n71697 = n71692 & n74756;
  assign n71683 = ~n74211;
  assign n74749 = ~n74464 | ~n60496;
  assign n71692 = n71693 | n74458;
  assign n71175 = n71180 | n69000;
  assign n69996 = ~n69999 | ~n68982;
  assign n74446 = ~n75007 ^ n71667;
  assign n67920 = n67919 | n67918;
  assign n71390 = n71386 | n71385;
  assign n67197 = ~n61346 | ~n61347;
  assign n74248 = ~n74249 ^ n74250;
  assign n68956 = ~n60266 ^ n68949;
  assign n61319 = ~n68784 | ~n68783;
  assign n60283 = n67746 & n67745;
  assign n60281 = ~n60098 ^ n59970;
  assign n68782 = ~n61323 ^ n61322;
  assign n64115 = ~n64127 ^ n61348;
  assign n64795 = n67205 | n67214;
  assign n64472 = n64471 & n59974;
  assign n64463 = n64530 | n64470;
  assign n60090 = n60088 & n59972;
  assign n67236 = n67233 & n59972;
  assign n60103 = ~n59904 | ~n64348;
  assign n60089 = n64775 & n59980;
  assign n60915 = ~n67346 | ~n64765;
  assign n64460 = n64459 & n64458;
  assign n61442 = ~n60091 ^ n61487;
  assign n60136 = ~n59862 ^ n64757;
  assign n64549 = n60403 & n60400;
  assign n63924 = ~n63920 ^ n64100;
  assign n70107 = ~n60037 | ~n68917;
  assign n60037 = n68914 & n68913;
  assign n60233 = ~n63672 | ~n63671;
  assign n70022 = ~n70102 | ~n60016;
  assign n64209 = ~n63985 | ~n63984;
  assign n60928 = n63917 | n63916;
  assign n68891 = ~n70098 ^ n70099;
  assign n63488 = n63117 | n63486;
  assign n67321 = ~n59954 | ~n60076;
  assign n63837 = ~n60226 | ~n63296;
  assign n67849 = n61357 & n67843;
  assign n61159 = ~n64220 ^ n60405;
  assign n63226 = n63225 & n63296;
  assign n64282 = n64058 & n64057;
  assign n60225 = n63646 & n59984;
  assign n60451 = ~n60174 ^ n59993;
  assign n63390 = ~n60506 | ~n60509;
  assign n60506 = n60507 & n60508;
  assign n63351 = ~n61365 | ~n63346;
  assign n63337 = ~n63427 ^ n63426;
  assign n60492 = n64699 | n64698;
  assign n67278 = ~n60949 | ~n60947;
  assign n60264 = ~n60265 & ~n59896;
  assign n60417 = n63327 | n63241;
  assign n63247 = ~n63327 ^ n63242;
  assign n63246 = n63153 | n63152;
  assign n64817 = P1_P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | n100123;
  assign n60465 = n60466 & n59991;
  assign n67781 = n59991 & n67778;
  assign n59976 = ~n67214;
  assign n64577 = ~n64718 ^ n64717;
  assign n60497 = ~n60498 | ~n59991;
  assign n64065 = ~n71230 & ~n59984;
  assign n71483 = ~n74771 & ~n76055;
  assign n59980 = ~n64350;
  assign n74798 = ~n76012;
  assign n74730 = ~n74729 & ~n74728;
  assign n59984 = ~n74315;
  assign n59930 = ~n63706;
  assign n76054 = n76028 & DIN_12_;
  assign n76037 = n76028 & DIN_13_;
  assign n74315 = n76028 & DIN_7_;
  assign n59935 = ~n61527;
  assign n59936 = ~n65136;
  assign n59937 = ~n64827;
  assign n59938 = ~n60788;
  assign n60500 = ~n64701 & ~n60501;
  assign n76051 = n76028 & DIN_17_;
  assign n64694 = ~n60722 | ~P4_DATAO_REG_19__SCAN_IN;
  assign n64697 = n71293 | n64572;
  assign n64369 = ~DIN_0_ | ~P4_DATAO_REG_20__SCAN_IN;
  assign n59940 = ~n64572;
  assign n74747 = n61577 | n74746;
  assign n76213 = ~n60413 | ~n74757;
  assign n61577 = ~n74738 | ~n74737;
  assign n71684 = ~n71683 ^ n71682;
  assign n61491 = ~n74738;
  assign n60467 = ~n71696 | ~n71697;
  assign n60414 = n74754 & n60415;
  assign n74754 = n74753 | n74752;
  assign n71691 = n71687 & n71686;
  assign n71694 = ~n71184 | ~n71183;
  assign n71183 = n71182 & n71181;
  assign n71172 = ~n71176;
  assign n71176 = ~n71676 ^ n61440;
  assign n60188 = n71186 & n74204;
  assign n71478 = n71477 & n74451;
  assign n69992 = ~n60456 | ~n68765;
  assign n71678 = n71674 & n71673;
  assign n74769 = n74768 | n74767;
  assign n69991 = n71180 & n69000;
  assign n60231 = n61444 & n61261;
  assign n61444 = ~n61443 | ~n60934;
  assign n67940 = n68765 & n67927;
  assign n71180 = ~n61443 ^ n60131;
  assign n60131 = ~n69996 ^ n69995;
  assign n71403 = ~n71405 ^ n70197;
  assign n67927 = n67926 | n67925;
  assign n61261 = ~n69996 | ~n69995;
  assign n59942 = ~n71474;
  assign n68765 = n67923 | n67924;
  assign n74785 = ~n74246 | ~n74245;
  assign n67933 = n67932 | n67931;
  assign n67937 = n67936 & n67935;
  assign n68998 = ~n68997 | ~n68996;
  assign n68996 = ~n67732 | ~n68983;
  assign n75941 = ~n61574 | ~n74982;
  assign n68997 = n68995 & n68994;
  assign n67935 = n67929 | n67930;
  assign n74246 = n60865 & n74236;
  assign n68993 = n68991 & n68990;
  assign n74222 = n74221 & n75004;
  assign n67929 = ~n67380 ^ n68989;
  assign n68980 = ~n68974 | ~n68973;
  assign n68995 = n68989 | n68985;
  assign n67928 = n67391 & n67390;
  assign n67936 = n67385 & n67384;
  assign n68974 = ~n67921 | ~n67920;
  assign n67380 = ~n68985 ^ n67202;
  assign n68976 = n68975 | n76044;
  assign n67382 = n67387 | n64658;
  assign n61131 = ~n67378 | ~n67379;
  assign n60469 = n60470 & n78645;
  assign n74254 = n74248 | n74247;
  assign n74253 = n74252 | n74251;
  assign n67193 = ~n67197 | ~n67195;
  assign n71657 = ~n60395 | ~n60394;
  assign n75933 = ~n74441 | ~n74440;
  assign n60395 = ~n60392 | ~n60391;
  assign n67375 = ~n67367;
  assign n67367 = ~n64801 ^ n67203;
  assign n74430 = ~n74434 ^ n74432;
  assign n68771 = ~n67738 | ~n67737;
  assign n74437 = ~n71645 | ~n74440;
  assign n64332 = n64331 | n64330;
  assign n70190 = n70189 | n70188;
  assign n60462 = n76793 & n60463;
  assign n67371 = n64663 & n64662;
  assign n76793 = ~n64329 ^ n64330;
  assign n64800 = ~n60209;
  assign n64508 = n64502 & n64501;
  assign n64663 = ~n64486 | ~n64485;
  assign n74945 = n74944 | n74943;
  assign n67899 = n67897 & n67904;
  assign n60209 = ~n60056 | ~n61138;
  assign n64329 = ~n64328 ^ n64489;
  assign n74960 = ~n71495 | ~n71494;
  assign n64661 = ~n64650 ^ n64649;
  assign n68949 = ~n68782 ^ n67895;
  assign n64487 = ~n64504 | ~n64662;
  assign n67219 = n67212 & n67211;
  assign n73153 = ~n64125 ^ n64124;
  assign n64125 = ~n63941 | ~n63940;
  assign n60050 = ~n67364;
  assign n67216 = n67215 & n67214;
  assign n67215 = ~n60234 | ~n60223;
  assign n71492 = ~n71500 | ~n60995;
  assign n72804 = ~n63939 ^ n63938;
  assign n67748 = ~n60281 ^ n67889;
  assign n64325 = n64130 & n64116;
  assign n63939 = ~n63792 | ~n63791;
  assign n64116 = n64115 | n60806;
  assign n64130 = ~n64115 | ~n60806;
  assign n64481 = ~n64512 ^ n64515;
  assign n63792 = n70254 | n70255;
  assign n70145 = ~n71213 ^ n71212;
  assign n64321 = n64122 | n64121;
  assign n61322 = ~n68789;
  assign n61323 = ~n61324 ^ n68793;
  assign n70254 = ~n60458 ^ n63790;
  assign n64127 = ~n64114 | ~n64113;
  assign n64336 = n64335 & n64334;
  assign n64122 = ~n63931 ^ n63930;
  assign n71496 = ~n71229 | ~n71228;
  assign n68789 = ~n67885 ^ n67884;
  assign n60458 = ~n63933 ^ n63932;
  assign n64343 = n64342 | n61535;
  assign n63933 = ~n63935 ^ n63934;
  assign n75991 = n74912 | n74911;
  assign n67223 = ~n64675 | ~n60093;
  assign n60123 = ~n64342 ^ n61535;
  assign n71210 = ~n71227 ^ n70144;
  assign n64517 = n64516 & n64515;
  assign n74920 = ~n74917 ^ n61452;
  assign n64112 = ~n63809 | ~n61573;
  assign n64132 = ~n64133 ^ n64134;
  assign n64790 = n64783 & n64782;
  assign n71358 = n71221 | n71220;
  assign n64533 = n64532 & n64531;
  assign n63809 = n63805 & n63804;
  assign n63934 = ~n63692 ^ n63691;
  assign n63585 = n63584 | n63583;
  assign n70011 = ~n60191 ^ n61358;
  assign n68822 = ~n68806 | ~n68805;
  assign n63584 = ~n63589 | ~n63477;
  assign n64477 = n64530 & n64470;
  assign n60102 = ~n60103 | ~n64526;
  assign n60235 = ~n64316 ^ n64530;
  assign n60191 = ~n68828 | ~n68827;
  assign n63802 = n63801 & n63800;
  assign n63589 = n63796 | n63475;
  assign n64531 = n64530 | n64529;
  assign n60040 = ~n64530 | ~n64525;
  assign n63477 = n63798 | n63476;
  assign n64133 = ~n60513 | ~n63953;
  assign n74903 = ~n61457 | ~n61455;
  assign n61452 = ~n74916;
  assign n63799 = ~n61439 | ~n63588;
  assign n61455 = n74789 | n61456;
  assign n61090 = ~n60097 ^ n64537;
  assign n67228 = ~n64768 ^ n60136;
  assign n64775 = ~n64537 | ~n64536;
  assign n60513 = ~n60514 | ~n63947;
  assign n63570 = n63699 | n63698;
  assign n63928 = n63825 | n63824;
  assign n74902 = ~n74900 | ~n74901;
  assign n71221 = ~n71217 ^ n71349;
  assign n64105 = n64166 | n64104;
  assign n63952 = n63949 & n63948;
  assign n60097 = ~n64635 ^ n64352;
  assign n60091 = ~n64207 & ~n64206;
  assign n71349 = ~n71335 | ~n70123;
  assign n76137 = ~n76139 ^ n76138;
  assign n61367 = ~n64163 ^ n64104;
  assign n63946 = n60095 | n63945;
  assign n64166 = ~n64163;
  assign n60086 = ~n60267 | ~n64549;
  assign n64165 = ~n63834 | ~n63833;
  assign n64182 = n64185 | n64181;
  assign n71343 = ~n70132 | ~n70125;
  assign n60083 = ~n60085 | ~n60084;
  assign n63303 = ~n63213 | ~n63212;
  assign n60400 = ~n60402 | ~n60401;
  assign n60403 = ~n64356 | ~n64355;
  assign n71603 = ~n74261 ^ n61002;
  assign n64761 = ~n64748 | ~n64629;
  assign n63834 = ~n63831 | ~n63830;
  assign n63831 = ~n60232 | ~n63672;
  assign n60402 = ~n64353;
  assign n60459 = ~n63557 | ~n63556;
  assign n63587 = ~n63474 ^ n63473;
  assign n64180 = ~n63924 | ~n63923;
  assign n64759 = n64634 & n64633;
  assign n60232 = n63666 & n63671;
  assign n74269 = n71585 | n71584;
  assign n64633 = ~n60273 | ~n64632;
  assign n63685 = n63684 & n63683;
  assign n70119 = ~n71327 ^ n70106;
  assign n61002 = ~n74262 ^ n71595;
  assign n71327 = ~n70105 | ~n71237;
  assign n60033 = n63993 & n60212;
  assign n60271 = ~n60268 | ~n64632;
  assign n63829 = ~n60233 ^ n63673;
  assign n60270 = n64452 & n60272;
  assign n60212 = ~n64211 | ~n60213;
  assign n74885 = n74884 | n74883;
  assign n70124 = ~n68923 | ~n68922;
  assign n63681 = ~n63472 | ~n63471;
  assign n68926 = ~n67873 ^ n67872;
  assign n63554 = n63553 & n63552;
  assign n71237 = ~n60386 | ~n60387;
  assign n63552 = n63551 | n63550;
  assign n64100 = ~n60927 | ~n63919;
  assign n63666 = ~n61134 | ~n61133;
  assign n63993 = n63988 & n63987;
  assign n63591 = ~n61343 | ~n63467;
  assign n60629 = ~n68899 | ~n68900;
  assign n60058 = ~n64450;
  assign n64626 = n64625 & n64624;
  assign n64450 = ~n64313 | ~n64312;
  assign n60927 = ~n60928 | ~n63918;
  assign n68918 = n67871 & n67870;
  assign n60213 = ~n64209 & ~n63992;
  assign n68917 = ~n70108 | ~n68916;
  assign n68919 = n68921 | n68920;
  assign n74880 = ~n74343 | ~n74344;
  assign n63470 = ~n63376 ^ n63375;
  assign n63465 = n63464 & n63463;
  assign n64088 = n64087 | n64086;
  assign n60376 = ~n64445;
  assign n64312 = n64311 | n64310;
  assign n64235 = n64228 & n64229;
  assign n70097 = n60381 | n70096;
  assign n71313 = n70102 & n70101;
  assign n60183 = ~n70110 ^ n70113;
  assign n60016 = ~n60018 | ~n60017;
  assign n70112 = ~n70108;
  assign n63219 = n63215 | n63214;
  assign n74797 = n74333 | n74334;
  assign n64446 = ~n64444 ^ n64443;
  assign n60018 = ~n68891;
  assign n63460 = ~n63374 ^ n63373;
  assign n61019 = n71556 & n71555;
  assign n60382 = ~n71307;
  assign n63669 = ~n63455 | ~n63454;
  assign n63968 = ~n60224;
  assign n60224 = ~n63847 | ~n60211;
  assign n60043 = ~n60045 | ~n60044;
  assign n63454 = n63453 | n63452;
  assign n60017 = ~n68890;
  assign n60210 = n60211 & n61158;
  assign n64301 = ~n64300 | ~n64299;
  assign n63216 = ~n63222 ^ n60853;
  assign n71559 = ~n71558 | ~n74335;
  assign n60277 = ~n64676 | ~n64677;
  assign n74865 = n74326 | n74327;
  assign n60044 = ~n63907;
  assign n63222 = ~n63140 & ~n63139;
  assign n61141 = ~n67322 | ~n67321;
  assign n63449 = n63450 | n63451;
  assign n60211 = ~n63846 | ~n63998;
  assign n60045 = ~n63908;
  assign n63448 = n63369 & n63368;
  assign n63450 = ~n63359 ^ n63358;
  assign n64679 = ~n60389 | ~n64610;
  assign n71289 = n71298 & n71241;
  assign n63139 = n63224 & n63138;
  assign n74863 = ~n74314 | ~n74858;
  assign n61372 = ~n60895 ^ n64427;
  assign n60404 = ~n61159;
  assign n63445 = n63438 | n63439;
  assign n63358 = ~n63438;
  assign n63117 = ~n63112 ^ n63111;
  assign n74332 = n71546 | n71545;
  assign n67855 = n67315 & n67316;
  assign n71546 = n71506 & n71505;
  assign n63439 = ~n63441 ^ n63354;
  assign n63438 = n61136 & n63357;
  assign n63111 = ~n63110 | ~n63109;
  assign n60218 = n60216 & n61383;
  assign n60226 = ~n60225 | ~n61383;
  assign n61357 = ~n67839 | ~n67840;
  assign n70087 = ~n60446 | ~n60445;
  assign n63651 = ~n61383 | ~n61129;
  assign n60895 = ~n64288 | ~n64287;
  assign n71295 = ~n70077 | ~n70032;
  assign n64288 = ~n64283 | ~n64282;
  assign n60446 = n60447 & n68834;
  assign n63368 = n63367 | n63366;
  assign n67309 = ~n67312;
  assign n70077 = n70074 | n70027;
  assign n64063 = n60180 & n64065;
  assign n59954 = ~n67320;
  assign n63106 = ~n63108 ^ n60051;
  assign n63355 = n63365 | n63356;
  assign n63433 = ~n63315 | ~n63314;
  assign n63223 = ~n63020 ^ n63019;
  assign n61130 = ~n63431 | ~n63430;
  assign n63365 = ~n63282 ^ n63310;
  assign n60216 = n63646 & n60217;
  assign n63495 = n63490 | n63491;
  assign n63431 = n63401 & n63400;
  assign n67845 = ~n67255 | ~n67254;
  assign n63019 = ~n63018 & ~n63017;
  assign n68837 = n68835 & n74315;
  assign n60182 = ~n61474 | ~n63858;
  assign n64608 = n60451 | n64416;
  assign n63386 = ~n63390 ^ n63389;
  assign n70080 = ~n67833 | ~n67834;
  assign n59955 = ~n68836;
  assign n64010 = ~n63895 | ~n64054;
  assign n63055 = n63104 | n63103;
  assign n67837 = ~n67830 ^ n67829;
  assign n68877 = ~n60443 | ~n60442;
  assign n68873 = ~n61359 | ~n67828;
  assign n60115 = ~n63642 ^ n63404;
  assign n60509 = ~n60510 | ~n63349;
  assign n71507 = ~n60840 | ~n71516;
  assign n74834 = n74293 | n74294;
  assign n63858 = ~n61511 | ~n63854;
  assign n60636 = ~n70069 ^ n60637;
  assign n61359 = ~n60858 | ~n67825;
  assign n63635 = n63424 & n63630;
  assign n60840 = ~n60985 | ~n60984;
  assign n60638 = ~n70068 ^ n68872;
  assign n60510 = ~n63351;
  assign n64054 = n63894 | n63893;
  assign n70066 = ~n71274 ^ n71275;
  assign n60637 = ~n70068;
  assign n63642 = ~n60096 | ~n63338;
  assign n64407 = n64276 & n64275;
  assign n70068 = n68871 & n68870;
  assign n63862 = n63861 & n63860;
  assign n67289 = ~n67284 | ~n67283;
  assign n71274 = ~n60379 ^ n71264;
  assign n70062 = n68865 | n68864;
  assign n63424 = n63423 | n63422;
  assign n63631 = ~n64052 ^ n63622;
  assign n63338 = ~n60219 | ~n63337;
  assign n63347 = n61365 & n63348;
  assign n67830 = ~n61150 ^ n67827;
  assign n62913 = n63026 | n63024;
  assign n62970 = ~n62966;
  assign n67284 = n67260 & n67282;
  assign n67283 = ~n67261 ^ n67262;
  assign n61249 = n64404 & n61251;
  assign n67831 = ~n67827 ^ n67826;
  assign n67822 = n67821 | n67820;
  assign n60924 = ~n64019 | ~n61259;
  assign n63277 = ~n63143 | ~n60847;
  assign n62966 = n62919 & n62918;
  assign n62984 = n62983 | n62982;
  assign n67261 = ~n60175 | ~n64700;
  assign n67282 = ~n67256 | ~n67257;
  assign n63093 = ~n63521 | ~n63088;
  assign n60175 = ~n60492 | ~n64697;
  assign n62918 = n62917 | n62916;
  assign n62964 = n62963 | n62962;
  assign n62911 = ~n60457 ^ n62891;
  assign n70052 = n70051 | n70050;
  assign n63268 = n63267 | n63266;
  assign n64273 = n64269 & n64268;
  assign n62979 = ~n62965 | ~n62958;
  assign n62981 = ~n62995 ^ n62994;
  assign n63255 = n63263 | n63250;
  assign n61362 = n63887 & n61363;
  assign n60457 = ~n62915 ^ n62917;
  assign n67824 = ~n60201 ^ n60200;
  assign n63521 = n63516 | n63517;
  assign n63343 = n63342 | n63341;
  assign n60877 = n64401 & n60878;
  assign n67256 = ~n67278 ^ n67279;
  assign n74799 = n74824 & n74287;
  assign n60201 = ~n67808 ^ n67813;
  assign n67801 = ~n68851 | ~n67785;
  assign n67808 = ~n60202 | ~n67276;
  assign n60200 = ~n67807 | ~n67805;
  assign n64699 = ~n64720 | ~n64696;
  assign n62994 = ~n62947 | ~n62946;
  assign n71520 = ~n60842 | ~n60841;
  assign n63340 = ~n63331 ^ n63247;
  assign n63160 = ~n63162 | ~n63163;
  assign n63167 = ~n63162 ^ n60039;
  assign n63263 = ~n63246 | ~n63154;
  assign n62917 = ~n62920 ^ n59893;
  assign n60202 = ~n67275 | ~n67274;
  assign n63624 = ~n60417 | ~n63330;
  assign n62995 = ~n62997 ^ n62955;
  assign n64587 = ~n64698;
  assign n60454 = n64610 & n64677;
  assign n60949 = n64712 & n60950;
  assign n62893 = ~n60464 | ~n59893;
  assign n62924 = n62920 | n59893;
  assign n63076 = ~n63039 | ~n63038;
  assign n61320 = ~n60134;
  assign n62920 = ~n62922 ^ n62921;
  assign n63039 = n63037 | n63036;
  assign n97991 = ~n64817;
  assign n60448 = n60450 & n60449;
  assign n67812 = ~n68857 ^ n68858;
  assign n60039 = ~n63163;
  assign n60577 = n63330 & n59911;
  assign n60464 = n60465 & n62884;
  assign n63157 = ~n61569 | ~n63152;
  assign n64581 = n60489 & n60488;
  assign n64712 = n64711 | n64710;
  assign n60084 = ~n60802;
  assign n61496 = ~n64577;
  assign n60082 = ~n64769;
  assign n60051 = ~n63107;
  assign n60450 = n67782 & n67780;
  assign n60631 = n60632 & n68842;
  assign n60265 = ~n64044 | ~n64035;
  assign n63841 = n63838 & P4_DATAO_REG_9__SCAN_IN;
  assign n60490 = ~n60184;
  assign n64632 = ~n59930 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n64196 = n59930 & P4_DATAO_REG_7__SCAN_IN;
  assign n97185 = ~n97204;
  assign n71197 = ~n71654 ^ n74238;
  assign n98007 = ~n64808;
  assign n70176 = ~n71192 ^ n71193;
  assign n70096 = n74798 & P4_DATAO_REG_17__SCAN_IN;
  assign n67752 = n74416 | n74367;
  assign n63152 = ~n62948 | ~n62986;
  assign n60221 = ~n63623;
  assign n97988 = ~n60796;
  assign n71212 = ~n74416 & ~n76061;
  assign n97987 = ~n61500;
  assign n98011 = ~n60792;
  assign n59967 = ~n67747;
  assign n97999 = ~n61526;
  assign n68928 = ~n76054 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n59969 = ~n71193;
  assign n98008 = ~n60788;
  assign n98002 = ~n65129;
  assign n71203 = ~n76051 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n97982 = ~n60799;
  assign n67880 = ~n63929 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n60630 = ~n68848 ^ n70038;
  assign n70043 = ~n60375 | ~P4_DATAO_REG_25__SCAN_IN;
  assign n59970 = ~n67890;
  assign n60449 = ~n67783;
  assign n67780 = n67779 | P4_DATAO_REG_24__SCAN_IN;
  assign n59972 = ~n67226;
  assign n74360 = ~n76054;
  assign n64249 = ~n60483;
  assign n64710 = n64709 & n60178;
  assign n67272 = ~n64709;
  assign n60262 = ~n64045;
  assign n60498 = ~n60499 | ~n74353;
  assign n63860 = n63856 & P4_DATAO_REG_12__SCAN_IN;
  assign n59974 = ~n64525;
  assign n76000 = ~n74881;
  assign n74367 = ~n76037;
  assign n60184 = ~n64694 ^ n64697;
  assign n60047 = ~n63496;
  assign n76067 = n76028 & DIN_18_;
  assign n64376 = n64367 & P4_DATAO_REG_18__SCAN_IN;
  assign n60483 = ~n64375 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n65136 = P1_P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | n100056;
  assign n64390 = ~n59940 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n65129 = n64836 | n64832;
  assign n97866 = ~n97998;
  assign n64808 = n100090 | n64832;
  assign n61527 = n96865 | n64824;
  assign n98052 = ~n100090 & ~n64824;
  assign n64827 = n64837 | n96865;
  assign n61526 = n64837 | n64835;
  assign n61500 = n64835 | n64832;
  assign n67287 = ~n74361 & ~n63855;
  assign n74806 = ~n74804;
  assign n64709 = n64367 & n60179;
  assign n60723 = ~n63317;
  assign n63874 = ~n74276 | ~n63412;
  assign n76012 = ~n76028 | ~DIN_9_;
  assign n74881 = ~n76028 | ~DIN_10_;
  assign n60375 = ~n63317;
  assign n71521 = ~n63317;
  assign n68848 = ~n67777 | ~n60634;
  assign n64706 = ~n64367;
  assign n64832 = ~P1_P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n100087;
  assign n100056 = n65089 | n99991;
  assign n71192 = n76076 & P4_DATAO_REG_6__SCAN_IN;
  assign n59986 = ~n74758;
  assign n64824 = ~P1_P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~n100136;
  assign n59988 = ~n74463;
  assign n64375 = ~n60721;
  assign n60517 = ~n74416;
  assign n61062 = ~DIN_1_ | ~n61063;
  assign n60179 = ~n74882;
  assign n60634 = n60715 & P4_DATAO_REG_24__SCAN_IN;
  assign n60501 = ~n71293;
  assign n68904 = ~P4_DATAO_REG_14__SCAN_IN;
  assign n63412 = P4_DATAO_REG_14__SCAN_IN & P4_DATAO_REG_15__SCAN_IN;
  assign n64250 = DIN_0_ & P4_DATAO_REG_16__SCAN_IN;
  assign n62986 = P4_DATAO_REG_10__SCAN_IN & P4_DATAO_REG_11__SCAN_IN;
  assign n67777 = SEL & P4_DATAO_REG_23__SCAN_IN;
  assign n59992 = ~n76076;
  assign n71171 = ~P4_DATAO_REG_0__SCAN_IN;
  assign n64572 = ~SEL | ~DIN_3_;
  assign n74763 = ~P4_DATAO_REG_3__SCAN_IN;
  assign n60721 = ~SEL | ~DIN_2_;
  assign n100090 = ~P1_P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n100136 = ~P1_P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n63855 = ~SEL | ~DIN_5_;
  assign n100087 = ~P1_P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n99991 = ~P1_P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n65089 = ~P1_P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n100072 = ~P1_P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n61063 = SEL & P4_DATAO_REG_19__SCAN_IN;
  assign n60715 = DIN_0_ & DIN_1_;
  assign n62928 = P4_DATAO_REG_9__SCAN_IN & P4_DATAO_REG_8__SCAN_IN;
  assign n60178 = ~P4_DATAO_REG_22__SCAN_IN;
  assign n60493 = ~P4_DATAO_REG_20__SCAN_IN;
  assign n60904 = ~SEL;
  assign n71188 = ~P4_DATAO_REG_1__SCAN_IN;
  assign n64607 = ~n60174 | ~n59993;
  assign n59993 = ~n64600 ^ n61065;
  assign n60079 = ~n67756 ^ n60650;
  assign n67756 = ~n59994 ^ n67762;
  assign n59996 = ~n67759;
  assign n67332 = ~n59997 | ~n60672;
  assign n67329 = ~n59998 | ~n67328;
  assign n64742 = ~n64736 ^ n59998;
  assign n59998 = ~n60819 ^ n64735;
  assign n64613 = n59999 | n64609;
  assign n64612 = ~n59999 | ~n64611;
  assign n59999 = ~n64685 ^ n64684;
  assign n71394 = ~n59942 | ~n60025;
  assign n70023 = ~n68898 | ~n68897;
  assign n67898 = ~n60836 | ~n59992;
  assign n71205 = ~n70153 | ~n70152;
  assign n68965 = ~n68964 | ~n68963;
  assign n67312 = ~n64733 | ~n64732;
  assign n64669 = ~n64534 | ~n64533;
  assign n64527 = n60006 & n64543;
  assign n60006 = ~n61371 | ~n64348;
  assign n68774 = ~n68773 & ~n68772;
  assign n63406 = ~n60007 | ~n63320;
  assign n60411 = ~n61082 | ~n63625;
  assign n60505 = n60008 & n64343;
  assign n60008 = ~n60099 | ~n64341;
  assign n64424 = n60132 | n64423;
  assign n63596 = ~n60009 ^ n63651;
  assign n60009 = ~n63652 ^ n63649;
  assign n60507 = ~n63347 | ~n63346;
  assign n64414 = ~n59892 | ~n64413;
  assign n64247 = ~n64251;
  assign n64252 = ~n64251 | ~n64250;
  assign n64251 = n64259 & P4_DATAO_REG_17__SCAN_IN;
  assign n64244 = ~n60013 | ~n60262;
  assign n60013 = ~n64242 ^ n60264;
  assign n64032 = ~SEL | ~DIN_0_;
  assign n60642 = ~n60643 | ~n74450;
  assign n60484 = ~n75002 ^ n74782;
  assign n60015 = ~n60861 | ~n74225;
  assign n61150 = ~n67824 ^ n67277;
  assign n70098 = ~n60019 | ~n70095;
  assign n60019 = ~n60198 | ~n60199;
  assign n67266 = ~n60020 | ~n67265;
  assign n60020 = ~n74804 | ~n75996;
  assign n75002 = ~n60485 | ~n60486;
  assign n64721 = ~n60021 ^ n67278;
  assign n60021 = ~n64716 ^ n64715;
  assign n74761 = ~n74760 | ~n60022;
  assign n74759 = ~n60022 ^ n74760;
  assign n60023 = ~n74735 | ~n74743;
  assign n60026 = ~n71475;
  assign n71479 = ~n60026 | ~n60025;
  assign n60487 = ~n60027 | ~n60625;
  assign n60027 = ~n60624 | ~n60028;
  assign n60028 = ~n60627 | ~n60816;
  assign n60627 = ~n60628 | ~n61436;
  assign n60624 = ~n60029 ^ n61491;
  assign n60639 = n70160 | n70159;
  assign n68779 = ~n60101 | ~n61254;
  assign n64089 = ~n60033 | ~n63994;
  assign n68768 = ~n68771;
  assign n74831 = ~n74802 | ~n60035;
  assign n60035 = ~n74288 | ~n74289;
  assign n74288 = ~n74800 ^ n74799;
  assign n74314 = ~n74312 | ~n74313;
  assign n60038 = ~n67850 | ~n67851;
  assign n61569 = n60518 & n60515;
  assign n60508 = ~n63349 | ~n63348;
  assign n63349 = ~n60846 | ~n63268;
  assign n60516 = ~n64701 & ~n60517;
  assign n60892 = ~n67740 | ~n67739;
  assign n64314 = ~n64457 ^ n61442;
  assign n64522 = ~n64527 | ~n60040;
  assign n64348 = n64314 | n61146;
  assign n68952 = ~n60041 | ~n67749;
  assign n60041 = ~n60282 | ~n60283;
  assign n60722 = ~n60721;
  assign n64512 = ~n60042 | ~n60746;
  assign n60042 = ~n64468 | ~n64469;
  assign n63910 = ~n60043 | ~n63906;
  assign n64662 = ~n64484 | ~n61572;
  assign n60046 = ~n64031 | ~n61570;
  assign n71240 = ~n60844 | ~n71287;
  assign n63097 = ~n60048 | ~n60047;
  assign n60048 = ~n63497;
  assign n63121 = ~n63120 | ~n60049;
  assign n60049 = ~n63483 | ~n63117;
  assign n60261 = ~n60050 ^ n67365;
  assign n67365 = ~n67360 ^ n67889;
  assign n63798 = ~n63588 ^ n63587;
  assign n60644 = ~n60484 ^ n60747;
  assign n63092 = ~n63093;
  assign n70071 = ~n60636 | ~n60635;
  assign n60056 = ~n60080 | ~n64666;
  assign n60336 = ~n67754 | ~n67755;
  assign n68939 = ~n60336 | ~n67757;
  assign n64565 = ~n60132 | ~n64423;
  assign n60132 = ~n64561 ^ n64562;
  assign n67800 = ~n67801;
  assign n60399 = ~n64455 ^ n61162;
  assign n67743 = ~n64672 | ~n60057;
  assign n60057 = ~n64671 | ~n60100;
  assign n60220 = ~n60229 ^ n60221;
  assign n61089 = ~n68971 | ~n61143;
  assign n61318 = ~n68965 | ~n68966;
  assign n60255 = ~n60874 | ~n70194;
  assign n61095 = ~n61486 | ~n61487;
  assign n61487 = ~n60253 ^ n59897;
  assign n64354 = ~n60058 ^ n64451;
  assign n64451 = ~n64305 ^ n64445;
  assign n60409 = ~n60411 | ~n60410;
  assign n61479 = ~n67909 | ~n67908;
  assign n71200 = n71199 | n71198;
  assign n61390 = ~n71652;
  assign n63845 = ~n60218 & ~n63842;
  assign n68773 = n68767 & n68766;
  assign n70192 = ~n60101 | ~n61253;
  assign n60080 = ~n64643 | ~n64642;
  assign n67735 = n60081 & n67914;
  assign n71364 = ~n60328 ^ n71197;
  assign n76218 = ~n75019 ^ n76211;
  assign n64593 = ~n60065 | ~n64566;
  assign n60065 = ~n64590;
  assign n64590 = ~n64568 ^ n64567;
  assign n61411 = ~n64565 | ~n64564;
  assign n67744 = ~n64792 ^ n64791;
  assign n63415 = ~n63601 ^ n63600;
  assign n63601 = ~n63413 | ~n63874;
  assign n67762 = ~n61038 | ~n67340;
  assign n68938 = ~n68826 ^ n60073;
  assign n60073 = ~n68825 | ~n68827;
  assign n67760 = ~n67758 | ~n67761;
  assign n70016 = ~n68942 | ~n68941;
  assign n74733 = ~n74749 | ~n74732;
  assign n67319 = ~n60077 | ~n67320;
  assign n60076 = ~n60077;
  assign n61164 = ~n59850 ^ n67318;
  assign n64682 = ~n61411 | ~n60078;
  assign n68798 = ~n60079 ^ n67753;
  assign n64650 = ~n61138 | ~n60080;
  assign n67738 = ~n60081 | ~n67736;
  assign n60081 = ~n60209 | ~n60208;
  assign n64768 = ~n60863;
  assign n60085 = ~n61161;
  assign n60098 = ~n60087 | ~n67886;
  assign n67888 = ~n67887 | ~n60087;
  assign n64774 = ~n64775 | ~n64776;
  assign n60088 = ~n60089 | ~n64776;
  assign n64783 = ~n60090 | ~n67228;
  assign n68957 = ~n60092;
  assign n67907 = ~n67903 | ~n60092;
  assign n60092 = ~n67219 | ~n67218;
  assign n64640 = ~n60093 | ~n64673;
  assign n68968 = ~n60094 | ~n61318;
  assign n71387 = ~n61142 | ~n60094;
  assign n61143 = ~n68970 | ~n60094;
  assign n63951 = ~n60095 | ~n63950;
  assign n63807 = n60095 & n63806;
  assign n63691 = ~n60095 ^ n63690;
  assign n63797 = ~n63795 & ~n60095;
  assign n60095 = ~n63810 ^ n63943;
  assign n63636 = ~n60096 | ~n63428;
  assign n67891 = ~n60098 | ~n59970;
  assign n64335 = ~n60123 ^ n60099;
  assign n60100 = ~n64670;
  assign n64347 = ~n64457 | ~n61442;
  assign n64532 = ~n64527 | ~n60102;
  assign n63345 = ~n60114 | ~n60116;
  assign n60114 = ~n60115;
  assign n63644 = ~n60115 | ~n63344;
  assign n60116 = ~n63344;
  assign n67377 = ~n60117 & ~n64661;
  assign n64342 = ~n64513 ^ n60736;
  assign n60252 = ~n60173 ^ n60134;
  assign n64384 = ~n60133 | ~n64263;
  assign n64389 = ~n64386 | ~n60134;
  assign n64629 = n60135 | n64628;
  assign n60135 = ~n64745 ^ n64744;
  assign n64772 = ~n60863 | ~n60136;
  assign n60230 = ~n71672;
  assign n67324 = ~n64683 | ~n64682;
  assign n67328 = ~n60275 | ~n64681;
  assign n64364 = ~n64362 & ~n64369;
  assign n71481 = ~n71380 | ~n71379;
  assign n67875 = n68802 | n68798;
  assign n64401 = ~n61320 | ~n60173;
  assign n64400 = ~n61320 & ~n60173;
  assign n60173 = ~n60851 | ~n64258;
  assign n60174 = ~n64415 | ~n64414;
  assign n67881 = ~n60899 | ~n60176;
  assign n67883 = n60899 | n60176;
  assign n60176 = ~n67356 | ~n67357;
  assign n63618 = ~n63617 | ~n60177;
  assign n63625 = ~n60177 | ~n63326;
  assign n60177 = ~n63325 | ~n63324;
  assign n60936 = ~n60182;
  assign n60180 = ~n64068 | ~n64066;
  assign n64068 = ~n60182 ^ n60181;
  assign n60181 = ~n64056;
  assign n68921 = ~n70108 ^ n60183;
  assign n64513 = ~n60185 ^ n60235;
  assign n64514 = ~n60235 | ~n60185;
  assign n60189 = ~n60186 | ~n71673;
  assign n60186 = ~n71187 | ~n71186;
  assign n71412 = ~n60189 | ~n60187;
  assign n60187 = ~n71187 | ~n60188;
  assign n74206 = ~n74205 | ~n60190;
  assign n60190 = ~n60882;
  assign n70020 = ~n61358 | ~n60191;
  assign n61365 = n63258 | n63257;
  assign n63257 = ~n63256 & ~n60192;
  assign n63258 = ~n63340 ^ n63248;
  assign n64367 = ~n60721;
  assign n70102 = ~n68891 | ~n68890;
  assign n70095 = ~n68885 | ~n68884;
  assign n60198 = ~n68884;
  assign n60199 = ~n68885;
  assign n60208 = ~n61441;
  assign n64211 = n60215 & n60214;
  assign n60215 = ~n63970 | ~n60404;
  assign n61383 = ~n60228 | ~n60227;
  assign n60217 = ~n63296;
  assign n60219 = ~n60220;
  assign n60222 = ~n63337;
  assign n64796 = ~n67205 | ~n67214;
  assign n60223 = ~n67205;
  assign n67205 = ~n61149 ^ n64670;
  assign n63972 = ~n60224 | ~n61158;
  assign n60763 = n60224 & n63980;
  assign n60227 = ~n63432;
  assign n60228 = ~n61130;
  assign n63627 = ~n60229 | ~n63623;
  assign n60229 = ~n63625 ^ n63624;
  assign n71672 = ~n71402 ^ n71403;
  assign n63833 = ~n60233 | ~n63832;
  assign n60234 = ~n61135;
  assign n61135 = ~n60931 | ~n64519;
  assign n63836 = n60249 | n63835;
  assign n63647 = ~n60249 ^ n63640;
  assign n60249 = ~n63849 ^ n63848;
  assign n64405 = n60252 | n60878;
  assign n60657 = ~n64403 ^ n60252;
  assign n61489 = ~n60253 ^ n61490;
  assign n60253 = ~n64353 ^ n64354;
  assign n71190 = ~n60255 | ~n71404;
  assign n71405 = ~n60255 | ~n71189;
  assign n60258 = ~n68966;
  assign n60259 = ~n68965;
  assign n67902 = ~n60261 | ~n76076;
  assign n67897 = ~n60261 | ~n60260;
  assign n60260 = ~n67901;
  assign n64242 = ~n60263 ^ n64034;
  assign n68954 = ~n60266 | ~n68949;
  assign n60266 = ~n68952 ^ n68950;
  assign n60267 = ~n61161 | ~n60802;
  assign n60268 = ~n64453 | ~n64452;
  assign n64548 = ~n60271 | ~n60269;
  assign n60269 = ~n60270 | ~n64453;
  assign n60272 = ~n64632;
  assign n64631 = ~n60274 | ~n59930;
  assign n60273 = ~n60274;
  assign n64455 = ~n60274 ^ n64454;
  assign n60278 = ~n61321;
  assign n60275 = ~n60276 | ~n60277;
  assign n63633 = ~n60279 | ~n63632;
  assign n60282 = ~n60280 | ~n59967;
  assign n60280 = ~n67748;
  assign n71648 = n60328 | n71649;
  assign n71650 = ~n60328 | ~n71649;
  assign n71655 = ~n60328 ^ n71654;
  assign n60328 = ~n71195 | ~n71196;
  assign n71363 = ~n71647 | ~n60334;
  assign n74434 = ~n60994 | ~n60334;
  assign n60334 = ~n71202 | ~n71201;
  assign n68821 = ~n60335 ^ n68938;
  assign n60335 = ~n68939 ^ n68936;
  assign n67238 = ~n60337 | ~n67232;
  assign n67224 = ~n67220 ^ n60337;
  assign n64792 = ~n67223 ^ n60337;
  assign n60337 = ~n64773 ^ n60651;
  assign n60519 = ~n71521 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n63077 = ~n60375 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n62879 = ~n60375 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n71251 = ~n60723 | ~P4_DATAO_REG_26__SCAN_IN;
  assign n62883 = ~n60375 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n64440 = ~n60376 | ~n64443;
  assign n64449 = ~n64446 ^ n60376;
  assign n71500 = ~n71361 | ~n60377;
  assign n60995 = n71361 | n60377;
  assign n60377 = ~n71360 ^ n60996;
  assign n64283 = ~n64286 ^ n64284;
  assign n60379 = ~n71265 ^ n70058;
  assign n71268 = ~n60378 | ~n70058;
  assign n60378 = ~n71264 ^ n71265;
  assign n64275 = ~n60380 | ~n64274;
  assign n60380 = ~n64270;
  assign n71310 = ~n60381 | ~n70096;
  assign n60381 = ~n71308 ^ n60382;
  assign n74436 = ~n71635 ^ n74411;
  assign n71384 = ~n71372 ^ n71373;
  assign n60383 = ~n71368;
  assign n70049 = ~n60384 | ~n70048;
  assign n60384 = ~n70047;
  assign n60385 = ~n70044 | ~n71517;
  assign n60386 = ~n70104;
  assign n60387 = ~n70103;
  assign n70122 = ~n70119;
  assign n71473 = n76038 & n60388;
  assign n71392 = ~n71394 | ~n60388;
  assign n74452 = ~n61036 | ~n60388;
  assign n64678 = ~n60389 | ~n60454;
  assign n67333 = ~n64626 | ~n60390;
  assign n64627 = n64626 | n60390;
  assign n60390 = ~n64738 ^ n64616;
  assign n60393 = ~n71368;
  assign n60392 = ~n60393 | ~n60396;
  assign n60394 = ~n71368 | ~n71192;
  assign n60396 = ~n71192;
  assign n60401 = ~n64354;
  assign n60405 = ~n64006;
  assign n63630 = ~n63423 | ~n63422;
  assign n63423 = ~n60409 & ~n60408;
  assign n60410 = ~n61080 | ~n63421;
  assign n60413 = ~n74755 | ~n74754;
  assign n76210 = ~n60414 | ~n74755;
  assign n60415 = ~n74757;
  assign n60859 = ~n60577 | ~n60417;
  assign n60889 = n60441 & n74206;
  assign n74210 = ~n74203 | ~n60441;
  assign n60441 = ~n71670 | ~n74463;
  assign n60442 = ~n68876;
  assign n60443 = ~n60444;
  assign n60445 = ~n68837 | ~n68836;
  assign n60447 = ~n59955 | ~n61392;
  assign n67784 = ~n67781 | ~n60450;
  assign n68851 = ~n60448 | ~n67781;
  assign n64417 = ~n60451 | ~n64416;
  assign n74735 = ~n74740 & ~n60453;
  assign n60453 = ~n60623 | ~n74219;
  assign n77917 = ~n60455 ^ n75020;
  assign n60456 = ~n67939 | ~n67940;
  assign n62919 = ~n60457 | ~n62914;
  assign n63487 = ~n63117 | ~n63486;
  assign n63112 = ~n63073 ^ n63072;
  assign n63791 = n60458 | n63790;
  assign n63562 = ~n60459 | ~n63700;
  assign n63772 = ~n60459 ^ n63701;
  assign n64333 = ~n60462 | ~n60461;
  assign n60461 = ~n73153 | ~n64126;
  assign n60463 = ~n64126 | ~n73154;
  assign n60466 = ~n59915 | ~n71660;
  assign n60628 = ~n60467 | ~n74466;
  assign n60471 = ~n74119 | ~n64497;
  assign n60470 = ~n64497 | ~n74120;
  assign n64391 = ~n60478 | ~n64249;
  assign n60480 = n64248 & n64247;
  assign n60479 = ~n60480 | ~n64252;
  assign n60482 = ~n60483 | ~n64252;
  assign n74782 = ~n74785 ^ n74783;
  assign n60485 = ~n60876 | ~n75007;
  assign n61446 = ~n60487;
  assign n75899 = ~n60487 | ~n74730;
  assign n67327 = ~n67865 ^ n67326;
  assign n67865 = ~n67866 ^ n67867;
  assign n60488 = ~n60490 | ~n64578;
  assign n60489 = ~n60490 | ~n64577;
  assign n70128 = ~n60491 ^ n70124;
  assign n60491 = ~n60937 ^ n70107;
  assign n70125 = n70124 | n60491;
  assign n60494 = ~n60816;
  assign n60496 = ~n74462 | ~n59988;
  assign n74804 = ~n64259;
  assign n74812 = ~n65183 | ~SEL;
  assign n60499 = ~n74806 | ~n60501;
  assign n67915 = ~n60716 | ~n60502;
  assign n68767 = ~n67735 | ~n60502;
  assign n64647 = ~n60504 | ~n64646;
  assign n60504 = ~n60505;
  assign n61572 = ~n60505 ^ n64483;
  assign n63350 = ~n63349;
  assign n64134 = ~n60511 ^ n59903;
  assign n60511 = ~n63964 | ~n59902;
  assign n60512 = ~n63967 | ~n63966;
  assign n60514 = ~n63946 | ~n61528;
  assign n60515 = ~n60516 & ~n74812;
  assign n60518 = ~n60519 | ~n71230;
  assign n71182 = ~n71176 | ~n60534;
  assign n60534 = ~n71175 | ~n71177;
  assign n71676 = ~n61350;
  assign n74216 = n60623 & n74215;
  assign n60625 = ~n60626 | ~n60628;
  assign n71234 = ~n60629 | ~n70025;
  assign n68846 = ~n60631 | ~n60630;
  assign n60632 = ~n60633 | ~n76007;
  assign n60633 = ~n59914 | ~P4_DATAO_REG_24__SCAN_IN;
  assign n60635 = ~n68872;
  assign n71202 = ~n71200 | ~n60639;
  assign n75007 = ~n60641;
  assign n60641 = ~n60944 ^ n61389;
  assign n75005 = ~n75007 | ~n60640;
  assign n60640 = ~n75006;
  assign n74226 = ~n60641 | ~n74222;
  assign n74770 = ~n60644 | ~n61478;
  assign n60643 = ~n60644;
  assign n76206 = ~n60647 | ~n74761;
  assign n60647 = ~n60648 | ~n59986;
  assign n60648 = ~n74759;
  assign n67755 = n67756 | n67752;
  assign n60650 = ~n67752;
  assign n67353 = ~n60651 | ~n60915;
  assign n67347 = ~n60651 | ~n60720;
  assign n60651 = ~n64772 | ~n64771;
  assign n70001 = n60652 | n61319;
  assign n60652 = ~n70184 ^ n68947;
  assign n70002 = ~n60652 | ~n61319;
  assign n71389 = ~n71388 | ~n60656;
  assign n70196 = ~n60656 ^ n71387;
  assign n60656 = ~n70191 ^ n71383;
  assign n63316 = ~n63504 & ~P4_DATAO_REG_13__SCAN_IN;
  assign n68841 = ~n63504 & ~P4_DATAO_REG_24__SCAN_IN;
  assign n64412 = n60657 | n64409;
  assign n64408 = n60657 & n64409;
  assign n64406 = ~n60657 ^ n64409;
  assign n60672 = ~n67330;
  assign n60673 = ~n67328;
  assign n60716 = n64800 | n61441;
  assign n67325 = ~n61164 ^ n59954;
  assign n60718 = ~n64218 | ~n64217;
  assign n64232 = ~n64218 | ~n64217;
  assign n60950 = n67273 | n64707;
  assign n60720 = n67346 & n64765;
  assign n67866 = ~n61243 | ~n61242;
  assign n63353 = ~n63387;
  assign n64019 = ~n61362 | ~n63888;
  assign n63156 = ~n74276 | ~n61554;
  assign n74822 = n62948 & n60774;
  assign n71381 = ~n71481 ^ n71483;
  assign n61412 = ~n64756 | ~n64755;
  assign n61137 = ~n63592 ^ n63591;
  assign n63592 = ~n63668 ^ n63456;
  assign n70173 = ~n70175;
  assign n68899 = ~n70022 ^ n70023;
  assign n64270 = n64244 & n64047;
  assign n60908 = ~n64303 | ~n64302;
  assign n64303 = ~n64357 ^ n64301;
  assign n74760 = ~n74456 | ~n74455;
  assign n63672 = n63668 | n63667;
  assign n68947 = ~n70182 ^ n70180;
  assign n74466 = ~n59869 ^ n71684;
  assign n61075 = ~n64742 ^ n67339;
  assign n64745 = ~n61475 | ~n64554;
  assign n64365 = ~n61062 | ~n61061;
  assign n61061 = ~SEL | ~P4_DATAO_REG_20__SCAN_IN;
  assign n64260 = n64259 & P4_DATAO_REG_19__SCAN_IN;
  assign n67295 = ~n67291;
  assign n64075 = ~n64011 | ~n64010;
  assign n61387 = ~n67831 ^ n67825;
  assign n61393 = ~n68830;
  assign n61394 = ~n61395 | ~n59984;
  assign n67847 = ~n61151 | ~n61152;
  assign n64557 = ~n60832;
  assign n67320 = ~n67312 ^ n64734;
  assign n61038 = ~n61039 | ~n67332;
  assign n74295 = ~n60998 | ~n71532;
  assign n67343 = ~n67341;
  assign n63144 = ~n62993 ^ n63164;
  assign n60856 = ~n60857 | ~n62994;
  assign n74326 = ~n74863 ^ n74862;
  assign n64183 = ~n64180;
  assign n74346 = ~n74797 | ~n61471;
  assign n64537 = ~n61095 | ~n61485;
  assign n63363 = ~n63295 | ~n63294;
  assign n63292 = n63291 & n63290;
  assign n64177 = n64174 & n64173;
  assign n71616 = ~n61009 | ~n61007;
  assign n61009 = ~n61014 | ~n61010;
  assign n61007 = ~n74373 | ~n61008;
  assign n70186 = ~n68954 | ~n68953;
  assign n61344 = ~n63458 | ~n63457;
  assign n71647 = n71202 | n71201;
  assign n71646 = ~n71636 ^ n71638;
  assign n63676 = ~n63679 | ~n63469;
  assign n69997 = ~n68980 | ~n68979;
  assign n61350 = ~n61444 | ~n61261;
  assign n64337 = ~n64130 | ~n64129;
  assign n64496 = ~n64333 | ~n64332;
  assign n64318 = ~n64323 | ~n64321;
  assign n76211 = ~n75018 ^ n76204;
  assign n61436 = ~n71691 | ~n71690;
  assign n64033 = ~n64250;
  assign n60893 = ~n64022;
  assign n64386 = n64385 & n64392;
  assign n61259 = ~n64018 | ~n64017;
  assign n64693 = ~n64694;
  assign n67791 = n68856 | n67788;
  assign n67273 = ~n64705 | ~n68856;
  assign n60948 = ~n67276;
  assign n61247 = ~n64405 | ~n64404;
  assign n67292 = n64593 & n64569;
  assign n63864 = ~n63863 | ~n63862;
  assign n60900 = ~n64376;
  assign n63407 = ~n64051 & ~n64706;
  assign n63878 = ~n63883;
  assign n63323 = ~n74276 | ~n61549;
  assign n63321 = P4_DATAO_REG_13__SCAN_IN & P4_DATAO_REG_14__SCAN_IN;
  assign n64051 = ~P4_DATAO_REG_12__SCAN_IN;
  assign n60858 = ~n67831;
  assign n67310 = ~n67248 ^ n67247;
  assign n64359 = ~n61372 ^ n64297;
  assign n64426 = ~n64297;
  assign n67833 = ~n61387 | ~n61386;
  assign n61386 = ~n67832;
  assign n71269 = ~n71507 ^ n71508;
  assign n61023 = ~n63504 & ~P4_DATAO_REG_27__SCAN_IN;
  assign n71545 = ~n74330 ^ n74329;
  assign n62942 = n74276 & n61555;
  assign n67339 = ~n67333 | ~n67335;
  assign n61243 = ~n61166 | ~n61165;
  assign n61165 = ~n67324;
  assign n71526 = ~n74270 ^ n74271;
  assign n71561 = ~n71506 | ~n60988;
  assign n60988 = ~n60990 | ~n60989;
  assign n60989 = ~n71280;
  assign n60990 = ~n71281;
  assign n61470 = ~n74821;
  assign n64753 = n61075 | n67338;
  assign n64755 = ~n74416 & ~n74360;
  assign n63432 = ~n63429 ^ n63636;
  assign n63429 = ~n63635 ^ n63634;
  assign n70135 = ~n61385 | ~n68931;
  assign n61385 = ~n68926 | ~n68925;
  assign n60841 = ~n71255;
  assign n61018 = ~n74349;
  assign n64204 = ~n64194 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n61485 = ~n61489 | ~n61488;
  assign n61490 = ~n64355;
  assign n64200 = ~n61492 | ~n64096;
  assign n63279 = n63276 & n63275;
  assign n74824 = ~n61450 | ~n61449;
  assign n61449 = ~n74285;
  assign n61450 = ~n74286;
  assign n74328 = ~n74326 | ~n74327;
  assign n62888 = n62897 | n63724;
  assign n63180 = ~n62973 | ~n62972;
  assign n61454 = ~n61462 | ~n60734;
  assign n71600 = ~n71603;
  assign n74368 = ~n74903 ^ n74904;
  assign n63657 = ~n63437 ^ n63908;
  assign n63437 = ~n63596 ^ n63597;
  assign n63447 = ~n63657 ^ n63658;
  assign n61017 = ~n71616;
  assign n74255 = ~n74393 ^ n61021;
  assign n61021 = ~n74391 ^ n71623;
  assign n63662 = n63447 | n63446;
  assign n63832 = ~n63666;
  assign n63373 = ~n63361 ^ n63300;
  assign n60875 = ~n60855 | ~n60854;
  assign n60854 = ~n63224;
  assign n60994 = ~n71646 | ~n71647;
  assign n71633 = ~n74255 ^ n74256;
  assign n74260 = n71633 | n71632;
  assign n61020 = ~n74393 ^ n74391;
  assign n74948 = ~n61463 | ~n74935;
  assign n61463 = ~n61464 | ~n61465;
  assign n61465 = ~n74397;
  assign n68948 = ~n61319 ^ n68786;
  assign n60945 = ~n61391 | ~n71663;
  assign n61477 = ~n71665 | ~n71664;
  assign n68958 = ~n60835 ^ n68959;
  assign n74445 = ~n61482 | ~n61481;
  assign n68982 = ~n61125 | ~n68981;
  assign n64484 = ~n61126 | ~n64340;
  assign n61126 = ~n61127 | ~n64130;
  assign n61127 = ~n64336 & ~n61128;
  assign n64128 = ~n64132 ^ n61124;
  assign n61124 = ~n64131;
  assign n63588 = ~n63385 | ~n63384;
  assign n63473 = ~n63676 | ~n63681;
  assign n63474 = ~n63677 ^ n63682;
  assign n61346 = ~n64659 ^ n60814;
  assign n61347 = ~n61345 | ~n64656;
  assign n61345 = ~n64652 | ~n64651;
  assign n76076 = n76028 & DIN_20_;
  assign n64109 = ~n64112 ^ n64110;
  assign n74738 = ~n74750 ^ n74749;
  assign n71186 = ~n61350 | ~n71672;
  assign n68992 = ~n67922 ^ n68974;
  assign n64328 = ~n64490;
  assign n64117 = ~n64325;
  assign n61445 = ~n74730;
  assign n60881 = ~n64036;
  assign n64576 = ~n74812 & ~n64573;
  assign n64361 = ~DIN_0_;
  assign n63888 = ~n63877 ^ n64022;
  assign n63877 = ~n64267 ^ n63870;
  assign n64592 = ~n64396 | ~n64395;
  assign n64395 = ~n61320 | ~n64394;
  assign n64396 = n64389 & n64388;
  assign n60947 = ~n60948 | ~n67274;
  assign n61484 = ~n67291 ^ n59901;
  assign n61250 = ~n61247 | ~n64601;
  assign n67250 = ~n64692 | ~n64691;
  assign n61360 = ~n64431;
  assign n63148 = ~n64032 | ~n71230;
  assign n63150 = P4_DATAO_REG_11__SCAN_IN & P4_DATAO_REG_12__SCAN_IN;
  assign n67841 = ~n60940 ^ n68836;
  assign n60940 = ~n70080 ^ n67835;
  assign n64677 = ~n74798 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n64081 = ~n64060 ^ n64059;
  assign n64059 = ~n64282;
  assign n64052 = ~n63882 | ~n63612;
  assign n63623 = ~n71230 & ~n74820;
  assign n71533 = ~n71257 | ~n71520;
  assign n68843 = ~n68845;
  assign n61262 = ~n67847 | ~n67846;
  assign n67848 = ~n61262 ^ n68886;
  assign n64432 = ~n64431 ^ n64430;
  assign n64224 = n64223 & n64306;
  assign n63980 = ~n63981 | ~n63982;
  assign n63417 = ~n63619 ^ n63613;
  assign n63163 = ~n63156;
  assign n63158 = ~n76045 & ~n63724;
  assign n62997 = ~n60852 | ~n62953;
  assign n60852 = ~n62989 ^ n63156;
  assign n70082 = ~n60740 | ~n60939;
  assign n60939 = ~n67835;
  assign n67330 = ~n76000 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n64437 = ~n64232 | ~n64231;
  assign n64304 = ~n64291 | ~n64290;
  assign n67862 = ~n61140 | ~n61246;
  assign n68915 = n70110 | n76000;
  assign n61263 = ~n68892;
  assign n71288 = ~n60991 ^ n71561;
  assign n60991 = ~n71549 ^ n71282;
  assign n74330 = ~n71544 ^ n74319;
  assign n61022 = ~n61023 & ~n74812;
  assign n64628 = n59930 & P4_DATAO_REG_10__SCAN_IN;
  assign n64447 = ~n76000 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n63981 = ~n63897 | ~n63898;
  assign n63905 = ~n61369 | ~n61368;
  assign n61369 = ~n63912;
  assign n63276 = ~n63144 | ~n63141;
  assign n74284 = ~n61470 ^ n74822;
  assign n74300 = ~n74841 ^ n74842;
  assign n71315 = ~n71310 | ~n70097;
  assign n62922 = ~n62926 | ~n62881;
  assign n67233 = n67228 | n67227;
  assign n67350 = n64350 & P4_DATAO_REG_8__SCAN_IN;
  assign n64756 = ~n64754 ^ n67342;
  assign n64754 = ~n64753 | ~n64752;
  assign n63649 = ~n76056 & ~n59984;
  assign n63174 = ~n63002 ^ n63144;
  assign n60847 = ~n63144;
  assign n70149 = ~n68943 ^ n70016;
  assign n60998 = ~n61000 | ~n60999;
  assign n74343 = ~n74346;
  assign n63603 = ~P4_DATAO_REG_16__SCAN_IN;
  assign n64546 = n63929 & P4_DATAO_REG_6__SCAN_IN;
  assign n60968 = ~n67243 | ~n61412;
  assign n64206 = n64205 & n64204;
  assign n61001 = ~n74261 ^ n61004;
  assign n61003 = ~n71595;
  assign n68787 = ~n68790 | ~n67750;
  assign n63923 = n59930 & P4_DATAO_REG_6__SCAN_IN;
  assign n63357 = ~n63365 | ~n63356;
  assign n63014 = ~n63181 | ~n61553;
  assign n63006 = n63181 | n63005;
  assign n60996 = ~n71359;
  assign n71361 = ~n71496 ^ n71497;
  assign n61458 = ~n61453 | ~n61459;
  assign n74376 = ~n61015 | ~n71609;
  assign n67890 = ~n76051 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n64156 = ~n64147;
  assign n74939 = ~n74260 | ~n74259;
  assign n70187 = ~n70186;
  assign n62909 = ~n63028 | ~n62904;
  assign n64671 = ~n64669;
  assign n61480 = ~n67221;
  assign n64316 = ~n64523 ^ n64525;
  assign n63956 = n64157 & n63954;
  assign n61133 = ~n63918 | ~n63664;
  assign n61343 = ~n61344 | ~n63459;
  assign n63022 = ~n63223 ^ n63224;
  assign n71660 = ~P4_DATAO_REG_6__SCAN_IN;
  assign n71658 = ~n71656 ^ n71655;
  assign n74976 = ~n60992 | ~n74435;
  assign n74395 = ~n61020 | ~n71623;
  assign n71388 = ~n71387;
  assign n63026 = ~n62911 ^ n62910;
  assign n64511 = n64513 | n60736;
  assign n60853 = ~n63221;
  assign n74447 = ~n74771 & ~n76063;
  assign n64506 = n64662 & n64505;
  assign n61138 = ~n61139 | ~n64641;
  assign n74221 = ~n61477 | ~n61476;
  assign n61476 = n71666 & n76055;
  assign n61373 = ~n68777 ^ n68776;
  assign n63574 = ~n63303 | ~n63302;
  assign n74219 = ~n74214 | ~n74213;
  assign n61241 = ~n74208 | ~n74207;
  assign n76038 = n76028 & DIN_25_;
  assign n67913 = ~n67366 ^ n61256;
  assign n61256 = ~n67916;
  assign n61348 = ~n64128;
  assign n61439 = ~n63587;
  assign n76061 = ~n76028 | ~DIN_16_;
  assign n63575 = ~n63379 | ~n63563;
  assign n63706 = ~n76028 | ~DIN_11_;
  assign n64837 = ~n100087 | ~n100136;
  assign n64835 = ~P1_P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~n65089;
  assign n76046 = n76028 & DIN_21_;
  assign n76043 = n76028 & DIN_19_;
  assign n61437 = ~n61346;
  assign n63931 = ~n64109;
  assign n75033 = ~n64827;
  assign n97746 = ~n65136;
  assign n67923 = ~n67734 ^ n60873;
  assign n60873 = ~n68992 ^ n67733;
  assign n68989 = ~n68984;
  assign n78645 = ~n64657 ^ n64658;
  assign n99992 = ~P1_P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P1_P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n96865 = ~n99992;
  assign n76802 = ~n64905 & ~n64904;
  assign n71174 = ~n69992 & ~n69991;
  assign n99201 = ~n65059 & ~n65058;
  assign n97648 = n62435 | n62434;
  assign n62435 = n62433 & n62432;
  assign n76224 = n97636 & n97648;
  assign n98061 = ~n97971;
  assign n97645 = ~n97648;
  assign n60728 = n61485 & n64351;
  assign n75006 = ~n61477 | ~n71666;
  assign n60862 = ~n75006;
  assign n60729 = n64287 & n60803;
  assign n60730 = n64092 & n64091;
  assign n60731 = n68982 & n60933;
  assign n61012 = ~n71609;
  assign n60734 = n74361 | n74360;
  assign n60736 = ~n63929 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n74820 = ~n59940;
  assign n74882 = ~P4_DATAO_REG_20__SCAN_IN;
  assign n60740 = n68836 ^ n70080;
  assign n61251 = ~n64601;
  assign n60747 = n74764 ^ n74444;
  assign n60878 = ~n64409;
  assign n64056 = n63889 & n64019;
  assign n61004 = ~n74262;
  assign n60750 = n63393 | n74846;
  assign n60752 = n67337 | n67336;
  assign n60759 = n74777 | n74776;
  assign n60761 = n63847 & n60210;
  assign n63885 = ~n74396 & ~n64572;
  assign n60762 = n64579 & n64693;
  assign n61162 = ~n64630;
  assign n60764 = n61255 & n64271;
  assign n75994 = ~P4_DATAO_REG_27__SCAN_IN;
  assign n64266 = ~n59940 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n60926 = ~n64266;
  assign n61395 = ~n70080;
  assign n60768 = n64287 & n64427;
  assign n60769 = n63419 & P4_DATAO_REG_11__SCAN_IN;
  assign n60773 = n64404 & n64405;
  assign n60774 = P4_DATAO_REG_27__SCAN_IN & P4_DATAO_REG_28__SCAN_IN;
  assign n60776 = ~n71371 | ~n71370;
  assign n60778 = ~n71360 | ~n71359;
  assign n63296 = n76028 & DIN_8_;
  assign n97204 = ~n98052;
  assign n60788 = n64837 | n64836;
  assign n60790 = n64835 | n64824;
  assign n60791 = n64835 | n99991;
  assign n60792 = n96865 | n99991;
  assign n60796 = n64837 | n100090;
  assign n60799 = n96865 | n64832;
  assign n60802 = n76056 | n74360;
  assign n61246 = ~n67861;
  assign n64536 = ~n76064 & ~n74367;
  assign n61160 = ~n63982;
  assign n64456 = ~n71660 & ~n74367;
  assign n61146 = ~n64456;
  assign n61460 = ~n60734;
  assign n60803 = P4_DATAO_REG_12__SCAN_IN & DIN_7_;
  assign n60805 = n74937 ^ n74950;
  assign n60806 = n74930 & P4_DATAO_REG_2__SCAN_IN;
  assign n60808 = n71660 | n76044;
  assign n60810 = n71659 & P4_DATAO_REG_3__SCAN_IN;
  assign n60811 = n74223 & P4_DATAO_REG_5__SCAN_IN;
  assign n60812 = ~n71659 | ~n76046;
  assign n60814 = n76076 & P4_DATAO_REG_1__SCAN_IN;
  assign n60933 = ~n69995;
  assign n60816 = n74465 | n74728;
  assign n60819 = ~n67324 ^ n67323;
  assign n61364 = ~n59858;
  assign n61142 = ~n61318 | ~n68969;
  assign n67884 = ~n68813;
  assign n61132 = ~n63662 | ~n63663;
  assign n68803 = ~n68802;
  assign n64397 = ~n64590 ^ n64566;
  assign n61163 = ~n64397 ^ n64592;
  assign n61144 = ~n61145 | ~n61148;
  assign n63638 = ~n61078 | ~n63425;
  assign n61078 = ~n61079 ^ n63635;
  assign n60834 = ~n61367 ^ n64165;
  assign n64147 = ~n61367 ^ n64165;
  assign n60835 = ~n67365 ^ n67364;
  assign n60836 = ~n67364 ^ n67365;
  assign n63066 = ~n63061 | ~n63060;
  assign n68804 = ~n68798 | ~n68799;
  assign n68801 = ~n68798;
  assign n60838 = ~n67345 ^ n61361;
  assign n64731 = ~n60839 | ~n64729;
  assign n61462 = ~n74790;
  assign n71572 = ~n71575;
  assign n74261 = ~n74269 | ~n71586;
  assign n60842 = ~n71256;
  assign n74793 = ~n61461 | ~n61460;
  assign n61151 = ~n67306;
  assign n64596 = n61163 | n64398;
  assign n71264 = ~n70052 | ~n71246;
  assign n70144 = ~n70143 ^ n71219;
  assign n70105 = ~n70104 | ~n70103;
  assign n60846 = ~n63260 | ~n63261;
  assign n63165 = n63167 | n63166;
  assign n63281 = ~n60848 | ~n63273;
  assign n60848 = ~n63272 | ~n63271;
  assign n61349 = ~n63312;
  assign n60851 = ~n64254 | ~n64255;
  assign n60855 = ~n63131 | ~n63132;
  assign n63143 = ~n63000 | ~n60856;
  assign n60857 = ~n62995;
  assign n61079 = ~n63636;
  assign n61492 = ~n61494 | ~n61493;
  assign n64352 = ~n64539 ^ n64351;
  assign n67225 = ~n67890 ^ n59967;
  assign n63828 = ~n63594 | ~n63593;
  assign n68878 = n68875 | n68874;
  assign n61094 = ~n64204;
  assign n61082 = ~n60859 | ~n60769;
  assign n60876 = ~n60860 | ~n60811;
  assign n60860 = ~n60640 | ~n76063;
  assign n60861 = ~n60862 | ~n60811;
  assign n64431 = ~n64429 | ~n64428;
  assign n68970 = ~n61142;
  assign n60865 = ~n74248 | ~n74231;
  assign n71325 = ~n71324 | ~n71323;
  assign n74391 = ~n71629 | ~n71622;
  assign n63970 = ~n63969 | ~n60871;
  assign n60871 = ~n63968 | ~n63980;
  assign n68797 = ~n60872 | ~n68789;
  assign n60872 = ~n68788 | ~n68787;
  assign n70195 = ~n70193 | ~n61366;
  assign n63199 = n63202 | n63070;
  assign n63827 = ~n63828 ^ n63829;
  assign n63810 = ~n63827 ^ n63674;
  assign n60874 = ~n70195;
  assign n63950 = ~n63810 | ~n63943;
  assign n63140 = ~n63135 | ~n60875;
  assign n64588 = ~n64581 | ~n64580;
  assign n71681 = ~n60882 | ~n74204;
  assign n71635 = ~n74960 ^ n71501;
  assign n75000 = ~n74788 ^ n76197;
  assign n68815 = ~n68824 | ~n68822;
  assign n64402 = ~n60879 | ~n60877;
  assign n60879 = ~n64400;
  assign n68824 = ~n60880 | ~n68810;
  assign n67761 = ~n67770 ^ n67771;
  assign n64044 = ~n60881 | ~n74361;
  assign n64776 = ~n64636 | ~n64635;
  assign n68884 = ~n61357 | ~n68883;
  assign n60938 = n67304 | n67303;
  assign n68819 = ~n68814 | ~n68813;
  assign n68813 = n67882 & n67883;
  assign n64366 = ~n64363 & ~n64364;
  assign n74208 = ~n74203 | ~n60889;
  assign n64801 = ~n68769 | ~n60716;
  assign n64415 = ~n60890 | ~n64407;
  assign n60890 = ~n64406 | ~n64410;
  assign n68775 = ~n60892 | ~n68777;
  assign n67911 = ~n61373 ^ n60892;
  assign n64024 = ~n60893 | ~n64020;
  assign n64028 = ~n64022 | ~n60926;
  assign n60925 = ~n64022 ^ n64266;
  assign n64269 = ~n64265 | ~n60893;
  assign n64296 = ~n64288 | ~n60768;
  assign n60894 = ~n60895;
  assign n64292 = ~n64288 | ~n60729;
  assign n64425 = ~n60895 | ~n64427;
  assign n64295 = ~n60895 | ~n60803;
  assign n64428 = ~n60894 | ~n64294;
  assign n61104 = ~n67358 ^ n60838;
  assign n64586 = ~n64582 | ~n60900;
  assign n64618 = ~n60908 | ~n64622;
  assign n64445 = ~n64304 | ~n60908;
  assign n64624 = ~n64623 | ~n60908;
  assign n64767 = ~n67348 | ~n60915;
  assign n67207 = ~n67205 | ~n61135;
  assign n71391 = ~n71482 ^ n71381;
  assign n64239 = ~n64238 | ~n60924;
  assign n64018 = ~n64267 ^ n60925;
  assign n63917 = ~n63915 ^ n63914;
  assign n69998 = ~n69997 | ~n60929;
  assign n61125 = ~n69997 ^ n60929;
  assign n68978 = ~n68977 ^ n60929;
  assign n60929 = ~n68972 ^ n61089;
  assign n60931 = ~n60932 | ~n64512;
  assign n60932 = ~n64511 | ~n64510;
  assign n60934 = ~n60731 | ~n69999;
  assign n61475 = ~n64441 | ~n60935;
  assign n64442 = n60935 | n64441;
  assign n60935 = ~n64434 ^ n64433;
  assign n64057 = ~n60936 | ~n64056;
  assign n67867 = ~n61245 ^ n67860;
  assign n70118 = n70107 | n60937;
  assign n67306 = ~n67305 | ~n60938;
  assign n68836 = ~n68875 ^ n68873;
  assign n60943 = ~n74240;
  assign n60946 = ~n60942 | ~n60941;
  assign n60941 = ~n74240 | ~n60812;
  assign n60942 = ~n60943 | ~n71659;
  assign n60944 = ~n60946 | ~n60945;
  assign n67241 = ~n60968 | ~n67239;
  assign n67354 = ~n60968 ^ n67242;
  assign n60984 = ~n71263;
  assign n60985 = ~n60986;
  assign n71516 = ~n60986 | ~n71263;
  assign n71256 = ~n71253 | ~n60987;
  assign n60987 = n71254 & n71252;
  assign n60992 = ~n74430 | ~n60993;
  assign n60993 = ~n74431;
  assign n74407 = ~n60997 ^ n74948;
  assign n60997 = ~n74939 ^ n60805;
  assign n74832 = n60998 & n74292;
  assign n60999 = ~n71531;
  assign n61000 = ~n71530;
  assign n74265 = ~n61001 | ~n61003;
  assign n61008 = ~n61006 | ~n61005;
  assign n61005 = n74374 | n71609;
  assign n61006 = ~n74374 | ~n71609;
  assign n61014 = ~n74373;
  assign n61016 = ~n71615;
  assign n61010 = ~n61013 | ~n61011;
  assign n61011 = n74374 | n61012;
  assign n61013 = ~n74374 | ~n61012;
  assign n61015 = ~n74373 ^ n74374;
  assign n74380 = ~n61017 | ~n61016;
  assign n71524 = ~n71523 | ~n61022;
  assign n71547 = ~n71545 | ~n71546;
  assign n71506 = ~n71281 | ~n71280;
  assign n74456 = ~n61036 | ~n71473;
  assign n71401 = ~n71395 | ~n61036;
  assign n61036 = ~n61410 | ~n71394;
  assign n67771 = ~n67327;
  assign n61039 = n67331 & n60752;
  assign n64603 = ~n64600 | ~n61065;
  assign n61065 = ~n61248 | ~n61250;
  assign n64752 = ~n61075 | ~n61522;
  assign n64743 = ~n61075 | ~n67338;
  assign n61080 = ~n59923 | ~n60769;
  assign n61081 = ~n59923 | ~n74820;
  assign n70193 = ~n61089 | ~n70192;
  assign n61371 = n61090 & n64347;
  assign n61093 = ~n64794 ^ n64793;
  assign n67213 = ~n61093;
  assign n67212 = ~n67206 | ~n61093;
  assign n61441 = ~n64799 ^ n61093;
  assign n64198 = ~n61094 | ~n64195;
  assign n64636 = ~n60728 | ~n61095;
  assign n68791 = n61104 | n67751;
  assign n68790 = ~n61104 | ~n67751;
  assign n67889 = ~n67359 ^ n61104;
  assign n61128 = ~n64129;
  assign n61129 = ~n63432 | ~n61130;
  assign n67921 = ~n61131 | ~n67913;
  assign n68984 = ~n61131 ^ n67913;
  assign n61134 = ~n61132 | ~n63661;
  assign n64797 = ~n64795 | ~n61135;
  assign n61136 = ~n63355 | ~n63363;
  assign n63594 = n61137 | n63590;
  assign n63677 = ~n61137 ^ n63468;
  assign n61139 = ~n64643;
  assign n67859 = ~n61141 | ~n67861;
  assign n61140 = ~n61141;
  assign n61245 = ~n61141 ^ n61246;
  assign n63334 = ~n63247;
  assign n64459 = ~n61442 | ~n61144;
  assign n67829 = ~n67289 | ~n67264;
  assign n61152 = ~n67307;
  assign n61158 = ~n63974;
  assign n64005 = ~n61159 | ~n63968;
  assign n63903 = ~n63968 ^ n61160;
  assign n64399 = ~n61163 | ~n64398;
  assign n61166 = ~n67325 | ~n61244;
  assign n74217 = ~n74216 | ~n61241;
  assign n74209 = ~n61241;
  assign n74743 = n74734 & n61241;
  assign n61242 = n67325 | n61244;
  assign n61244 = ~n67323;
  assign n64735 = ~n67325;
  assign n61248 = ~n61249 | ~n64405;
  assign n64357 = ~n61252 | ~n64237;
  assign n61252 = ~n64082 | ~n64081;
  assign n61253 = ~n68778 & ~n60810;
  assign n61254 = ~n68778;
  assign n64026 = ~n60764 | ~n64029;
  assign n61258 = ~n71283 ^ n71284;
  assign n71287 = ~n61258 | ~n70072;
  assign n71582 = ~n61260 | ~n71581;
  assign n71675 = ~n71672 | ~n71671;
  assign n61440 = ~n71672 ^ n71671;
  assign n68888 = ~n61262 | ~n68887;
  assign n70108 = ~n68893 ^ n61263;
  assign n68893 = ~n68895 ^ n68894;
  assign n64720 = ~n60762 | ~n61496;
  assign n64695 = ~n61496 | ~n64579;
  assign n71371 = ~n70185 ^ n61319;
  assign n64616 = ~n61321 ^ n64560;
  assign n64737 = ~n61321 ^ n59961;
  assign n61321 = ~n64558 | ~n64559;
  assign n61324 = ~n68787 | ~n68791;
  assign n63668 = ~n63670 ^ n63669;
  assign n63313 = ~n63270 ^ n63269;
  assign n61358 = ~n61384 ^ n70135;
  assign n64556 = ~n60832 | ~n64431;
  assign n64558 = ~n61360 | ~n64557;
  assign n61363 = ~n61364 | ~n63610;
  assign n63404 = ~n61365 | ~n63343;
  assign n68972 = ~n61366 | ~n70192;
  assign n61368 = ~n61370;
  assign n63915 = ~n61370 ^ n63912;
  assign n64289 = ~n64357 ^ n64359;
  assign n68777 = ~n67910 ^ n61479;
  assign n61384 = ~n70128 ^ n68924;
  assign n61388 = ~n74232;
  assign n61391 = ~n61388 | ~n60808;
  assign n61392 = ~n61394 | ~n61393;
  assign n71474 = n71190 & n71189;
  assign n67753 = ~n61412 | ~n67344;
  assign n67244 = n61412 & n67242;
  assign n67368 = ~n61435 | ~n67374;
  assign n64657 = ~n61347 ^ n61437;
  assign n61438 = ~n63447 | ~n63446;
  assign n63803 = ~n63796 | ~n63799;
  assign n64478 = ~n64476 | ~n61447;
  assign n61447 = ~n64527 | ~n71345;
  assign n63899 = ~n63897;
  assign n74787 = ~n61448 | ~n74782;
  assign n75001 = ~n61448 ^ n74765;
  assign n61448 = ~n74764 ^ n74776;
  assign n74915 = ~n74920;
  assign n74932 = ~n74390 | ~n61451;
  assign n61451 = ~n74920 | ~n74389;
  assign n61456 = ~n61454 | ~n61453;
  assign n61453 = ~n74790 | ~n61460;
  assign n61461 = ~n74789 ^ n74790;
  assign n61457 = ~n74789 | ~n61458;
  assign n61459 = ~n61462 | ~n60734;
  assign n74404 = ~n74407;
  assign n61464 = ~n74398;
  assign n61471 = ~n74333 | ~n74334;
  assign n74841 = ~n74834 | ~n61472;
  assign n61472 = ~n74293 | ~n74294;
  assign n64766 = ~n67354 | ~n60720;
  assign n61473 = n63415 | n63414;
  assign n64630 = ~n64442 | ~n61475;
  assign n61478 = ~n74450;
  assign n68964 = n61479 | n68956;
  assign n64791 = ~n67220 ^ n61480;
  assign n67220 = n64790 & n64789;
  assign n61481 = ~n74447;
  assign n61482 = ~n59867;
  assign n74448 = ~n59867 | ~n74447;
  assign n71668 = ~n61483 ^ n74447;
  assign n61486 = ~n60091;
  assign n61488 = ~n64349;
  assign n61493 = ~n64090 | ~n60730;
  assign n61494 = ~n64093;
  assign n64093 = ~n63902 ^ n63903;
  assign n64580 = ~n61496 | ~n61495;
  assign n63902 = ~n61159 ^ n63901;
  assign n74240 = n71658 | n71657;
  assign n67240 = ~n67351;
  assign n63611 = ~n63886 ^ n63878;
  assign n64718 = ~n74276 | ~n64570;
  assign n64225 = ~n64220 | ~n64221;
  assign n64218 = n64220 | n64006;
  assign n67362 = ~n67744 | ~n67741;
  assign n63896 = ~n64068 ^ n64066;
  assign n61511 = n63853 & n74835;
  assign n61519 = ~n70189 | ~n70188;
  assign n61522 = P4_DATAO_REG_11__SCAN_IN & DIN_11_;
  assign n71345 = ~n63929;
  assign n68776 = n76046 & P4_DATAO_REG_3__SCAN_IN;
  assign n61528 = n63950 & n63944;
  assign n61534 = n63799 & n59980;
  assign n61535 = n74763 | n76061;
  assign n68816 = ~n76056 & ~n76061;
  assign n64015 = ~n64065;
  assign n61549 = P4_DATAO_REG_13__SCAN_IN & P4_DATAO_REG_12__SCAN_IN;
  assign n61551 = n63914 ^ n63916;
  assign n64528 = ~n64526;
  assign n61553 = n63178 | n74846;
  assign n97723 = n97928 & n97620;
  assign n61554 = P4_DATAO_REG_10__SCAN_IN & P4_DATAO_REG_9__SCAN_IN;
  assign n61555 = P4_DATAO_REG_7__SCAN_IN & P4_DATAO_REG_8__SCAN_IN;
  assign n76028 = ~n60904;
  assign n62954 = ~n64572;
  assign n61571 = ~n63874 | ~n63873;
  assign n61573 = ~n63808 | ~n63807;
  assign n63796 = ~n63798;
  assign n61574 = n74975 & n74974;
  assign n61575 = ~n71484 | ~n71483;
  assign n64261 = DIN_1_ & P4_DATAO_REG_17__SCAN_IN;
  assign n68856 = ~n74276 | ~n64704;
  assign n64380 = ~n64392;
  assign n64255 = ~n64246 | ~n64245;
  assign n64589 = ~n64566;
  assign n63607 = P4_DATAO_REG_15__SCAN_IN & P4_DATAO_REG_16__SCAN_IN;
  assign n68852 = ~n70053 ^ n70054;
  assign n64074 = ~n64068;
  assign n71279 = ~P4_DATAO_REG_21__SCAN_IN;
  assign n67840 = ~n67841;
  assign n68880 = ~n70074 ^ n68879;
  assign n71293 = ~P4_DATAO_REG_18__SCAN_IN;
  assign n64061 = ~n64081;
  assign n64221 = ~n64008 | ~n64007;
  assign n63402 = n63395 & P4_DATAO_REG_9__SCAN_IN;
  assign n74353 = ~P4_DATAO_REG_19__SCAN_IN;
  assign n64443 = ~n64435;
  assign n67872 = ~n68918;
  assign n68935 = ~n68939;
  assign n63653 = ~n63651;
  assign n67878 = ~n68810 | ~n68809;
  assign n63907 = ~n63596;
  assign n70170 = n70163 & n70162;
  assign n63444 = n63443 | n63442;
  assign n68944 = ~n70149;
  assign n63663 = n63660 | n63659;
  assign n71501 = ~n74409 ^ n74962;
  assign n68781 = ~n68780;
  assign n64473 = ~n64527 ^ n63929;
  assign n64173 = ~n64164;
  assign n63466 = ~n63460 | ~n63461;
  assign n76081 = ~P4_DATAO_REG_5__SCAN_IN;
  assign n63671 = n63670 | n63669;
  assign n63023 = ~n63022 | ~n63021;
  assign n63468 = ~n63590;
  assign n63308 = n63307 | n74881;
  assign n63221 = ~n63196 ^ n63230;
  assign n74245 = ~n74244 | ~n74243;
  assign n74982 = ~n74981 | ~n74980;
  assign n63382 = n63381 & n63380;
  assign n63808 = ~n61534 | ~n63796;
  assign n76056 = ~P4_DATAO_REG_8__SCAN_IN;
  assign n68778 = n68777 & n68776;
  assign n64642 = ~n64641;
  assign n74788 = ~n75921 ^ n74781;
  assign n74771 = ~P4_DATAO_REG_4__SCAN_IN;
  assign n63929 = n76028 & DIN_15_;
  assign n64491 = ~n64327 | ~n64326;
  assign n71398 = ~n71400;
  assign n74780 = ~n76055;
  assign n68979 = ~n67911 | ~n67912;
  assign n74930 = ~n76061;
  assign n71181 = n71180 | n71179;
  assign n67379 = n67373 & n67372;
  assign n64651 = ~n64494 | ~n64493;
  assign n75055 = ~n60791;
  assign n97761 = ~n60792;
  assign n97225 = ~n60796;
  assign n63775 = n63774 | n63773;
  assign n71469 = ~n71410 | ~n71409;
  assign n99178 = ~n99179 & ~n96896;
  assign n100130 = ~n65079 & ~n65078;
  assign n70255 = n63789 & n63788;
  assign n62410 = P1_P1_ADDRESS_REG_25__SCAN_IN | P1_P1_ADDRESS_REG_24__SCAN_IN;
  assign n99199 = ~n65119 & ~n65118;
  assign n97747 = ~n64817;
  assign n74470 = n63776 & n63775;
  assign n71419 = n63767 & n63766;
  assign n71693 = ~n71412 ^ n74212;
  assign n75022 = n63780 & n63779;
  assign n99221 = ~n64935 | ~n64934;
  assign n99213 = ~n97620 & ~n100066;
  assign n100048 = ~n65110 & ~n65118;
  assign n97895 = ~n97866;
  assign n70278 = ~P1_P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n96896 = ~n99221;
  assign n99179 = n64997 & n64996;
  assign n97620 = ~n97556;
  assign n97930 = ~n98024;
  assign n100479 = ~n100184 & ~n96193;
  assign n96895 = ~n99179;
  assign n97928 = ~n100164 & ~n65125;
  assign n99180 = ~n64875 & ~n64874;
  assign n100164 = ~n100479;
  assign n62434 = ~P1_P1_ADDRESS_REG_29__SCAN_IN;
  assign n96899 = ~n65029 & ~n65028;
  assign n97556 = ~n64845 & ~n64844;
  assign n97636 = n97723 & n96895;
  assign n97929 = ~n97723;
  assign n97971 = n97928 & n65126;
  assign n100044 = ~P1_P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n62412 = ~P1_P1_ADDRESS_REG_27__SCAN_IN & ~P1_P1_ADDRESS_REG_26__SCAN_IN;
  assign n62408 = ~P1_P1_ADDRESS_REG_23__SCAN_IN & ~P1_P1_ADDRESS_REG_22__SCAN_IN;
  assign n62407 = ~P1_P1_ADDRESS_REG_21__SCAN_IN & ~P1_P1_ADDRESS_REG_20__SCAN_IN;
  assign n62409 = ~n62408 | ~n62407;
  assign n62411 = ~n62410 & ~n62409;
  assign n62428 = ~n62412 | ~n62411;
  assign n62414 = ~P1_P1_ADDRESS_REG_15__SCAN_IN & ~P1_P1_ADDRESS_REG_14__SCAN_IN;
  assign n62413 = ~P1_P1_ADDRESS_REG_13__SCAN_IN & ~P1_P1_ADDRESS_REG_12__SCAN_IN;
  assign n62418 = ~n62414 | ~n62413;
  assign n62416 = ~P1_P1_ADDRESS_REG_19__SCAN_IN & ~P1_P1_ADDRESS_REG_18__SCAN_IN;
  assign n62415 = ~P1_P1_ADDRESS_REG_17__SCAN_IN & ~P1_P1_ADDRESS_REG_16__SCAN_IN;
  assign n62417 = ~n62416 | ~n62415;
  assign n62426 = ~n62418 & ~n62417;
  assign n62420 = ~P1_P1_ADDRESS_REG_7__SCAN_IN & ~P1_P1_ADDRESS_REG_6__SCAN_IN;
  assign n62419 = ~P1_P1_ADDRESS_REG_5__SCAN_IN & ~P1_P1_ADDRESS_REG_4__SCAN_IN;
  assign n62424 = ~n62420 | ~n62419;
  assign n62422 = ~P1_P1_ADDRESS_REG_11__SCAN_IN & ~P1_P1_ADDRESS_REG_10__SCAN_IN;
  assign n62421 = ~P1_P1_ADDRESS_REG_9__SCAN_IN & ~P1_P1_ADDRESS_REG_8__SCAN_IN;
  assign n62423 = ~n62422 | ~n62421;
  assign n62425 = ~n62424 & ~n62423;
  assign n62427 = ~n62426 | ~n62425;
  assign n62433 = ~n62428 & ~n62427;
  assign n62430 = ~P1_P1_ADDRESS_REG_0__SCAN_IN & ~P1_P1_ADDRESS_REG_28__SCAN_IN;
  assign n62429 = ~P1_P1_ADDRESS_REG_2__SCAN_IN & ~P1_P1_ADDRESS_REG_1__SCAN_IN;
  assign n62431 = ~n62430 | ~n62429;
  assign n62432 = ~n62431 & ~P1_P1_ADDRESS_REG_3__SCAN_IN;
  assign n74276 = n71248 & SEL;
  assign n62926 = ~n62942;
  assign n62880 = ~n64701 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n64259 = SEL & DIN_1_;
  assign n62881 = ~n62880 | ~n62879;
  assign n62921 = ~n59870 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n62882 = ~P4_DATAO_REG_7__SCAN_IN | ~P4_DATAO_REG_6__SCAN_IN;
  assign n62884 = ~n62883 | ~n76064;
  assign n62885 = P4_DATAO_REG_6__SCAN_IN & P4_DATAO_REG_5__SCAN_IN;
  assign n62897 = ~n74276 | ~n62885;
  assign n62886 = ~n59870 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n62887 = ~n62897 | ~n62886;
  assign n62892 = ~n62888 | ~n62887;
  assign n62890 = ~n62893 & ~n62892;
  assign n62889 = ~n62888;
  assign n62914 = ~n76081 & ~n74820;
  assign n62891 = ~n62914;
  assign n62907 = ~n62893 ^ n62892;
  assign n62895 = ~n64701 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n62894 = ~n71521 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n62896 = ~n62895 | ~n62894;
  assign n63029 = n62897 & n62896;
  assign n62898 = P4_DATAO_REG_5__SCAN_IN & P4_DATAO_REG_4__SCAN_IN;
  assign n63040 = ~n74276 | ~n62898;
  assign n62901 = n63040 | n60722;
  assign n62899 = ~n74771 & ~n64706;
  assign n62900 = ~n63040 | ~n62899;
  assign n63031 = ~n62901 | ~n62900;
  assign n62903 = ~n63029 | ~n63031;
  assign n62902 = n63040 | n63724;
  assign n62905 = ~n62903 | ~n62902;
  assign n63028 = ~n62907 ^ n62905;
  assign n63027 = ~n62954 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n62904 = ~n63027;
  assign n62906 = ~n62905;
  assign n62908 = n62907 | n62906;
  assign n62910 = ~n62909 | ~n62908;
  assign n63024 = ~n59905 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n62912 = ~n62911 | ~n62910;
  assign n62939 = ~n62913 | ~n62912;
  assign n62916 = ~n62915;
  assign n62923 = n62922 | n62921;
  assign n62957 = ~n62924 | ~n62923;
  assign n62944 = ~n60722 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n62925 = ~n62944;
  assign n62932 = ~n62926 ^ n62925;
  assign n62927 = ~n74276;
  assign n62948 = ~n62927;
  assign n62989 = ~n62948 | ~n62928;
  assign n62930 = ~n64701 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n62929 = ~n60375 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n62931 = ~n62930 | ~n62929;
  assign n62945 = ~n62989 | ~n62931;
  assign n62956 = ~n62932 ^ n62945;
  assign n62960 = ~n62957 ^ n62956;
  assign n62961 = ~n62954 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n62967 = ~n76081 & ~n59912;
  assign n62933 = ~n62967;
  assign n62934 = ~n62961 ^ n62933;
  assign n62935 = ~n62960 ^ n62934;
  assign n62938 = ~n62970 ^ n62935;
  assign n63057 = ~n74835 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n62936 = ~n63057;
  assign n62941 = ~n62937 | ~n62936;
  assign n62940 = ~n62939 | ~n62938;
  assign n62976 = ~n62941 | ~n62940;
  assign n63005 = n76028 & DIN_6_;
  assign n62974 = ~n63005 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63064 = ~n62976 ^ n62974;
  assign n62943 = ~n62945 | ~n62944;
  assign n62947 = ~n62943 | ~n62942;
  assign n62946 = n62945 | n62944;
  assign n62949 = ~n76045 | ~n74277;
  assign n62952 = ~n59991 | ~n62949;
  assign n62950 = ~n76045 & ~n63317;
  assign n62951 = ~n62950 & ~P4_DATAO_REG_10__SCAN_IN;
  assign n62953 = ~n62952 & ~n62951;
  assign n62996 = ~n59870 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n62998 = ~n59940 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n62955 = ~n62996 ^ n62998;
  assign n62982 = ~n59908 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n62980 = ~n62981 ^ n62982;
  assign n62959 = ~n62980;
  assign n62958 = ~n62957 | ~n62956;
  assign n63181 = ~n62959 ^ n62979;
  assign n62963 = ~n62960;
  assign n62962 = ~n62961;
  assign n62969 = ~n62965 | ~n62964;
  assign n62968 = ~n62966 | ~n62969;
  assign n62973 = ~n62968 | ~n62967;
  assign n62971 = ~n62969;
  assign n62972 = ~n62971 | ~n62970;
  assign n63179 = ~n63181 ^ n63180;
  assign n63188 = ~n63179;
  assign n63178 = ~n74835 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n63062 = ~n63188 ^ n63178;
  assign n62978 = ~n63064 | ~n63062;
  assign n62975 = ~n62974;
  assign n62977 = ~n62976 | ~n62975;
  assign n63224 = ~n62978 | ~n62977;
  assign n62985 = ~n62980 | ~n62979;
  assign n62983 = ~n62981;
  assign n63175 = ~n62985 | ~n62984;
  assign n63166 = ~n76056 & ~n74820;
  assign n62987 = ~n63166;
  assign n62988 = ~n63156 ^ n62987;
  assign n62993 = ~n63162 ^ n62988;
  assign n62992 = n62997 | n62996;
  assign n62990 = ~n62989;
  assign n62991 = ~n62990 | ~n63156;
  assign n63164 = ~n62992 | ~n62991;
  assign n62999 = ~n62997 ^ n62996;
  assign n63142 = ~n76064 & ~n59912;
  assign n63001 = ~n63142;
  assign n63002 = ~n63143 ^ n63001;
  assign n63003 = ~n74835 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n63004 = ~n63287 | ~n63003;
  assign n63020 = ~n63186;
  assign n63395 = ~n63855 | ~n74846;
  assign n63011 = n63395 & P4_DATAO_REG_5__SCAN_IN;
  assign n63008 = ~n63006 | ~n63011;
  assign n63007 = ~n63180;
  assign n63018 = n63008 & n63007;
  assign n63182 = ~n63005 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n63190 = ~n63182;
  assign n63010 = n63180 & n63190;
  assign n63009 = n63181 | n74835;
  assign n63016 = ~n63010 | ~n63009;
  assign n63012 = ~n63011;
  assign n63013 = n63181 | n63012;
  assign n63015 = ~n63014 | ~n63013;
  assign n63017 = ~n63016 | ~n63015;
  assign n63021 = ~n74771 & ~n59984;
  assign n63227 = n63022 | n63021;
  assign n63197 = ~n63296 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63204 = ~n63197;
  assign n63025 = ~n63024;
  assign n63053 = ~n63026 ^ n63025;
  assign n63049 = ~n63028 ^ n63027;
  assign n63030 = ~n63029;
  assign n63045 = ~n63031 ^ n63030;
  assign n63032 = P4_DATAO_REG_4__SCAN_IN & P4_DATAO_REG_3__SCAN_IN;
  assign n63080 = ~n62948 | ~n63032;
  assign n63034 = ~n64701 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n63033 = ~n60375 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63035 = ~n63034 | ~n63033;
  assign n63037 = ~n63080 | ~n63035;
  assign n63036 = ~n63040;
  assign n63038 = n63040 | n63080;
  assign n63074 = ~n74763 & ~n63724;
  assign n63043 = ~n63076 | ~n63074;
  assign n63041 = ~n63080;
  assign n63042 = ~n63041 | ~n63040;
  assign n63044 = ~n63043 | ~n63042;
  assign n63090 = ~n63045 ^ n63044;
  assign n63089 = ~n62954 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63047 = n63090 | n63089;
  assign n63046 = ~n63045 | ~n63044;
  assign n63048 = ~n63047 | ~n63046;
  assign n63099 = ~n63049 ^ n63048;
  assign n63098 = ~n59906 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63051 = n63099 | n63098;
  assign n63050 = ~n63049 | ~n63048;
  assign n63052 = ~n63051 | ~n63050;
  assign n63104 = ~n63053 ^ n63052;
  assign n63103 = ~n74835 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63054 = ~n63053 | ~n63052;
  assign n63058 = ~n63055 | ~n63054;
  assign n63059 = ~n62937 ^ n63057;
  assign n63071 = ~n63058 ^ n63059;
  assign n63072 = ~n63005 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63061 = n63071 | n63072;
  assign n63060 = ~n63059 | ~n63058;
  assign n63063 = ~n63062;
  assign n63067 = ~n63064 ^ n63063;
  assign n63065 = ~n63202;
  assign n63070 = ~n74315 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63203 = ~n63067 | ~n63066;
  assign n63068 = ~n63199 | ~n63203;
  assign n63482 = ~n63065 ^ n63070;
  assign n63073 = ~n63071;
  assign n63075 = ~n63074;
  assign n63087 = ~n63076 ^ n63075;
  assign n63078 = ~n63504 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63079 = ~n63078 | ~n63077;
  assign n63083 = ~n63080 | ~n63079;
  assign n63082 = ~n60722 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63511 = ~n63083 ^ n63082;
  assign n63081 = P4_DATAO_REG_3__SCAN_IN & P4_DATAO_REG_2__SCAN_IN;
  assign n63502 = ~n62948 | ~n63081;
  assign n63085 = n63511 | n63502;
  assign n63084 = n63083 | n63082;
  assign n63086 = ~n63085 | ~n63084;
  assign n63516 = ~n63087 ^ n63086;
  assign n63517 = ~n62954 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63088 = ~n63087 | ~n63086;
  assign n63091 = ~n63090 ^ n63089;
  assign n63096 = ~n63092 | ~n63091;
  assign n63094 = ~n63091;
  assign n63095 = ~n63094 | ~n63093;
  assign n63497 = ~n63096 | ~n63095;
  assign n63496 = ~n71397 & ~n59912;
  assign n63101 = ~n63097 | ~n63096;
  assign n63100 = ~n63099 ^ n63098;
  assign n63490 = ~n63101 ^ n63100;
  assign n63491 = ~n74835 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63102 = n63101 | n63100;
  assign n63108 = ~n63495 | ~n63102;
  assign n63107 = ~n71397 & ~n74846;
  assign n63489 = ~n63104 ^ n63103;
  assign n63105 = ~n63489;
  assign n63110 = ~n63106 | ~n63105;
  assign n63109 = ~n63108 | ~n63107;
  assign n63486 = ~n74315 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63114 = ~n63111;
  assign n63113 = ~n63112;
  assign n63481 = ~n63296 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63115 = n63483 & n63481;
  assign n63116 = ~n63488 | ~n63115;
  assign n63122 = ~n63482 | ~n63116;
  assign n63119 = ~n63483 | ~n59984;
  assign n63118 = ~n63481;
  assign n63120 = n63119 & n63118;
  assign n63123 = ~n63122 | ~n63121;
  assign n63548 = ~n63124 ^ n63123;
  assign n63549 = ~n74798 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63553 = n63548 | n63549;
  assign n63125 = ~n63124 | ~n63123;
  assign n63127 = ~n63129;
  assign n63128 = ~n71397 & ~n74881;
  assign n63126 = ~n63128;
  assign n63130 = ~n63127 | ~n63126;
  assign n63212 = ~n63129 | ~n63128;
  assign n63136 = ~n63223;
  assign n63131 = ~n63136 | ~n60217;
  assign n63838 = ~n60217 | ~n59984;
  assign n63132 = n63838 & P4_DATAO_REG_4__SCAN_IN;
  assign n63843 = ~n60217 & ~n59984;
  assign n63133 = ~n63136 | ~n63132;
  assign n63135 = ~n63134 | ~n63133;
  assign n63137 = ~n63136 | ~n59984;
  assign n63138 = n63137 & n63296;
  assign n63141 = ~n63143;
  assign n63271 = ~n63276 | ~n63142;
  assign n63145 = ~n63271 | ~n63277;
  assign n63274 = ~n74835 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n63172 = ~n63145 ^ n63274;
  assign n63146 = ~P4_DATAO_REG_11__SCAN_IN | ~DIN_1_;
  assign n63147 = ~n64051 | ~n63146;
  assign n63149 = ~n63148 | ~n63147;
  assign n63151 = ~n74812 & ~n63149;
  assign n63241 = ~n74276 | ~n63150;
  assign n63244 = ~n63151 | ~n63241;
  assign n63243 = ~n59870 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n63153 = ~n63244 ^ n63243;
  assign n63154 = ~n63153 | ~n63152;
  assign n63252 = ~n62954 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n63266 = ~n59907 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n63155 = ~n63252 ^ n63266;
  assign n63161 = ~n63263 ^ n63155;
  assign n63159 = ~n63157;
  assign n63251 = ~n63159 | ~n63158;
  assign n63265 = ~n63160 | ~n63251;
  assign n63261 = ~n63161 ^ n63265;
  assign n63170 = ~n63261;
  assign n63169 = ~n63165 | ~n63164;
  assign n63168 = ~n63167 | ~n63166;
  assign n63260 = ~n63169 | ~n63168;
  assign n63273 = ~n63170 ^ n63260;
  assign n63171 = ~n63273;
  assign n63285 = ~n63172 ^ n63171;
  assign n63173 = ~n63285;
  assign n63289 = ~n63005 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n63177 = ~n63173 ^ n63289;
  assign n63288 = ~n63175 | ~n63174;
  assign n63176 = ~n63284 | ~n63288;
  assign n63233 = ~n63177 ^ n63176;
  assign n63184 = n63179 | n63178;
  assign n63189 = ~n63181 | ~n63180;
  assign n63183 = n63189 & n63182;
  assign n63185 = ~n63184 | ~n63183;
  assign n63195 = ~n63186 | ~n63185;
  assign n63187 = ~n63189;
  assign n63193 = n63188 | n63187;
  assign n63191 = ~n63189 | ~n63855;
  assign n63192 = n63191 & n63190;
  assign n63194 = ~n63193 | ~n63192;
  assign n63232 = ~n63195 | ~n63194;
  assign n63231 = ~n63233 ^ n63232;
  assign n63196 = ~n63231;
  assign n63230 = ~n74315 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n63198 = n63203 & n63197;
  assign n63201 = ~n63199 | ~n63198;
  assign n63209 = ~n63201 | ~n63200;
  assign n63207 = ~n63202 | ~n63203;
  assign n63205 = ~n63203 | ~n59984;
  assign n63206 = n63205 & n63204;
  assign n63208 = ~n63207 | ~n63206;
  assign n63217 = ~n63209 | ~n63208;
  assign n63215 = ~n63216 ^ n63217;
  assign n63211 = ~n63215;
  assign n63214 = ~n74763 & ~n76012;
  assign n63210 = ~n63214;
  assign n63479 = ~n63211 ^ n63210;
  assign n63213 = ~n63478 | ~n63479;
  assign n63218 = n63217 | n63216;
  assign n63307 = ~n63219 | ~n63218;
  assign n63220 = ~n76000 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63306 = ~n63307 ^ n63220;
  assign n63225 = n63224 | n63223;
  assign n63228 = ~n63227 | ~n63226;
  assign n63235 = n63231 | n63230;
  assign n63234 = ~n63233 | ~n63232;
  assign n63361 = ~n63235 | ~n63234;
  assign n63238 = ~n64051 | ~n64032;
  assign n63236 = ~DIN_1_ | ~P4_DATAO_REG_12__SCAN_IN;
  assign n63237 = ~n74396 | ~n63236;
  assign n63239 = ~n63238 | ~n63237;
  assign n63240 = ~n74812 & ~n63239;
  assign n63328 = ~n60722 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n63242 = ~n63241;
  assign n63245 = n63244 | n63243;
  assign n63333 = ~n62954 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n63339 = ~n63333;
  assign n63341 = ~n59908 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n63248 = ~n63339 ^ n63341;
  assign n63249 = ~n63263 | ~n63252;
  assign n63250 = n63251 & n63252;
  assign n63253 = ~n63251;
  assign n63262 = ~n63252;
  assign n63254 = ~n63253 | ~n63262;
  assign n63256 = ~n63255 | ~n63254;
  assign n63346 = ~n63258 | ~n63257;
  assign n63348 = ~n76056 & ~n63855;
  assign n63259 = ~n63348;
  assign n63264 = ~n63263 ^ n63262;
  assign n63267 = ~n63265 ^ n63264;
  assign n63269 = ~n63350;
  assign n63272 = n63277 & n63274;
  assign n63275 = ~n63274;
  assign n63278 = ~n63277 | ~n59912;
  assign n63280 = ~n63279 | ~n63278;
  assign n63312 = ~n63281 | ~n63280;
  assign n63310 = ~n63005 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n63299 = ~n63365;
  assign n63283 = n63288 & n63289;
  assign n63286 = ~n63284 | ~n63283;
  assign n63295 = ~n63286 | ~n63285;
  assign n63293 = ~n63287 | ~n63288;
  assign n63291 = ~n63288 | ~n63855;
  assign n63290 = ~n63289;
  assign n63294 = ~n63293 | ~n63292;
  assign n63356 = ~n71660 & ~n59984;
  assign n63362 = ~n63356;
  assign n63366 = ~n63296 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n63297 = ~n63362 ^ n63366;
  assign n63298 = ~n63363 ^ n63297;
  assign n63360 = ~n63299 ^ n63298;
  assign n63300 = ~n63360;
  assign n63372 = ~n74798 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63305 = ~n63460 ^ n63372;
  assign n63301 = ~n63306 ^ n63305;
  assign n63379 = ~n63303 ^ n63301;
  assign n63563 = n59930 & P4_DATAO_REG_2__SCAN_IN;
  assign n63302 = ~n63301;
  assign n63572 = ~n76054 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63304 = n63574 & n63572;
  assign n63378 = ~n63575 | ~n63304;
  assign n63309 = n63306 | n63305;
  assign n63472 = ~n63309 | ~n63308;
  assign n63311 = ~n63310;
  assign n63315 = ~n63282 | ~n63311;
  assign n63314 = ~n63313 | ~n63312;
  assign n63320 = ~n63316 & ~n74812;
  assign n63318 = ~n74806 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n63319 = ~n63318 | ~n68904;
  assign n63414 = ~n74276 | ~n63321;
  assign n63325 = ~n63406 ^ n63407;
  assign n63322 = ~n63325;
  assign n63326 = ~n63322 | ~n63323;
  assign n63324 = ~n63323;
  assign n63330 = n63329 | n63328;
  assign n63332 = ~n63247 | ~n63339;
  assign n63336 = ~n63332 | ~n63331;
  assign n63335 = ~n63334 | ~n63333;
  assign n63427 = ~n63336 | ~n63335;
  assign n63426 = ~n59905 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n63342 = ~n63340 ^ n63339;
  assign n63393 = ~n74835 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n63344 = ~n63393;
  assign n63389 = ~n76056 & ~n74846;
  assign n63352 = ~n63386;
  assign n63440 = ~n74315 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n63442 = ~n63296 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n63354 = ~n63440 ^ n63442;
  assign n63359 = ~n63439;
  assign n63369 = ~n63361 | ~n63360;
  assign n63364 = ~n63363 ^ n63362;
  assign n63367 = ~n63365 ^ n63364;
  assign n63370 = ~n63448;
  assign n63451 = ~n74798 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n63371 = ~n63370 ^ n63451;
  assign n63459 = ~n63450 ^ n63371;
  assign n63462 = ~n76000 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63376 = ~n63459 ^ n63462;
  assign n63461 = ~n63374 | ~n63373;
  assign n63375 = ~n63458 | ~n63461;
  assign n63679 = ~n63472 ^ n63470;
  assign n63469 = n59930 & P4_DATAO_REG_3__SCAN_IN;
  assign n63377 = ~n63469;
  assign n63571 = ~n63679 ^ n63377;
  assign n63385 = ~n63378 | ~n63571;
  assign n63565 = ~n63379;
  assign n63383 = ~n63565 | ~n63574;
  assign n63381 = ~n63574 | ~n63706;
  assign n63380 = ~n63572;
  assign n63384 = ~n63383 | ~n63382;
  assign n63388 = ~n63386;
  assign n63392 = ~n63388 | ~n63387;
  assign n63391 = ~n63390 | ~n63389;
  assign n63652 = ~n63392 | ~n63391;
  assign n63394 = ~n63642;
  assign n63397 = ~n63394 | ~n60750;
  assign n63396 = ~n63642 | ~n63402;
  assign n63401 = ~n63397 | ~n63396;
  assign n63399 = ~n63642 | ~n63855;
  assign n63398 = n63404 & n63005;
  assign n63400 = ~n63399 | ~n63398;
  assign n63403 = ~n63642 | ~n74846;
  assign n63405 = ~n63403 | ~n63402;
  assign n63641 = ~n63404;
  assign n63430 = ~n63405 | ~n63641;
  assign n63408 = ~n63406;
  assign n63616 = ~n63408 | ~n63407;
  assign n63410 = P4_DATAO_REG_15__SCAN_IN | n64259;
  assign n63867 = ~DIN_0_ | ~P4_DATAO_REG_15__SCAN_IN;
  assign n63409 = ~n68904 | ~n63867;
  assign n63411 = ~n63410 | ~n63409;
  assign n63413 = ~n74812 & ~n63411;
  assign n63600 = ~n59870 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n63416 = ~n63415 | ~n63414;
  assign n63615 = ~n63613;
  assign n63422 = ~n63614 ^ n63417;
  assign n63418 = ~n63625 & ~n59912;
  assign n63419 = ~n64572 | ~n59911;
  assign n63420 = ~n62954 | ~n59909;
  assign n63421 = ~n63624 | ~n63420;
  assign n63634 = ~n74835 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n63425 = ~n63634;
  assign n63428 = n63427 | n63426;
  assign n63597 = ~n63296 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n63435 = ~n63434 | ~n63433;
  assign n63908 = ~n63436 | ~n63435;
  assign n63443 = ~n63441 ^ n63440;
  assign n63658 = ~n63445 | ~n63444;
  assign n63446 = ~n74798 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n63455 = ~n63449 | ~n63448;
  assign n63453 = ~n63450;
  assign n63452 = ~n63451;
  assign n63667 = ~n76000 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n63456 = ~n63667;
  assign n63457 = n63461 & n63462;
  assign n63464 = ~n63461 | ~n76012;
  assign n63463 = ~n63462;
  assign n63467 = ~n63466 | ~n63465;
  assign n63590 = ~n59930 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63682 = ~n76054 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63471 = ~n63470;
  assign n63475 = ~n76037 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63476 = ~n63475;
  assign n63582 = n64350 & P4_DATAO_REG_1__SCAN_IN;
  assign n63693 = ~n63584 ^ n63582;
  assign n63480 = ~n63478;
  assign n63560 = ~n63480 ^ n63479;
  assign n63558 = ~n59930 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63700 = ~n63560 ^ n63558;
  assign n63485 = ~n63482 ^ n63481;
  assign n63484 = ~n63488 | ~n63483;
  assign n63544 = ~n63485 ^ n63484;
  assign n63541 = ~n63488 | ~n63487;
  assign n63540 = ~n63296 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63709 = ~n63541 ^ n63540;
  assign n63537 = ~n63106 ^ n63489;
  assign n63493 = ~n63490;
  assign n63492 = ~n63491;
  assign n63494 = n63493 | n63492;
  assign n63531 = ~n63495 | ~n63494;
  assign n63527 = ~n63497 ^ n63496;
  assign n63498 = n71397 & n74277;
  assign n63501 = ~n74812 & ~n63498;
  assign n63499 = ~n60375 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63500 = ~n63499 | ~n74763;
  assign n63503 = ~n63501 | ~n63500;
  assign n63510 = ~n63502;
  assign n63505 = n63503 | n63510;
  assign n63506 = ~n71188 & ~n63724;
  assign n63717 = ~n63505 ^ n63506;
  assign n72811 = ~n71188 & ~n74277;
  assign n63723 = ~n72811 | ~n60375;
  assign n63716 = ~n63723 & ~n71397;
  assign n63509 = ~n63717 | ~n63716;
  assign n63507 = ~n63505;
  assign n63508 = ~n63507 | ~n63506;
  assign n63512 = ~n63509 | ~n63508;
  assign n63513 = ~n63511 ^ n63510;
  assign n63732 = ~n63512 ^ n63513;
  assign n63731 = ~n59940 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63515 = n63732 | n63731;
  assign n63514 = ~n63513 | ~n63512;
  assign n63523 = ~n63515 | ~n63514;
  assign n63522 = ~n71188 & ~n59910;
  assign n63715 = ~n63523 ^ n63522;
  assign n63519 = ~n63516;
  assign n63518 = ~n63517;
  assign n63520 = n63519 | n63518;
  assign n63714 = ~n63521 | ~n63520;
  assign n63525 = n63715 | n63714;
  assign n63524 = ~n63523 | ~n63522;
  assign n63526 = ~n63525 | ~n63524;
  assign n63742 = ~n63527 ^ n63526;
  assign n63741 = ~n74835 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63529 = n63742 | n63741;
  assign n63528 = ~n63527 | ~n63526;
  assign n63532 = ~n63529 | ~n63528;
  assign n63713 = ~n63531 ^ n63532;
  assign n63712 = ~n63005 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63530 = ~n63712;
  assign n63535 = ~n63713 | ~n63530;
  assign n63533 = ~n63531;
  assign n63534 = ~n63533 | ~n63532;
  assign n63536 = ~n63535 | ~n63534;
  assign n63755 = ~n63537 ^ n63536;
  assign n63754 = ~n74315 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63539 = n63755 | n63754;
  assign n63538 = ~n63537 | ~n63536;
  assign n63710 = ~n63539 | ~n63538;
  assign n63543 = n63709 | n63710;
  assign n63542 = ~n63541 | ~n63540;
  assign n63545 = ~n63543 | ~n63542;
  assign n63708 = ~n63544 ^ n63545;
  assign n63707 = ~n74798 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63547 = n63708 | n63707;
  assign n63546 = n63545 | n63544;
  assign n63555 = ~n63547 | ~n63546;
  assign n63551 = ~n63548;
  assign n63550 = ~n63549;
  assign n63702 = ~n63555 ^ n63554;
  assign n63703 = ~n76000 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63557 = n63702 | n63703;
  assign n63556 = ~n63555 | ~n63554;
  assign n63559 = ~n63558;
  assign n63561 = ~n63560 | ~n63559;
  assign n63568 = ~n63562 | ~n63561;
  assign n63567 = ~n71188 & ~n74360;
  assign n63699 = ~n63568 ^ n63567;
  assign n63564 = ~n63563;
  assign n63566 = ~n63565 | ~n63564;
  assign n63698 = ~n63575 | ~n63566;
  assign n63569 = ~n63568 | ~n63567;
  assign n63579 = ~n63570 | ~n63569;
  assign n63573 = ~n63571;
  assign n63577 = ~n63573 ^ n63572;
  assign n63576 = ~n63575 | ~n63574;
  assign n63578 = ~n63577 ^ n63576;
  assign n63697 = ~n63579 ^ n63578;
  assign n63696 = ~n76037 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63580 = ~n63579 | ~n63578;
  assign n63694 = ~n63581 | ~n63580;
  assign n63583 = ~n63582;
  assign n63692 = ~n63589 | ~n63799;
  assign n63593 = ~n63592 | ~n63591;
  assign n63595 = ~n63596 | ~n63597;
  assign n63599 = ~n63595 | ~n63908;
  assign n63906 = ~n63597;
  assign n63598 = ~n63907 | ~n63906;
  assign n63602 = n63601 | n63600;
  assign n63605 = ~n63603 | ~n63317;
  assign n76062 = ~P4_DATAO_REG_15__SCAN_IN;
  assign n63604 = ~n76062 | ~n64033;
  assign n63606 = ~n63605 | ~n63604;
  assign n63608 = ~n74812 & ~n63606;
  assign n64036 = ~n74276 | ~n63607;
  assign n63871 = ~n63608 | ~n64036;
  assign n63873 = ~n60722 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n63609 = ~n63874 ^ n63873;
  assign n63883 = ~n63871 ^ n63609;
  assign n63610 = ~n63885;
  assign n63612 = ~n63611 | ~n63610;
  assign n63621 = ~n63614 | ~n63613;
  assign n63617 = n63616 & n63615;
  assign n63890 = ~n63621 | ~n63620;
  assign n63893 = ~n59906 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n63622 = ~n63890 ^ n63893;
  assign n63626 = n63625 | n59923;
  assign n63628 = ~n63627 | ~n63626;
  assign n63629 = ~n63628 | ~n59909;
  assign n63891 = ~n63630 | ~n63629;
  assign n63848 = ~n64011 | ~n63633;
  assign n63637 = ~n63636 | ~n63635;
  assign n63996 = ~n76045 & ~n59984;
  assign n63835 = ~n74416 & ~n74846;
  assign n63639 = ~n63835;
  assign n63640 = ~n63996 ^ n63639;
  assign n63643 = n63642 | n63641;
  assign n63645 = ~n63644 | ~n63643;
  assign n63646 = ~n63645 | ~n63005;
  assign n63648 = ~n63652;
  assign n63650 = ~n63648 | ~n63651;
  assign n63655 = ~n63650 | ~n63649;
  assign n63654 = ~n63653 | ~n63652;
  assign n63974 = ~n63296 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n63904 = ~n76064 & ~n76012;
  assign n63914 = ~n63904;
  assign n63916 = ~n76000 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n63661 = ~n63915 ^ n61551;
  assign n63660 = ~n63657;
  assign n63659 = ~n63658;
  assign n63664 = ~n63661;
  assign n63830 = n59930 & P4_DATAO_REG_5__SCAN_IN;
  assign n63665 = ~n63830;
  assign n63673 = ~n63666 ^ n63665;
  assign n63826 = ~n76054 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63674 = ~n63826;
  assign n63675 = n63681 & n63682;
  assign n63678 = ~n63676 | ~n63675;
  assign n63688 = ~n63678 | ~n63677;
  assign n63680 = ~n63679;
  assign n63686 = ~n63680 | ~n63681;
  assign n63684 = ~n63681 | ~n63706;
  assign n63683 = ~n63682;
  assign n63687 = ~n63686 | ~n63685;
  assign n63943 = ~n63688 | ~n63687;
  assign n63800 = n64350 & P4_DATAO_REG_2__SCAN_IN;
  assign n63689 = ~n63800;
  assign n63945 = ~n76037 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63690 = ~n63689 ^ n63945;
  assign n63932 = ~n63929 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63790 = ~n74930 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n63695 = ~n63693;
  assign n63787 = ~n63695 ^ n63694;
  assign n63785 = ~n63929 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n97644 = ~n63787 ^ n63785;
  assign n63782 = ~n63697 ^ n63696;
  assign n63781 = ~n64350 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n75021 = ~n63782 ^ n63781;
  assign n63778 = ~n63699 ^ n63698;
  assign n63777 = ~n76037 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n74469 = ~n63778 ^ n63777;
  assign n63701 = ~n63700;
  assign n63773 = ~n76054 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n71699 = ~n63772 ^ n63773;
  assign n63705 = ~n63702;
  assign n63704 = ~n63703;
  assign n63769 = ~n63705 ^ n63704;
  assign n63768 = ~n59930 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n71420 = ~n63769 ^ n63768;
  assign n63765 = ~n63708 ^ n63707;
  assign n63764 = ~n76000 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n70199 = ~n63765 ^ n63764;
  assign n63711 = ~n63709;
  assign n63761 = ~n63711 ^ n63710;
  assign n63760 = ~n74798 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n69006 = ~n63761 ^ n63760;
  assign n63749 = ~n63713 ^ n63712;
  assign n63750 = ~n74315 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n67465 = ~n63749 ^ n63750;
  assign n63748 = ~n67465;
  assign n63738 = ~n63715 ^ n63714;
  assign n63737 = ~n74835 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n78651 = ~n63738 ^ n63737;
  assign n63718 = ~n63717 ^ n63716;
  assign n63719 = ~n62954 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n63730 = n63718 | n63719;
  assign n76798 = n63719 ^ n63718;
  assign n63720 = ~n63723 ^ n63724;
  assign n73159 = ~n63720 & ~n71171;
  assign n63722 = ~n59914 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n63721 = ~n71397 & ~n74277;
  assign n73158 = ~n63722 ^ n63721;
  assign n63728 = ~n73159 | ~n73158;
  assign n63726 = ~n63723;
  assign n63725 = ~n71171 & ~n63724;
  assign n63727 = ~n63726 | ~n63725;
  assign n76797 = ~n63728 | ~n63727;
  assign n63729 = ~n76798 | ~n76797;
  assign n63734 = ~n63730 | ~n63729;
  assign n63733 = ~n71171 & ~n59911;
  assign n74125 = ~n63734 ^ n63733;
  assign n74124 = ~n63732 ^ n63731;
  assign n63736 = n74125 | n74124;
  assign n63735 = ~n63734 | ~n63733;
  assign n78650 = n63736 & n63735;
  assign n63740 = n78651 | n78650;
  assign n63739 = n63738 | n63737;
  assign n63744 = ~n63740 | ~n63739;
  assign n63743 = ~n71171 & ~n74846;
  assign n65162 = ~n63744 ^ n63743;
  assign n65161 = ~n63742 ^ n63741;
  assign n63746 = n65162 | n65161;
  assign n63745 = ~n63744 | ~n63743;
  assign n67466 = ~n63746 | ~n63745;
  assign n63747 = ~n67466;
  assign n63753 = n63748 | n63747;
  assign n63751 = ~n63749;
  assign n63752 = n63751 | n63750;
  assign n63757 = ~n63753 | ~n63752;
  assign n63756 = ~n71171 & ~n60217;
  assign n67984 = ~n63757 ^ n63756;
  assign n67985 = ~n63755 ^ n63754;
  assign n63759 = n67984 | n67985;
  assign n63758 = ~n63757 | ~n63756;
  assign n69007 = n63759 & n63758;
  assign n63763 = n69006 | n69007;
  assign n63762 = n63761 | n63760;
  assign n70200 = n63763 & n63762;
  assign n63767 = n70199 | n70200;
  assign n63766 = n63765 | n63764;
  assign n63771 = n71420 | n71419;
  assign n63770 = n63769 | n63768;
  assign n71700 = ~n63771 | ~n63770;
  assign n63776 = ~n71699 | ~n71700;
  assign n63774 = ~n63772;
  assign n63780 = n74469 | n74470;
  assign n63779 = n63778 | n63777;
  assign n63784 = n75021 | n75022;
  assign n63783 = n63782 | n63781;
  assign n97643 = ~n63784 | ~n63783;
  assign n63789 = ~n97644 | ~n97643;
  assign n63786 = ~n63785;
  assign n63788 = ~n63787 | ~n63786;
  assign n63938 = n76051 & P4_DATAO_REG_0__SCAN_IN;
  assign n63960 = ~n59980 | ~n74367;
  assign n63793 = ~n63960 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n63794 = ~n63799 | ~n63793;
  assign n63795 = ~n63794 | ~n63945;
  assign n63805 = ~n63797 | ~n63808;
  assign n63801 = ~n63799 | ~n74367;
  assign n63804 = ~n63803 | ~n63802;
  assign n63806 = ~n63945 & ~n71397;
  assign n63942 = ~n63810;
  assign n63811 = n63943 | n76037;
  assign n63944 = ~n64350 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n63948 = ~n63944;
  assign n63812 = ~n63811 | ~n63948;
  assign n63825 = ~n63942 & ~n63812;
  assign n63814 = n63943 | n64350;
  assign n63813 = ~n63960;
  assign n63816 = ~n63813 & ~n74763;
  assign n63815 = ~n63814 | ~n63816;
  assign n63823 = ~n63815 | ~n63942;
  assign n63817 = ~n63816;
  assign n63821 = n63943 | n63817;
  assign n63818 = ~n63945;
  assign n63819 = ~n63818 | ~n64350;
  assign n63820 = ~n63943 | ~n63819;
  assign n63822 = ~n63821 | ~n63820;
  assign n63824 = ~n63823 | ~n63822;
  assign n64142 = ~n63829 | ~n63828;
  assign n63998 = ~n63836 | ~n63852;
  assign n63840 = ~n63998 & ~n63837;
  assign n63839 = ~n63999 & ~n63841;
  assign n63842 = ~n63841;
  assign n63844 = ~n63999 | ~n63843;
  assign n63846 = ~n63845 | ~n63844;
  assign n63982 = ~n74798 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n63850 = ~n63848;
  assign n63851 = ~n63850 | ~n63849;
  assign n64007 = ~n63852 | ~n63851;
  assign n63853 = ~n59846 | ~n59912;
  assign n63854 = ~n64052;
  assign n63856 = ~n59910 | ~n63855;
  assign n63857 = n63890 | n63860;
  assign n63859 = ~n59912 & ~n63855;
  assign n63861 = ~n63890 | ~n63859;
  assign n63865 = ~n63864 | ~n64052;
  assign n64041 = ~n76062 & ~n60721;
  assign n63866 = ~n64041;
  assign n63869 = ~n64038 ^ n63866;
  assign n63868 = ~n63867 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n64037 = ~n63868 & ~n63317;
  assign n64267 = ~n63869 ^ n64037;
  assign n64016 = ~n59905 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n63870 = ~n64266 ^ n64016;
  assign n63872 = ~n63871;
  assign n63876 = ~n63872 | ~n61571;
  assign n63875 = n63874 | n63873;
  assign n63880 = ~n63888;
  assign n63879 = ~n59857 | ~n63878;
  assign n63881 = n63880 & n63879;
  assign n63889 = ~n63882 | ~n63881;
  assign n63884 = ~n59857 | ~n63885;
  assign n63887 = ~n63884 | ~n63883;
  assign n64066 = ~n63005 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n63894 = ~n64052 ^ n59846;
  assign n63892 = ~n63894 | ~n63893;
  assign n63895 = n63891 & n63892;
  assign n64220 = ~n64007 ^ n64008;
  assign n64006 = ~n74315 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n63900 = ~n63976 | ~n61158;
  assign n63901 = ~n63900 | ~n63981;
  assign n64090 = ~n63905 | ~n63904;
  assign n63909 = ~n63908 | ~n63907;
  assign n63911 = ~n63910 | ~n63909;
  assign n64092 = ~n63912 | ~n63911;
  assign n64091 = ~n76000 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n64094 = ~n64091;
  assign n63913 = ~n64095 ^ n64094;
  assign n64099 = ~n63913 ^ n64093;
  assign n63920 = ~n64099;
  assign n63919 = ~n63917 | ~n63916;
  assign n63922 = ~n63924;
  assign n63921 = ~n63923;
  assign n63925 = ~n63922 | ~n63921;
  assign n64168 = ~n76081 & ~n74360;
  assign n64104 = ~n64168;
  assign n63957 = ~n76037 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63926 = ~n60834 ^ n63957;
  assign n63947 = ~n63926 ^ n64157;
  assign n63927 = ~n63947;
  assign n64108 = n63929 & P4_DATAO_REG_2__SCAN_IN;
  assign n63930 = ~n64108;
  assign n64120 = ~n71188 & ~n76061;
  assign n64119 = ~n64122 ^ n64120;
  assign n63937 = n63933 | n63932;
  assign n63936 = ~n63935 | ~n63934;
  assign n64118 = ~n63937 | ~n63936;
  assign n72805 = ~n64119 ^ n64118;
  assign n63940 = ~n63939 | ~n63938;
  assign n64124 = n76067 & P4_DATAO_REG_0__SCAN_IN;
  assign n63949 = ~n63950 | ~n74367;
  assign n63953 = ~n63952 | ~n63951;
  assign n64154 = ~n64350 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63954 = ~n64154;
  assign n63955 = ~n60834 | ~n74367;
  assign n63964 = ~n63956 | ~n63955;
  assign n63958 = ~n63957;
  assign n63959 = ~n63958 | ~n64350;
  assign n63962 = ~n64156 | ~n63959;
  assign n64146 = ~n63960 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n63965 = ~n64146;
  assign n63961 = ~n60834 | ~n63965;
  assign n63963 = ~n63962 | ~n63961;
  assign n63967 = ~n64157;
  assign n64137 = ~n64147 | ~n59980;
  assign n63966 = ~n64137 | ~n63965;
  assign n63969 = ~n60761 | ~n63976;
  assign n63971 = ~n63976;
  assign n63973 = ~n63972 & ~n63971;
  assign n63975 = ~n63974 & ~n76012;
  assign n63977 = ~n63976 | ~n63975;
  assign n63979 = ~n64211;
  assign n64201 = ~n64196;
  assign n63986 = ~n64201 ^ n74881;
  assign n63994 = ~n63979 | ~n63986;
  assign n63985 = ~n60763 | ~n61159;
  assign n63983 = ~n63981;
  assign n63984 = ~n63983 | ~n61160;
  assign n63988 = ~n64209 | ~n63986;
  assign n63987 = ~n64196 | ~n76056;
  assign n63991 = ~n64196 | ~n74881;
  assign n63989 = ~n76056 & ~n74881;
  assign n63990 = ~n64201 | ~n63989;
  assign n63992 = n63991 & n63990;
  assign n63995 = ~n63998;
  assign n64002 = ~n63995 | ~n63996;
  assign n63997 = ~n63996;
  assign n64000 = ~n63998 | ~n63997;
  assign n64001 = ~n64000 | ~n63999;
  assign n64003 = ~n64002 | ~n64001;
  assign n64004 = ~n64003 | ~n63296;
  assign n64087 = ~n64005 | ~n64004;
  assign n64309 = ~n64218 | ~n64221;
  assign n64073 = ~n64066;
  assign n64009 = ~n64075 | ~n64073;
  assign n64014 = ~n64009 | ~n64068;
  assign n64012 = n64010 & n64066;
  assign n64013 = ~n64012 | ~n64011;
  assign n64236 = ~n64014 | ~n64013;
  assign n64062 = ~n64236 ^ n64015;
  assign n64017 = ~n64016;
  assign n64271 = ~n59906 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n64027 = ~n64271;
  assign n64029 = ~n64267;
  assign n64020 = ~n64027 | ~n64266;
  assign n64021 = ~n60926 | ~n64271;
  assign n64023 = ~n64022 | ~n64021;
  assign n64025 = ~n64024 | ~n64023;
  assign n64030 = ~n64028 | ~n64027;
  assign n64262 = ~n64032 & ~n71293;
  assign n64034 = ~n64251 | ~n64033;
  assign n64035 = ~n64038 | ~n59870;
  assign n64045 = ~n62954 | ~P4_DATAO_REG_15__SCAN_IN;
  assign n64040 = ~n64037;
  assign n64039 = ~n64038;
  assign n64042 = ~n64040 | ~n64039;
  assign n64043 = ~n64042 | ~n64041;
  assign n64241 = ~n64044 | ~n64043;
  assign n64046 = ~n64242 ^ n64241;
  assign n64047 = ~n64046 | ~n64045;
  assign n64048 = ~n74835 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n64050 = ~n64049 | ~n64048;
  assign n64286 = ~n64240 | ~n64050;
  assign n64284 = ~n64051 & ~n74846;
  assign n64060 = ~n64283;
  assign n64053 = n64052 | n59846;
  assign n64055 = ~n64054 | ~n64053;
  assign n64058 = ~n64055 | ~n74835;
  assign n64083 = ~n64062 | ~n64061;
  assign n64072 = ~n64063 | ~n64075;
  assign n64064 = ~n64065 | ~n64073;
  assign n64070 = ~n64074 | ~n64064;
  assign n64067 = ~n64015 | ~n64066;
  assign n64069 = ~n64068 | ~n64067;
  assign n64071 = ~n64070 | ~n64069;
  assign n64080 = ~n64072 | ~n64071;
  assign n64078 = n64074 & n64073;
  assign n64076 = ~n64075;
  assign n64077 = ~n64015 | ~n64076;
  assign n64079 = ~n64078 & ~n64077;
  assign n64082 = ~n64080 & ~n64079;
  assign n64222 = ~n63296 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n64310 = ~n74798 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n64084 = ~n64222 ^ n64310;
  assign n64085 = ~n64307 ^ n64084;
  assign n64086 = ~n64085 ^ n64309;
  assign n64313 = ~n64087 | ~n64086;
  assign n64199 = ~n64208;
  assign n64097 = ~n64089 ^ n64199;
  assign n64096 = ~n64095 | ~n64094;
  assign n64185 = ~n64097 ^ n64200;
  assign n64098 = ~n64185;
  assign n64187 = ~n76054 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n64102 = ~n64098 ^ n64187;
  assign n64186 = n64100 | n64099;
  assign n64101 = ~n64180 | ~n64186;
  assign n64171 = ~n64102 ^ n64101;
  assign n64103 = ~n64166 | ~n64104;
  assign n64106 = ~n64103 | ~n64165;
  assign n64107 = ~n64106 | ~n64105;
  assign n64139 = ~n64171 ^ n64107;
  assign n64150 = ~n64139;
  assign n64164 = ~n76037 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n64131 = ~n63929 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n64114 = ~n64109 | ~n64108;
  assign n64111 = ~n64110;
  assign n64113 = ~n64112 | ~n64111;
  assign n64319 = n76051 & P4_DATAO_REG_1__SCAN_IN;
  assign n64123 = ~n64117 ^ n64319;
  assign n64323 = ~n64119 | ~n64118;
  assign n64121 = ~n64120;
  assign n73154 = ~n64123 ^ n64318;
  assign n64126 = ~n64125 | ~n64124;
  assign n64129 = ~n64128 | ~n64127;
  assign n64135 = ~n64134 | ~n64133;
  assign n64141 = ~n64137 & ~n64157;
  assign n64138 = ~n64173 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n64140 = n64139 & n64138;
  assign n64153 = ~n64141 & ~n64140;
  assign n64143 = n64142 & n64146;
  assign n64145 = ~n64144 | ~n64143;
  assign n64149 = n64145 & n64164;
  assign n64148 = ~n60834 | ~n64146;
  assign n64151 = ~n64149 | ~n64148;
  assign n64152 = ~n64151 | ~n64150;
  assign n64162 = ~n64153 | ~n64152;
  assign n64155 = ~n64157 & ~n64156;
  assign n64160 = ~n64155 & ~n64154;
  assign n64158 = ~n64157 | ~n64156;
  assign n64159 = ~n64158 | ~n74367;
  assign n64161 = ~n64160 | ~n64159;
  assign n64175 = ~n64163 | ~n64165;
  assign n64170 = n64175 & n64164;
  assign n64167 = ~n64165;
  assign n64174 = ~n64167 | ~n64166;
  assign n64169 = ~n64174 | ~n64168;
  assign n64172 = ~n64170 | ~n64169;
  assign n64179 = ~n64172 | ~n64171;
  assign n64176 = ~n64175 | ~n74360;
  assign n64178 = ~n64177 | ~n64176;
  assign n64525 = ~n64350 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n64181 = ~n64187;
  assign n64184 = ~n64186 | ~n64187;
  assign n64188 = ~n64186;
  assign n64189 = ~n64188 | ~n64181;
  assign n64192 = ~n64200 | ~n64208;
  assign n64191 = ~n64208 | ~n64196;
  assign n64195 = ~n64192 | ~n64191;
  assign n64193 = ~n64209;
  assign n64194 = ~n64214 ^ n74881;
  assign n64197 = ~n64200 | ~n64196;
  assign n64207 = ~n64198 | ~n64197;
  assign n64203 = ~n64200 | ~n64199;
  assign n64202 = n64208 | n64201;
  assign n64205 = ~n64203 | ~n64202;
  assign n64213 = ~n64208 & ~n76056;
  assign n64210 = ~n64209 & ~n76000;
  assign n64212 = ~n64211 | ~n64210;
  assign n64216 = ~n64213 | ~n64212;
  assign n64215 = ~n64214 | ~n76000;
  assign n64353 = ~n64216 | ~n64215;
  assign n64217 = n64221 & n64222;
  assign n64435 = ~n74798 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n64230 = ~n64443 ^ n64447;
  assign n64219 = ~n64307 & ~n64230;
  assign n64229 = ~n60718 | ~n64219;
  assign n64223 = ~n64221 | ~n59984;
  assign n64306 = ~n64222;
  assign n64436 = ~n64225 | ~n64224;
  assign n64227 = ~n64436;
  assign n64226 = ~n64230;
  assign n64228 = ~n64227 | ~n64226;
  assign n64233 = n64436 & n64230;
  assign n64234 = ~n64233 | ~n64437;
  assign n64305 = ~n64235 | ~n64234;
  assign n64419 = ~n64240 | ~n64239;
  assign n64243 = ~n64242 | ~n64241;
  assign n64403 = ~n64244 | ~n64243;
  assign n64567 = ~n74361 & ~n64572;
  assign n64246 = ~n64567 | ~n59870;
  assign n64392 = ~n60722 | ~P4_DATAO_REG_17__SCAN_IN;
  assign n64245 = ~n64390 | ~n64392;
  assign n64248 = ~n64262;
  assign n64253 = ~n64262 | ~n60483;
  assign n64254 = ~n64387;
  assign n64256 = ~n64390;
  assign n64257 = ~n64256 ^ n64392;
  assign n64258 = ~n64257 | ~n64387;
  assign n64583 = ~n64262 | ~n64260;
  assign n64381 = ~n64262 | ~n64261;
  assign n64264 = ~n64583 ^ n64381;
  assign n64265 = n64267 | n64266;
  assign n64268 = ~n64267 | ~n64266;
  assign n64272 = ~n64270 | ~n64273;
  assign n64276 = ~n64272 | ~n64271;
  assign n64274 = ~n64273;
  assign n64277 = ~n64407;
  assign n64410 = ~n74835 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n64278 = ~n64277 ^ n64410;
  assign n64418 = ~n64406 ^ n64278;
  assign n64280 = ~n64419 ^ n64418;
  assign n64279 = ~n74396 & ~n74846;
  assign n64422 = ~n64280 | ~n64279;
  assign n64285 = ~n64284;
  assign n64287 = ~n64286 | ~n64285;
  assign n64427 = ~n74315 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n64291 = ~n64289;
  assign n64302 = ~n71230 & ~n60217;
  assign n64290 = ~n64302;
  assign n64293 = ~n64425 | ~n64292;
  assign n64300 = ~n64293 | ~n64297;
  assign n64294 = ~n64427;
  assign n64298 = ~n64296 | ~n64295;
  assign n64299 = ~n64298 | ~n64426;
  assign n64308 = ~n64307 ^ n64306;
  assign n64311 = ~n64309 ^ n64308;
  assign n64355 = ~n59930 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n64349 = ~n76054 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n64315 = ~n64314 | ~n61146;
  assign n64339 = ~n64335;
  assign n64334 = n76051 & P4_DATAO_REG_2__SCAN_IN;
  assign n64338 = ~n64334;
  assign n64317 = ~n64339 ^ n64338;
  assign n64492 = ~n64337 ^ n64317;
  assign n64327 = ~n64318 | ~n64319;
  assign n64320 = ~n64319;
  assign n64322 = n64321 & n64320;
  assign n64324 = ~n64323 | ~n64322;
  assign n64326 = ~n64325 | ~n64324;
  assign n64490 = ~n64492 ^ n64491;
  assign n64489 = ~n76067 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n64330 = ~n76043 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n64331 = ~n64329;
  assign n64495 = n76076 & P4_DATAO_REG_0__SCAN_IN;
  assign n64340 = ~n64339 | ~n64338;
  assign n64341 = ~n64342 | ~n61535;
  assign n64470 = ~n64523;
  assign n64526 = ~n63929 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n64346 = ~n64464 | ~n64526;
  assign n64777 = ~n64350 & ~n63929;
  assign n64344 = ~n64777 & ~n76081;
  assign n64345 = ~n64463 | ~n64344;
  assign n64461 = ~n64346 | ~n64345;
  assign n64539 = ~n64350 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n64351 = ~n64536;
  assign n64356 = ~n64354 | ~n64353;
  assign n64358 = ~n64357;
  assign n64622 = n64359 | n64358;
  assign n64617 = ~n71230 & ~n76012;
  assign n64551 = ~n76000 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n64360 = ~n64617 ^ n64551;
  assign n64434 = ~n64618 ^ n64360;
  assign n64363 = n64362 & n64361;
  assign n64584 = ~n64366 | ~n64365;
  assign n64368 = ~n64584;
  assign n64372 = ~n64368 | ~n59870;
  assign n64370 = ~n64369;
  assign n64371 = ~n64370 | ~n64706;
  assign n64374 = ~n64372 | ~n64371;
  assign n64373 = ~n64583;
  assign n64379 = ~n64374 | ~n64373;
  assign n64377 = ~n64584 ^ n64376;
  assign n64378 = ~n64377 | ~n64583;
  assign n64382 = ~n64381;
  assign n64383 = ~n64382 | ~n64583;
  assign n64385 = ~n64387 | ~n64390;
  assign n64388 = n64387 | n64390;
  assign n64393 = ~n64391 | ~n64390;
  assign n64394 = n64393 & n64380;
  assign n64398 = ~n59907 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n64600 = ~n64596 | ~n64399;
  assign n64404 = ~n64403 | ~n64402;
  assign n64601 = ~n74835 | ~P4_DATAO_REG_15__SCAN_IN;
  assign n64413 = ~n64408;
  assign n64411 = ~n64410;
  assign n64416 = ~n63005 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n64561 = ~n64608 | ~n64417;
  assign n64420 = ~n64418;
  assign n64421 = ~n64420 | ~n64419;
  assign n64423 = ~n64422 | ~n64421;
  assign n64429 = ~n64426 | ~n64425;
  assign n64555 = ~n63296 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n64430 = ~n64555;
  assign n64620 = ~n64557 ^ n64432;
  assign n64433 = ~n64620;
  assign n64438 = ~n64445 | ~n64435;
  assign n64439 = ~n64438 | ~n64444;
  assign n64441 = ~n64440 | ~n64439;
  assign n64448 = ~n64447;
  assign n64453 = ~n64449 | ~n64448;
  assign n64454 = ~n64632 ^ n60802;
  assign n64458 = ~n64457 | ~n64456;
  assign n64469 = ~n64461 | ~n64527;
  assign n64462 = ~n64528 | ~n59980;
  assign n64466 = ~n64463 | ~n64462;
  assign n64464 = ~n64463;
  assign n64465 = ~n64464 | ~n64528;
  assign n64467 = ~n64466 | ~n64465;
  assign n64468 = ~n64467 | ~n64475;
  assign n64471 = ~n64477;
  assign n64474 = ~n64473 | ~n64472;
  assign n64476 = ~n64475 | ~n64528;
  assign n64479 = ~n64478 | ~n64477;
  assign n64509 = ~n74930 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n64515 = ~n64509;
  assign n64480 = ~n64511 | ~n64514;
  assign n64644 = n76051 & P4_DATAO_REG_3__SCAN_IN;
  assign n64482 = ~n64644;
  assign n64483 = ~n60503 ^ n64482;
  assign n64486 = ~n64487;
  assign n64499 = n76067 & P4_DATAO_REG_2__SCAN_IN;
  assign n64485 = ~n64499;
  assign n64488 = ~n64487 | ~n64499;
  assign n64655 = ~n64663 | ~n64488;
  assign n64653 = ~n76043 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n64494 = n64490 | n64489;
  assign n64493 = ~n64492 | ~n64491;
  assign n74120 = ~n64652 ^ n64651;
  assign n64498 = ~n64662;
  assign n64505 = n76043 & P4_DATAO_REG_2__SCAN_IN;
  assign n67369 = ~n64505;
  assign n64502 = ~n64498 | ~n67369;
  assign n64500 = n67369 & n64485;
  assign n64501 = ~n64504 | ~n64500;
  assign n64503 = ~n76067;
  assign n64507 = ~n64504 | ~n64503;
  assign n64510 = n64514 & n64509;
  assign n64518 = ~n64513 | ~n64514;
  assign n64516 = ~n64514 | ~n71345;
  assign n64519 = ~n64518 | ~n64517;
  assign n67214 = n76051 & P4_DATAO_REG_4__SCAN_IN;
  assign n64520 = ~n64530 | ~n59980;
  assign n64521 = ~n64520 | ~n64528;
  assign n64524 = ~n64522 | ~n64521;
  assign n64534 = ~n64524 | ~n64523;
  assign n64529 = ~n64528 | ~n64350;
  assign n64667 = ~n74930 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n64535 = ~n64667;
  assign n64538 = ~n64636 | ~n64775;
  assign n64541 = ~n64635 ^ n64538;
  assign n64540 = ~n64539;
  assign n64542 = ~n64541 | ~n64540;
  assign n64547 = ~n64543 | ~n64542;
  assign n64545 = ~n64547;
  assign n64544 = ~n64546;
  assign n64673 = ~n64547 | ~n64546;
  assign n64769 = ~n76056 & ~n74367;
  assign n64621 = ~n64617;
  assign n64550 = ~n64618 ^ n64621;
  assign n64553 = ~n64550 ^ n64620;
  assign n64552 = ~n64551;
  assign n64554 = ~n64553 | ~n64552;
  assign n64559 = ~n64556 | ~n64555;
  assign n64739 = ~n76000 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n64560 = ~n59961 ^ n64739;
  assign n64563 = ~n64561;
  assign n64564 = ~n64563 | ~n64562;
  assign n64569 = ~n64568 | ~n64567;
  assign n64570 = P4_DATAO_REG_19__SCAN_IN & P4_DATAO_REG_20__SCAN_IN;
  assign n64571 = ~n71279 & ~n61061;
  assign n67274 = ~n64571 | ~n60715;
  assign n64575 = ~n64574 | ~n71279;
  assign n64582 = n64584 | n64583;
  assign n64585 = ~n64584 | ~n64583;
  assign n64698 = ~n64586 | ~n64585;
  assign n67291 = ~n64588 ^ n64587;
  assign n67293 = ~n74361 & ~n59911;
  assign n64725 = ~n74835 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n64591 = ~n64590 | ~n64589;
  assign n64594 = n64592 & n64591;
  assign n64595 = ~n64594 | ~n64593;
  assign n64598 = ~n64596 | ~n64595;
  assign n64597 = ~n64598;
  assign n64729 = ~n64598 | ~n64599;
  assign n64602 = ~n60773 | ~n64601;
  assign n64730 = ~n64603 | ~n64602;
  assign n64605 = ~n64731 ^ n64730;
  assign n64604 = ~n63005 | ~P4_DATAO_REG_15__SCAN_IN;
  assign n64733 = n64605 | n64604;
  assign n64606 = ~n64605 | ~n64604;
  assign n64684 = ~n64733 | ~n64606;
  assign n64685 = ~n64608 | ~n64607;
  assign n64609 = ~n68904 & ~n59984;
  assign n64610 = ~n63296 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n64611 = P4_DATAO_REG_14__SCAN_IN & DIN_7_;
  assign n64615 = DIN_8_ & P4_DATAO_REG_13__SCAN_IN;
  assign n64738 = ~n64679 | ~n64683;
  assign n64619 = ~n64618 | ~n64617;
  assign n64625 = ~n64620 | ~n64619;
  assign n64623 = n64622 & n64621;
  assign n64634 = ~n64631 | ~n64630;
  assign n64757 = ~n76054 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n67229 = n64350 & P4_DATAO_REG_7__SCAN_IN;
  assign n64637 = ~n67229;
  assign n64638 = ~n64774 ^ n64637;
  assign n64674 = ~n67228 ^ n64638;
  assign n64639 = ~n64674;
  assign n64670 = ~n64640 ^ n64639;
  assign n64641 = n76067 & P4_DATAO_REG_3__SCAN_IN;
  assign n64648 = ~n64645 | ~n64644;
  assign n64649 = ~n64666;
  assign n64654 = ~n64653;
  assign n64656 = ~n64655 | ~n64654;
  assign n64658 = ~n76046 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n67387 = ~n64657;
  assign n64660 = ~n64659;
  assign n67195 = ~n64660 | ~n60814;
  assign n64665 = ~n67377;
  assign n64664 = ~n67371 | ~n76043;
  assign n64803 = ~n64665 | ~n64664;
  assign n64668 = ~n64669 | ~n64670;
  assign n64672 = ~n64668 | ~n64667;
  assign n67741 = ~n76051 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n64794 = ~n67743 ^ n67741;
  assign n64675 = ~n64674 | ~n64673;
  assign n64676 = ~n64683;
  assign n64680 = n64683 & n59961;
  assign n64681 = ~n64680 | ~n64679;
  assign n64736 = ~n67328 ^ n67330;
  assign n67323 = ~n74798 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n64686 = ~n64684;
  assign n64687 = ~n64686 | ~n64685;
  assign n67318 = ~n63296 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n64692 = ~n67296 | ~n67293;
  assign n64689 = ~n67293;
  assign n64690 = ~n67292 | ~n64689;
  assign n64691 = ~n64690 | ~n67295;
  assign n67251 = ~n63005 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n64723 = ~n67250 ^ n67251;
  assign n64696 = ~n64695 | ~n64694;
  assign n64700 = ~n64699 | ~n64698;
  assign n64703 = ~n63504 | ~P4_DATAO_REG_22__SCAN_IN;
  assign n64702 = ~n59913 | ~P4_DATAO_REG_21__SCAN_IN;
  assign n64705 = ~n64703 | ~n64702;
  assign n64704 = P4_DATAO_REG_21__SCAN_IN & P4_DATAO_REG_22__SCAN_IN;
  assign n64707 = ~n67274 | ~n64709;
  assign n64708 = ~n63724 | ~P4_DATAO_REG_22__SCAN_IN;
  assign n64711 = ~n64717 | ~n64708;
  assign n67276 = ~n67273 | ~n67272;
  assign n67279 = ~n74353 & ~n64572;
  assign n64714 = ~n67279;
  assign n64713 = ~n67287;
  assign n64716 = ~n64714 ^ n64713;
  assign n67262 = ~n71293 & ~n59911;
  assign n64715 = ~n67262;
  assign n64719 = n64718 | n64717;
  assign n67257 = ~n64720 | ~n64719;
  assign n64722 = ~n64721 ^ n67257;
  assign n67299 = ~n67261 ^ n64722;
  assign n67248 = ~n67299 ^ n64723;
  assign n64724 = ~n67295 ^ n67293;
  assign n64727 = ~n67296 ^ n64724;
  assign n64726 = ~n64725;
  assign n64728 = ~n64727 | ~n64726;
  assign n67247 = n64729 & n64728;
  assign n67313 = ~n74315 | ~P4_DATAO_REG_15__SCAN_IN;
  assign n64734 = ~n67310 ^ n67313;
  assign n64732 = n64731 | n64730;
  assign n64741 = ~n64738 ^ n64737;
  assign n64740 = ~n64739;
  assign n67335 = ~n64741 | ~n64740;
  assign n67334 = ~n59930 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n67338 = ~n67334;
  assign n67341 = ~n64743 | ~n64753;
  assign n64746 = ~n64744;
  assign n64747 = ~n64746 | ~n64745;
  assign n67342 = ~n64748 | ~n64747;
  assign n64749 = ~n67342;
  assign n64751 = ~n67341 ^ n64749;
  assign n64750 = ~n64755;
  assign n67243 = ~n64751 | ~n64750;
  assign n67239 = ~n76037 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n67242 = ~n67239;
  assign n67348 = ~n67354;
  assign n64763 = ~n64758 | ~n64757;
  assign n64760 = ~n64759;
  assign n64762 = ~n64761 | ~n64760;
  assign n67351 = ~n64763 | ~n64762;
  assign n64764 = ~n67350;
  assign n67346 = n67351 | n64764;
  assign n64765 = ~n67351 | ~n64764;
  assign n64773 = ~n64767 | ~n64766;
  assign n64771 = ~n64770 | ~n64769;
  assign n67226 = ~n63929 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n64778 = ~n67227;
  assign n64784 = ~n64777 & ~n76064;
  assign n64781 = ~n64778 | ~n64784;
  assign n64779 = ~n59972 | ~n64350;
  assign n64780 = ~n67227 | ~n64779;
  assign n64782 = ~n64781 | ~n64780;
  assign n64788 = ~n67228;
  assign n64786 = ~n67227 & ~n63929;
  assign n64789 = ~n64788 | ~n64787;
  assign n67221 = ~n71660 & ~n76061;
  assign n64793 = ~n67744;
  assign n64798 = ~n64797 | ~n64796;
  assign n67208 = ~n76067 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n64799 = ~n64798 ^ n67208;
  assign n67203 = n76043 & P4_DATAO_REG_3__SCAN_IN;
  assign n67374 = ~n76076 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n64802 = ~n67375 ^ n67374;
  assign n67198 = ~n64803 ^ n64802;
  assign n64804 = ~n67198;
  assign n67192 = n76046 & P4_DATAO_REG_1__SCAN_IN;
  assign n67194 = ~n67192;
  assign n64805 = ~n64804 ^ n67194;
  assign n67384 = ~n67193 ^ n64805;
  assign n76044 = ~n76028 | ~DIN_22_;
  assign n67390 = ~n71171 & ~n76044;
  assign n67381 = ~n67390;
  assign n100184 = ~P1_P1_STATE2_REG_2__SCAN_IN;
  assign n100434 = ~P1_P1_STATE2_REG_1__SCAN_IN;
  assign n96193 = ~n100434 | ~P1_P1_STATE2_REG_0__SCAN_IN;
  assign n97203 = ~n60799;
  assign n64810 = ~n97203 | ~P1_P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n97743 = ~n64808;
  assign n64809 = ~n97743 | ~P1_P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n64814 = ~n64810 | ~n64809;
  assign n64812 = ~n97761 | ~P1_P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n97998 = ~n100090 & ~n99991;
  assign n64811 = ~n97895 | ~P1_P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n64813 = ~n64812 | ~n64811;
  assign n64823 = ~n64814 & ~n64813;
  assign n64816 = ~P1_P1_INSTQUEUE_REG_4__7__SCAN_IN | ~n59935;
  assign n97754 = ~n61500;
  assign n64815 = ~P1_P1_INSTQUEUE_REG_9__7__SCAN_IN | ~n97754;
  assign n64821 = ~n64816 | ~n64815;
  assign n100108 = ~n65089 & ~n64824;
  assign n100123 = ~n100108;
  assign n64819 = ~P1_P1_INSTQUEUE_REG_6__7__SCAN_IN | ~n97747;
  assign n64818 = ~P1_P1_INSTQUEUE_REG_14__7__SCAN_IN | ~n97746;
  assign n64820 = ~n64819 | ~n64818;
  assign n64822 = ~n64821 & ~n64820;
  assign n64845 = ~n64823 | ~n64822;
  assign n64826 = ~P1_P1_INSTQUEUE_REG_5__7__SCAN_IN | ~n97979;
  assign n64825 = ~P1_P1_INSTQUEUE_REG_7__7__SCAN_IN | ~n97185;
  assign n64831 = ~n64826 | ~n64825;
  assign n97303 = ~n61526;
  assign n64829 = ~P1_P1_INSTQUEUE_REG_1__7__SCAN_IN | ~n97303;
  assign n64828 = ~n75033 | ~P1_P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n64830 = ~n64829 | ~n64828;
  assign n64843 = ~n64831 & ~n64830;
  assign n64834 = ~n97225 | ~P1_P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n64836 = ~P1_P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~n100072;
  assign n75052 = ~n65129;
  assign n64833 = ~n75052 | ~P1_P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n64841 = ~n64834 | ~n64833;
  assign n64839 = ~P1_P1_INSTQUEUE_REG_13__7__SCAN_IN | ~n97978;
  assign n64838 = ~P1_P1_INSTQUEUE_REG_2__7__SCAN_IN | ~n59938;
  assign n64840 = ~n64839 | ~n64838;
  assign n64842 = ~n64841 & ~n64840;
  assign n64844 = ~n64843 | ~n64842;
  assign n64847 = ~P1_P1_INSTQUEUE_REG_9__1__SCAN_IN | ~n97754;
  assign n64846 = ~P1_P1_INSTQUEUE_REG_10__1__SCAN_IN | ~n75052;
  assign n64851 = ~n64847 | ~n64846;
  assign n64849 = ~P1_P1_INSTQUEUE_REG_4__1__SCAN_IN | ~n59935;
  assign n64848 = ~P1_P1_INSTQUEUE_REG_5__1__SCAN_IN | ~n98034;
  assign n64850 = ~n64849 | ~n64848;
  assign n64859 = ~n64851 & ~n64850;
  assign n64853 = ~P1_P1_INSTQUEUE_REG_11__1__SCAN_IN | ~n97743;
  assign n64852 = ~P1_P1_INSTQUEUE_REG_15__1__SCAN_IN | ~n97895;
  assign n64857 = ~n64853 | ~n64852;
  assign n64855 = ~P1_P1_INSTQUEUE_REG_6__1__SCAN_IN | ~n97747;
  assign n64854 = ~P1_P1_INSTQUEUE_REG_14__1__SCAN_IN | ~n97746;
  assign n64856 = ~n64855 | ~n64854;
  assign n64858 = ~n64857 & ~n64856;
  assign n64875 = ~n64859 | ~n64858;
  assign n64861 = ~P1_P1_INSTQUEUE_REG_8__1__SCAN_IN | ~n97203;
  assign n64860 = ~P1_P1_INSTQUEUE_REG_1__1__SCAN_IN | ~n97303;
  assign n64865 = ~n64861 | ~n64860;
  assign n64863 = ~P1_P1_INSTQUEUE_REG_12__1__SCAN_IN | ~n97761;
  assign n64862 = ~P1_P1_INSTQUEUE_REG_0__1__SCAN_IN | ~n75033;
  assign n64864 = ~n64863 | ~n64862;
  assign n64873 = ~n64865 & ~n64864;
  assign n64867 = ~P1_P1_INSTQUEUE_REG_2__1__SCAN_IN | ~n59938;
  assign n64866 = ~P1_P1_INSTQUEUE_REG_7__1__SCAN_IN | ~n97185;
  assign n64871 = ~n64867 | ~n64866;
  assign n64869 = ~P1_P1_INSTQUEUE_REG_13__1__SCAN_IN | ~n97978;
  assign n64868 = ~P1_P1_INSTQUEUE_REG_3__1__SCAN_IN | ~n97225;
  assign n64870 = ~n64869 | ~n64868;
  assign n64872 = ~n64871 & ~n64870;
  assign n64874 = ~n64873 | ~n64872;
  assign n64877 = ~P1_P1_INSTQUEUE_REG_8__3__SCAN_IN | ~n97203;
  assign n64876 = ~P1_P1_INSTQUEUE_REG_0__3__SCAN_IN | ~n75033;
  assign n64881 = ~n64877 | ~n64876;
  assign n64879 = ~P1_P1_INSTQUEUE_REG_4__3__SCAN_IN | ~n59935;
  assign n64878 = ~P1_P1_INSTQUEUE_REG_15__3__SCAN_IN | ~n97895;
  assign n64880 = ~n64879 | ~n64878;
  assign n64889 = ~n64881 & ~n64880;
  assign n64883 = ~P1_P1_INSTQUEUE_REG_10__3__SCAN_IN | ~n75052;
  assign n64882 = ~P1_P1_INSTQUEUE_REG_7__3__SCAN_IN | ~n97185;
  assign n64887 = ~n64883 | ~n64882;
  assign n64885 = ~P1_P1_INSTQUEUE_REG_6__3__SCAN_IN | ~n97747;
  assign n64884 = ~P1_P1_INSTQUEUE_REG_14__3__SCAN_IN | ~n97746;
  assign n64886 = ~n64885 | ~n64884;
  assign n64888 = ~n64887 & ~n64886;
  assign n64905 = ~n64889 | ~n64888;
  assign n64891 = ~P1_P1_INSTQUEUE_REG_11__3__SCAN_IN | ~n97743;
  assign n64890 = ~P1_P1_INSTQUEUE_REG_3__3__SCAN_IN | ~n97225;
  assign n64895 = ~n64891 | ~n64890;
  assign n64893 = ~P1_P1_INSTQUEUE_REG_5__3__SCAN_IN | ~n97979;
  assign n64892 = ~P1_P1_INSTQUEUE_REG_1__3__SCAN_IN | ~n97303;
  assign n64894 = ~n64893 | ~n64892;
  assign n64903 = ~n64895 & ~n64894;
  assign n64897 = ~P1_P1_INSTQUEUE_REG_9__3__SCAN_IN | ~n97754;
  assign n64896 = ~P1_P1_INSTQUEUE_REG_2__3__SCAN_IN | ~n59938;
  assign n64901 = ~n64897 | ~n64896;
  assign n64899 = ~P1_P1_INSTQUEUE_REG_12__3__SCAN_IN | ~n97761;
  assign n64898 = ~P1_P1_INSTQUEUE_REG_13__3__SCAN_IN | ~n75055;
  assign n64900 = ~n64899 | ~n64898;
  assign n64902 = ~n64901 & ~n64900;
  assign n64904 = ~n64903 | ~n64902;
  assign n64907 = ~P1_P1_INSTQUEUE_REG_5__5__SCAN_IN | ~n97979;
  assign n64906 = ~P1_P1_INSTQUEUE_REG_0__5__SCAN_IN | ~n75033;
  assign n64911 = ~n64907 | ~n64906;
  assign n64909 = ~P1_P1_INSTQUEUE_REG_4__5__SCAN_IN | ~n59935;
  assign n64908 = ~P1_P1_INSTQUEUE_REG_15__5__SCAN_IN | ~n97895;
  assign n64910 = ~n64909 | ~n64908;
  assign n64935 = ~n64911 & ~n64910;
  assign n64913 = ~P1_P1_INSTQUEUE_REG_13__5__SCAN_IN | ~n97978;
  assign n64912 = ~P1_P1_INSTQUEUE_REG_2__5__SCAN_IN | ~n59938;
  assign n64915 = ~n64913 | ~n64912;
  assign n64914 = n97303 & P1_P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n64917 = ~n64915 & ~n64914;
  assign n64916 = ~n97203 | ~P1_P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n64933 = ~n64917 | ~n64916;
  assign n64919 = ~P1_P1_INSTQUEUE_REG_9__5__SCAN_IN | ~n97754;
  assign n64918 = ~P1_P1_INSTQUEUE_REG_10__5__SCAN_IN | ~n75052;
  assign n64923 = ~n64919 | ~n64918;
  assign n64921 = ~P1_P1_INSTQUEUE_REG_12__5__SCAN_IN | ~n97761;
  assign n64920 = ~P1_P1_INSTQUEUE_REG_3__5__SCAN_IN | ~n97225;
  assign n64922 = ~n64921 | ~n64920;
  assign n64931 = ~n64923 & ~n64922;
  assign n64925 = ~P1_P1_INSTQUEUE_REG_11__5__SCAN_IN | ~n97743;
  assign n64924 = ~P1_P1_INSTQUEUE_REG_7__5__SCAN_IN | ~n97185;
  assign n64929 = ~n64925 | ~n64924;
  assign n64927 = ~P1_P1_INSTQUEUE_REG_6__5__SCAN_IN | ~n97747;
  assign n64926 = ~P1_P1_INSTQUEUE_REG_14__5__SCAN_IN | ~n97746;
  assign n64928 = ~n64927 | ~n64926;
  assign n64930 = ~n64929 & ~n64928;
  assign n64932 = ~n64931 | ~n64930;
  assign n64934 = ~n64933 & ~n64932;
  assign n65062 = ~n76802 | ~n99221;
  assign n64936 = ~n99180 | ~n65062;
  assign n64967 = ~n64936 | ~n97556;
  assign n64938 = ~P1_P1_INSTQUEUE_REG_9__4__SCAN_IN | ~n97987;
  assign n64937 = ~P1_P1_INSTQUEUE_REG_15__4__SCAN_IN | ~n97895;
  assign n64942 = ~n64938 | ~n64937;
  assign n64940 = ~P1_P1_INSTQUEUE_REG_11__4__SCAN_IN | ~n98007;
  assign n97979 = ~n60790;
  assign n64939 = ~P1_P1_INSTQUEUE_REG_5__4__SCAN_IN | ~n97979;
  assign n64941 = ~n64940 | ~n64939;
  assign n64950 = ~n64942 & ~n64941;
  assign n64944 = ~P1_P1_INSTQUEUE_REG_12__4__SCAN_IN | ~n98011;
  assign n64943 = ~P1_P1_INSTQUEUE_REG_3__4__SCAN_IN | ~n97988;
  assign n64948 = ~n64944 | ~n64943;
  assign n64946 = ~P1_P1_INSTQUEUE_REG_6__4__SCAN_IN | ~n97991;
  assign n64945 = ~P1_P1_INSTQUEUE_REG_14__4__SCAN_IN | ~n59936;
  assign n64947 = ~n64946 | ~n64945;
  assign n64949 = ~n64948 & ~n64947;
  assign n64966 = ~n64950 | ~n64949;
  assign n64952 = ~P1_P1_INSTQUEUE_REG_8__4__SCAN_IN | ~n97982;
  assign n64951 = ~P1_P1_INSTQUEUE_REG_10__4__SCAN_IN | ~n98002;
  assign n64956 = ~n64952 | ~n64951;
  assign n64954 = ~P1_P1_INSTQUEUE_REG_2__4__SCAN_IN | ~n98008;
  assign n64953 = ~P1_P1_INSTQUEUE_REG_0__4__SCAN_IN | ~n59937;
  assign n64955 = ~n64954 | ~n64953;
  assign n64964 = ~n64956 & ~n64955;
  assign n64958 = ~P1_P1_INSTQUEUE_REG_7__4__SCAN_IN | ~n97185;
  assign n64957 = ~P1_P1_INSTQUEUE_REG_1__4__SCAN_IN | ~n97999;
  assign n64962 = ~n64958 | ~n64957;
  assign n64960 = ~P1_P1_INSTQUEUE_REG_4__4__SCAN_IN | ~n59935;
  assign n64959 = ~P1_P1_INSTQUEUE_REG_13__4__SCAN_IN | ~n97978;
  assign n64961 = ~n64960 | ~n64959;
  assign n64963 = ~n64962 & ~n64961;
  assign n64965 = ~n64964 | ~n64963;
  assign n96898 = ~n64966 & ~n64965;
  assign n64999 = ~n64967 | ~n96898;
  assign n64969 = ~P1_P1_INSTQUEUE_REG_8__6__SCAN_IN | ~n97203;
  assign n64968 = ~P1_P1_INSTQUEUE_REG_3__6__SCAN_IN | ~n97225;
  assign n64973 = ~n64969 | ~n64968;
  assign n64971 = ~P1_P1_INSTQUEUE_REG_9__6__SCAN_IN | ~n97754;
  assign n64970 = ~P1_P1_INSTQUEUE_REG_13__6__SCAN_IN | ~n97978;
  assign n64972 = ~n64971 | ~n64970;
  assign n64981 = ~n64973 & ~n64972;
  assign n64975 = ~P1_P1_INSTQUEUE_REG_6__6__SCAN_IN | ~n97747;
  assign n64974 = ~P1_P1_INSTQUEUE_REG_1__6__SCAN_IN | ~n97303;
  assign n64979 = ~n64975 | ~n64974;
  assign n64977 = ~P1_P1_INSTQUEUE_REG_14__6__SCAN_IN | ~n97746;
  assign n64976 = ~P1_P1_INSTQUEUE_REG_5__6__SCAN_IN | ~n98034;
  assign n64978 = ~n64977 | ~n64976;
  assign n64980 = ~n64979 & ~n64978;
  assign n64997 = n64981 & n64980;
  assign n64983 = ~P1_P1_INSTQUEUE_REG_11__6__SCAN_IN | ~n97743;
  assign n64982 = ~P1_P1_INSTQUEUE_REG_7__6__SCAN_IN | ~n97185;
  assign n64987 = ~n64983 | ~n64982;
  assign n64985 = ~P1_P1_INSTQUEUE_REG_10__6__SCAN_IN | ~n75052;
  assign n64984 = ~P1_P1_INSTQUEUE_REG_0__6__SCAN_IN | ~n75033;
  assign n64986 = ~n64985 | ~n64984;
  assign n64995 = ~n64987 & ~n64986;
  assign n64989 = ~P1_P1_INSTQUEUE_REG_4__6__SCAN_IN | ~n59935;
  assign n64988 = ~P1_P1_INSTQUEUE_REG_2__6__SCAN_IN | ~n59938;
  assign n64993 = ~n64989 | ~n64988;
  assign n64991 = ~P1_P1_INSTQUEUE_REG_15__6__SCAN_IN | ~n97895;
  assign n64990 = ~P1_P1_INSTQUEUE_REG_12__6__SCAN_IN | ~n97761;
  assign n64992 = ~n64991 | ~n64990;
  assign n64994 = ~n64993 & ~n64992;
  assign n64996 = n64995 & n64994;
  assign n65071 = ~n99178;
  assign n64998 = ~n97620 | ~n65071;
  assign n65066 = ~n64999 | ~n64998;
  assign n65001 = ~P1_P1_INSTQUEUE_REG_11__0__SCAN_IN | ~n97743;
  assign n65000 = ~P1_P1_INSTQUEUE_REG_5__0__SCAN_IN | ~n98034;
  assign n65005 = ~n65001 | ~n65000;
  assign n65003 = ~P1_P1_INSTQUEUE_REG_8__0__SCAN_IN | ~n97203;
  assign n65002 = ~P1_P1_INSTQUEUE_REG_7__0__SCAN_IN | ~n97185;
  assign n65004 = ~n65003 | ~n65002;
  assign n65013 = ~n65005 & ~n65004;
  assign n65007 = ~P1_P1_INSTQUEUE_REG_4__0__SCAN_IN | ~n59935;
  assign n65006 = ~P1_P1_INSTQUEUE_REG_13__0__SCAN_IN | ~n97978;
  assign n65011 = ~n65007 | ~n65006;
  assign n65009 = ~P1_P1_INSTQUEUE_REG_6__0__SCAN_IN | ~n97747;
  assign n65008 = ~P1_P1_INSTQUEUE_REG_14__0__SCAN_IN | ~n97746;
  assign n65010 = ~n65009 | ~n65008;
  assign n65012 = ~n65011 & ~n65010;
  assign n65029 = ~n65013 | ~n65012;
  assign n65015 = ~P1_P1_INSTQUEUE_REG_9__0__SCAN_IN | ~n97754;
  assign n65014 = ~P1_P1_INSTQUEUE_REG_15__0__SCAN_IN | ~n97895;
  assign n65019 = ~n65015 | ~n65014;
  assign n65017 = ~P1_P1_INSTQUEUE_REG_3__0__SCAN_IN | ~n97225;
  assign n65016 = ~P1_P1_INSTQUEUE_REG_0__0__SCAN_IN | ~n75033;
  assign n65018 = ~n65017 | ~n65016;
  assign n65027 = ~n65019 & ~n65018;
  assign n65021 = ~P1_P1_INSTQUEUE_REG_12__0__SCAN_IN | ~n97761;
  assign n65020 = ~P1_P1_INSTQUEUE_REG_10__0__SCAN_IN | ~n75052;
  assign n65025 = ~n65021 | ~n65020;
  assign n65023 = ~P1_P1_INSTQUEUE_REG_2__0__SCAN_IN | ~n59938;
  assign n65022 = ~P1_P1_INSTQUEUE_REG_1__0__SCAN_IN | ~n97303;
  assign n65024 = ~n65023 | ~n65022;
  assign n65026 = ~n65025 & ~n65024;
  assign n65028 = ~n65027 | ~n65026;
  assign n98214 = ~n99180;
  assign n99186 = ~n96899 | ~n98214;
  assign n65031 = ~P1_P1_INSTQUEUE_REG_4__2__SCAN_IN | ~n59935;
  assign n65030 = ~P1_P1_INSTQUEUE_REG_7__2__SCAN_IN | ~n97185;
  assign n65035 = ~n65031 | ~n65030;
  assign n65033 = ~P1_P1_INSTQUEUE_REG_10__2__SCAN_IN | ~n75052;
  assign n65032 = ~P1_P1_INSTQUEUE_REG_3__2__SCAN_IN | ~n97225;
  assign n65034 = ~n65033 | ~n65032;
  assign n65043 = ~n65035 & ~n65034;
  assign n65037 = ~P1_P1_INSTQUEUE_REG_6__2__SCAN_IN | ~n97747;
  assign n65036 = ~P1_P1_INSTQUEUE_REG_2__2__SCAN_IN | ~n59938;
  assign n65041 = ~n65037 | ~n65036;
  assign n65039 = ~P1_P1_INSTQUEUE_REG_9__2__SCAN_IN | ~n97754;
  assign n65038 = ~P1_P1_INSTQUEUE_REG_14__2__SCAN_IN | ~n97746;
  assign n65040 = ~n65039 | ~n65038;
  assign n65042 = ~n65041 & ~n65040;
  assign n65059 = ~n65043 | ~n65042;
  assign n65045 = ~P1_P1_INSTQUEUE_REG_8__2__SCAN_IN | ~n97203;
  assign n65044 = ~P1_P1_INSTQUEUE_REG_5__2__SCAN_IN | ~n97979;
  assign n65049 = ~n65045 | ~n65044;
  assign n65047 = ~P1_P1_INSTQUEUE_REG_13__2__SCAN_IN | ~n97978;
  assign n65046 = ~P1_P1_INSTQUEUE_REG_0__2__SCAN_IN | ~n75033;
  assign n65048 = ~n65047 | ~n65046;
  assign n65057 = ~n65049 & ~n65048;
  assign n65051 = ~P1_P1_INSTQUEUE_REG_15__2__SCAN_IN | ~n97895;
  assign n65050 = ~P1_P1_INSTQUEUE_REG_1__2__SCAN_IN | ~n97303;
  assign n65055 = ~n65051 | ~n65050;
  assign n65053 = ~P1_P1_INSTQUEUE_REG_11__2__SCAN_IN | ~n97743;
  assign n65052 = ~P1_P1_INSTQUEUE_REG_12__2__SCAN_IN | ~n97761;
  assign n65054 = ~n65053 | ~n65052;
  assign n65056 = ~n65055 & ~n65054;
  assign n65058 = ~n65057 | ~n65056;
  assign n65060 = ~n99186 | ~n99201;
  assign n65061 = ~n65060 | ~n65071;
  assign n65120 = ~n99221 | ~n99179;
  assign n65126 = ~n65120;
  assign n99191 = ~n65126 | ~n96898;
  assign n65064 = ~n65061 | ~n99191;
  assign n65063 = ~n96899 & ~n65062;
  assign n65065 = ~n65064 & ~n65063;
  assign n65079 = ~n65066 | ~n65065;
  assign n100065 = ~n97620 | ~n65120;
  assign n97651 = ~n100065;
  assign n98071 = ~n96899;
  assign n100471 = ~n99180 | ~n98071;
  assign n99197 = ~n97651 & ~n100471;
  assign n65085 = ~n99179 | ~n96898;
  assign n65067 = n65085 & n96896;
  assign n65068 = ~n99197 & ~n65067;
  assign n65069 = ~n65068 | ~n99201;
  assign n65070 = ~n76802;
  assign n65077 = ~n65069 | ~n65070;
  assign n65122 = ~n98071 & ~n98214;
  assign n65074 = n65070 | n65122;
  assign n65072 = ~n65085 | ~n65071;
  assign n65073 = ~n96899 | ~n65072;
  assign n65075 = ~n65074 | ~n65073;
  assign n65076 = ~n65075 | ~n99201;
  assign n65078 = ~n65077 | ~n65076;
  assign n96897 = ~n76802 | ~n99201;
  assign n99214 = ~n96895 & ~n96897;
  assign n65080 = ~n99214;
  assign n100066 = ~n100130 | ~n65080;
  assign n100481 = ~P2_P1_ADS_N_REG_SCAN_IN | ~P1_READY11_REG_SCAN_IN;
  assign n96146 = ~n96898 | ~n99178;
  assign n65081 = ~n76802 | ~n96899;
  assign n65083 = ~n96146 & ~n65081;
  assign n65082 = ~n97556 & ~n99201;
  assign n96131 = ~n65083 | ~n65082;
  assign n100107 = ~n98214 & ~n96131;
  assign n65088 = ~n100481 | ~n100107;
  assign n65084 = ~n97556 & ~n76802;
  assign n99194 = ~n99201 | ~n65084;
  assign n65086 = ~n65085 & ~n99194;
  assign n96132 = ~n96896 | ~n65086;
  assign n96893 = ~n98071 | ~n98214;
  assign n65087 = ~n96132 & ~n96893;
  assign n98211 = ~n65087 | ~n100481;
  assign n65111 = ~n65088 | ~n98211;
  assign n100023 = ~P1_P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n65092 = ~P1_P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~n100023;
  assign n65103 = ~P1_P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n100072;
  assign n65090 = ~P1_P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n65089;
  assign n65091 = ~n65103 & ~n65090;
  assign n65093 = ~n65092 & ~n65091;
  assign n65094 = ~P1_P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ P1_P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n65113 = n65093 ^ n65094;
  assign n65100 = ~P1_P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~n100044;
  assign n100141 = ~P1_P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n65096 = ~P1_P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~n100141;
  assign n65095 = ~n65094 | ~n65093;
  assign n65098 = ~n65096 | ~n65095;
  assign n65105 = ~n70278 | ~n65098;
  assign n65097 = ~n65100 | ~n65105;
  assign n65102 = ~P1_P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n65097;
  assign n65099 = ~n70278 & ~n65098;
  assign n65106 = ~n65100 & ~n65099;
  assign n65101 = ~n65106;
  assign n65116 = ~n65102 | ~n65101;
  assign n96143 = ~n65113 | ~n65116;
  assign n65112 = n100023 ^ P1_P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n65104 = ~n65112 ^ n65103;
  assign n65110 = ~n96143 & ~n65104;
  assign n65107 = ~n65105 | ~n100136;
  assign n65109 = ~n65107 | ~n65106;
  assign n65108 = ~P1_P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n100044;
  assign n65118 = ~n65109 | ~n65108;
  assign n65124 = ~n65111 | ~n100048;
  assign n100076 = ~P1_P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n96141 = ~n100076 ^ n100072;
  assign n65115 = ~n65112 | ~n96141;
  assign n65114 = ~n65113;
  assign n65117 = ~n65115 | ~n65114;
  assign n65119 = n65117 & n65116;
  assign n100046 = ~n99199;
  assign n65121 = ~n99194;
  assign n99188 = ~n96898 & ~n65120;
  assign n99216 = ~n65121 | ~n99188;
  assign n96892 = ~n100046 & ~n99216;
  assign n65123 = ~n65122 | ~n96892;
  assign n100085 = ~n65124 | ~n65123;
  assign n65125 = ~n99213 & ~n100085;
  assign n71418 = ~n97636;
  assign n97564 = ~n71418 & ~n97648;
  assign n98034 = ~n60790;
  assign n98037 = ~n64817;
  assign n97591 = n97723 & n96896;
  assign n97630 = ~n97591;
  assign n97604 = ~P1_P1_EAX_REG_11__SCAN_IN | ~P1_P1_EAX_REG_10__SCAN_IN;
  assign n98337 = ~P1_P1_EAX_REG_9__SCAN_IN;
  assign n98326 = ~P1_P1_EAX_REG_7__SCAN_IN;
  assign n98291 = ~P1_P1_EAX_REG_0__SCAN_IN;
  assign n65168 = ~P1_P1_EAX_REG_2__SCAN_IN | ~P1_P1_EAX_REG_1__SCAN_IN;
  assign n97846 = ~n98291 & ~n65168;
  assign n65170 = ~P1_P1_EAX_REG_3__SCAN_IN | ~n97846;
  assign n65169 = ~P1_P1_EAX_REG_5__SCAN_IN | ~P1_P1_EAX_REG_4__SCAN_IN;
  assign n97808 = ~n65170 & ~n65169;
  assign n97730 = ~P1_P1_EAX_REG_6__SCAN_IN | ~n97808;
  assign n65171 = ~n98326 & ~n97730;
  assign n97708 = ~P1_P1_EAX_REG_8__SCAN_IN | ~n65171;
  assign n97698 = ~n98337 & ~n97708;
  assign n98362 = ~P1_P1_EAX_REG_14__SCAN_IN;
  assign n98357 = ~P1_P1_EAX_REG_13__SCAN_IN;
  assign n97655 = ~n98362 & ~n98357;
  assign n97621 = P1_P1_EAX_REG_15__SCAN_IN & n97655;
  assign n65173 = ~P1_P1_EAX_REG_16__SCAN_IN | ~n97621;
  assign n65172 = ~P1_P1_EAX_REG_12__SCAN_IN | ~P1_P1_EAX_REG_17__SCAN_IN;
  assign n97605 = ~n65173 & ~n65172;
  assign n65174 = ~n97698 | ~n97605;
  assign n65175 = ~n97604 & ~n65174;
  assign n97595 = ~P1_P1_EAX_REG_18__SCAN_IN | ~n65175;
  assign n97555 = ~P1_P1_EAX_REG_20__SCAN_IN | ~P1_P1_EAX_REG_19__SCAN_IN;
  assign n71742 = ~n97595 & ~n97555;
  assign n98024 = ~n97556 | ~n97928;
  assign n67201 = ~n67193 | ~n67192;
  assign n67196 = n67195 & n67194;
  assign n67199 = ~n67197 | ~n67196;
  assign n67200 = ~n67199 | ~n67198;
  assign n68985 = ~n67201 | ~n67200;
  assign n68983 = ~n71659 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n67202 = ~n68983;
  assign n67914 = ~n76076 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n67918 = ~n76046 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n67204 = ~n67914 ^ n67918;
  assign n67366 = ~n67915 ^ n67204;
  assign n67206 = ~n67207 | ~n67208;
  assign n67210 = ~n67207;
  assign n67209 = ~n67208;
  assign n67211 = ~n67210 | ~n67209;
  assign n67217 = ~n67213 | ~n64503;
  assign n67218 = ~n67217 | ~n67216;
  assign n67222 = ~n67224 | ~n67223;
  assign n67747 = n76067 & P4_DATAO_REG_5__SCAN_IN;
  assign n67234 = ~n67228 | ~n67227;
  assign n67231 = n67234 & n67226;
  assign n67230 = ~n67233 | ~n67229;
  assign n67232 = ~n67231 | ~n67230;
  assign n67235 = ~n67234 | ~n59980;
  assign n67237 = ~n67236 | ~n67235;
  assign n67750 = ~n76064 & ~n76061;
  assign n67246 = ~n67241 | ~n67240;
  assign n67245 = ~n67244 | ~n67243;
  assign n68799 = ~n64350 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n67345 = ~n68802 ^ n68800;
  assign n67249 = ~n67299;
  assign n67253 = ~n67250 ^ n67249;
  assign n67252 = ~n67251;
  assign n67254 = ~n67253 | ~n67252;
  assign n67844 = ~n63603 & ~n59984;
  assign n67307 = ~n67845 ^ n67844;
  assign n67259 = ~n67256;
  assign n67258 = ~n67257;
  assign n67260 = ~n67259 | ~n67258;
  assign n67263 = ~n67261;
  assign n67264 = ~n67263 | ~n67262;
  assign n75996 = ~P4_DATAO_REG_23__SCAN_IN;
  assign n67270 = ~DIN_0_ | ~P4_DATAO_REG_23__SCAN_IN;
  assign n67265 = ~n60178 | ~n67270;
  assign n67267 = P4_DATAO_REG_22__SCAN_IN & P4_DATAO_REG_23__SCAN_IN;
  assign n68849 = ~n74276 | ~n67267;
  assign n68857 = ~n67268 | ~n68849;
  assign n68858 = ~n59870 | ~P4_DATAO_REG_21__SCAN_IN;
  assign n67269 = ~n68856;
  assign n67814 = ~n68858 | ~n67270;
  assign n68845 = ~n59870 | ~P4_DATAO_REG_23__SCAN_IN;
  assign n67271 = ~n67814 | ~n68845;
  assign n67805 = n67271 | n68856;
  assign n67813 = ~n74882 & ~n74820;
  assign n67823 = ~n59909 | ~P4_DATAO_REG_19__SCAN_IN;
  assign n67832 = ~n74835 | ~P4_DATAO_REG_18__SCAN_IN;
  assign n67277 = ~n67823 ^ n67832;
  assign n67280 = ~n67278;
  assign n67281 = ~n67280 | ~n67279;
  assign n67836 = ~n63005 | ~P4_DATAO_REG_17__SCAN_IN;
  assign n67304 = ~n67837 ^ n67836;
  assign n67286 = ~n67283;
  assign n67285 = ~n67284;
  assign n67288 = ~n67286 | ~n67285;
  assign n67290 = n67288 & n67287;
  assign n67302 = ~n67290 | ~n67289;
  assign n67294 = ~n67292 | ~n67291;
  assign n67298 = ~n67294 | ~n67293;
  assign n67297 = ~n67296 | ~n67295;
  assign n67300 = ~n67298 | ~n67297;
  assign n67301 = ~n67300 | ~n67299;
  assign n67303 = n67302 & n67301;
  assign n67305 = ~n67304 | ~n67303;
  assign n67308 = ~n67307 | ~n67306;
  assign n67316 = ~n67309 | ~n67310;
  assign n67311 = ~n67310;
  assign n67314 = ~n67312 | ~n67311;
  assign n67315 = ~n67314 | ~n67313;
  assign n67852 = ~n76062 & ~n60217;
  assign n67317 = ~n67852;
  assign n67322 = ~n67319 | ~n67318;
  assign n67861 = ~n74798 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n67773 = ~n59930 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n67864 = ~n76000 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n67326 = ~n67773 ^ n67864;
  assign n67759 = ~n71230 & ~n74360;
  assign n67770 = ~n67332 | ~n67329;
  assign n67337 = ~n67333;
  assign n67336 = ~n67335 | ~n67334;
  assign n67340 = ~n67339 | ~n67338;
  assign n67344 = ~n67343 | ~n67342;
  assign n67349 = ~n67347 | ~n67346;
  assign n67357 = ~n67349 | ~n67348;
  assign n67352 = ~n67351 | ~n67350;
  assign n67355 = ~n67353 | ~n67352;
  assign n67356 = ~n67355 | ~n67354;
  assign n67363 = ~n67361 | ~n67743;
  assign n68959 = ~n76043 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n67373 = ~n67368 | ~n67367;
  assign n67370 = ~n59992 & ~n67369;
  assign n67372 = ~n67371 | ~n67370;
  assign n67376 = ~n67375 | ~n67374;
  assign n67378 = ~n67377 | ~n67376;
  assign n76055 = ~n76028 | ~DIN_23_;
  assign n67930 = ~n71171 & ~n76055;
  assign n67383 = n67382 & n67381;
  assign n67385 = ~n67389 | ~n67383;
  assign n67386 = ~n76046;
  assign n67388 = n67387 | n67386;
  assign n67391 = ~n67389 | ~n67388;
  assign n67397 = ~P1_P1_INSTQUEUE_REG_8__0__SCAN_IN | ~n59935;
  assign n67396 = ~P1_P1_INSTQUEUE_REG_11__0__SCAN_IN | ~n97185;
  assign n67401 = ~n67397 | ~n67396;
  assign n67399 = ~P1_P1_INSTQUEUE_REG_13__0__SCAN_IN | ~n97754;
  assign n67398 = ~P1_P1_INSTQUEUE_REG_1__0__SCAN_IN | ~n75055;
  assign n67400 = ~n67399 | ~n67398;
  assign n67409 = ~n67401 & ~n67400;
  assign n67403 = ~P1_P1_INSTQUEUE_REG_7__0__SCAN_IN | ~n97225;
  assign n67402 = ~P1_P1_INSTQUEUE_REG_9__0__SCAN_IN | ~n97979;
  assign n67407 = ~n67403 | ~n67402;
  assign n67405 = ~P1_P1_INSTQUEUE_REG_10__0__SCAN_IN | ~n97747;
  assign n67404 = ~P1_P1_INSTQUEUE_REG_2__0__SCAN_IN | ~n97746;
  assign n67406 = ~n67405 | ~n67404;
  assign n67408 = ~n67407 & ~n67406;
  assign n67425 = ~n67409 | ~n67408;
  assign n67411 = ~P1_P1_INSTQUEUE_REG_3__0__SCAN_IN | ~n97895;
  assign n67410 = ~P1_P1_INSTQUEUE_REG_5__0__SCAN_IN | ~n97303;
  assign n67415 = ~n67411 | ~n67410;
  assign n67413 = ~P1_P1_INSTQUEUE_REG_12__0__SCAN_IN | ~n97203;
  assign n67412 = ~P1_P1_INSTQUEUE_REG_4__0__SCAN_IN | ~n75033;
  assign n67414 = ~n67413 | ~n67412;
  assign n67423 = ~n67415 & ~n67414;
  assign n67417 = ~P1_P1_INSTQUEUE_REG_0__0__SCAN_IN | ~n97761;
  assign n67416 = ~P1_P1_INSTQUEUE_REG_14__0__SCAN_IN | ~n75052;
  assign n67421 = ~n67417 | ~n67416;
  assign n67419 = ~P1_P1_INSTQUEUE_REG_15__0__SCAN_IN | ~n97743;
  assign n67418 = ~P1_P1_INSTQUEUE_REG_6__0__SCAN_IN | ~n59938;
  assign n67420 = ~n67419 | ~n67418;
  assign n67422 = ~n67421 & ~n67420;
  assign n67424 = ~n67423 | ~n67422;
  assign n67943 = ~n67425 & ~n67424;
  assign n67427 = ~P1_P1_INSTQUEUE_REG_15__7__SCAN_IN | ~n97761;
  assign n67426 = ~n59938 | ~P1_P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n67431 = ~n67427 | ~n67426;
  assign n67429 = ~n75052 | ~P1_P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n67428 = ~n59935 | ~P1_P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n67430 = ~n67429 | ~n67428;
  assign n67439 = ~n67431 & ~n67430;
  assign n67433 = ~P1_P1_INSTQUEUE_REG_14__7__SCAN_IN | ~n97743;
  assign n67432 = ~P1_P1_INSTQUEUE_REG_11__7__SCAN_IN | ~n97203;
  assign n67437 = ~n67433 | ~n67432;
  assign n67435 = ~P1_P1_INSTQUEUE_REG_9__7__SCAN_IN | ~n98037;
  assign n67434 = ~n97746 | ~P1_P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n67436 = ~n67435 | ~n67434;
  assign n67438 = ~n67437 & ~n67436;
  assign n67455 = ~n67439 | ~n67438;
  assign n67441 = ~n97895 | ~P1_P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n67440 = ~P1_P1_INSTQUEUE_REG_10__7__SCAN_IN | ~n97185;
  assign n67445 = ~n67441 | ~n67440;
  assign n67443 = ~n97754 | ~P1_P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n67442 = ~n75055 | ~P1_P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n67444 = ~n67443 | ~n67442;
  assign n67453 = ~n67445 & ~n67444;
  assign n67447 = ~P1_P1_INSTQUEUE_REG_6__7__SCAN_IN | ~n97225;
  assign n67446 = ~P1_P1_INSTQUEUE_REG_4__7__SCAN_IN | ~n97303;
  assign n67451 = ~n67447 | ~n67446;
  assign n67449 = ~P1_P1_INSTQUEUE_REG_8__7__SCAN_IN | ~n97979;
  assign n67448 = ~P1_P1_INSTQUEUE_REG_3__7__SCAN_IN | ~n75033;
  assign n67450 = ~n67449 | ~n67448;
  assign n67452 = ~n67451 & ~n67450;
  assign n67454 = ~n67453 | ~n67452;
  assign n67942 = ~n67455 & ~n67454;
  assign n67732 = ~n68989 | ~n68985;
  assign n67734 = ~n68996 | ~n68995;
  assign n68994 = ~n71188 & ~n76055;
  assign n67733 = ~n68994;
  assign n67740 = ~n68767 | ~n67916;
  assign n67736 = ~n76043;
  assign n67737 = ~n67914;
  assign n67739 = ~n68768 | ~n68769;
  assign n67742 = n67743 | n67744;
  assign n67746 = ~n67742 | ~n67741;
  assign n67745 = ~n67744 | ~n67743;
  assign n67749 = ~n67748 | ~n67747;
  assign n68950 = ~n76043 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n68793 = ~n76051 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n67754 = ~n67753;
  assign n67757 = ~n67756 | ~n67752;
  assign n68936 = ~n64350 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n67758 = ~n67762;
  assign n67765 = ~n67760 | ~n67759;
  assign n67763 = ~n67761;
  assign n67764 = ~n67763 | ~n67762;
  assign n67769 = ~n67765 | ~n67764;
  assign n67767 = ~n67769;
  assign n67768 = ~n71230 & ~n74367;
  assign n67766 = ~n67768;
  assign n68825 = ~n67767 | ~n67766;
  assign n68827 = ~n67769 | ~n67768;
  assign n67772 = ~n67770;
  assign n67774 = ~n67865 ^ n67864;
  assign n67775 = ~n67774 | ~n67773;
  assign n67874 = ~n68927 ^ n68928;
  assign n76032 = ~P4_DATAO_REG_24__SCAN_IN;
  assign n67782 = ~n68849 ^ n68848;
  assign n67778 = ~n75996 | ~n74277;
  assign n67779 = ~n75996 & ~n63317;
  assign n67783 = ~n59870 | ~P4_DATAO_REG_22__SCAN_IN;
  assign n67785 = ~n67784 | ~n67783;
  assign n67786 = ~n68856 | ~n64706;
  assign n67787 = ~n67786 | ~n62954;
  assign n67793 = n67787 | n68857;
  assign n67788 = ~n63724 & ~n74820;
  assign n67789 = ~n63724 | ~n74820;
  assign n67794 = n67789 & P4_DATAO_REG_21__SCAN_IN;
  assign n67790 = ~n68856 | ~n67794;
  assign n67792 = ~n67791 | ~n67790;
  assign n67798 = ~n67793 | ~n67792;
  assign n67795 = ~n68856 | ~n74820;
  assign n67796 = ~n67795 | ~n67794;
  assign n67797 = n67796 & n68857;
  assign n68863 = ~n67800 | ~n67799;
  assign n67802 = ~n67799;
  assign n67803 = ~n67802 | ~n67801;
  assign n68868 = ~n68863 | ~n67803;
  assign n67804 = ~n67813;
  assign n67806 = n67805 & n67804;
  assign n67810 = ~n67807 | ~n67806;
  assign n67809 = ~n67808;
  assign n67819 = ~n67810 | ~n67809;
  assign n67811 = ~n68856 | ~n67813;
  assign n67817 = n67812 | n67811;
  assign n67815 = ~n67814 | ~n67813;
  assign n67816 = n67815 | n68856;
  assign n67818 = n67817 & n67816;
  assign n68867 = ~n67819 | ~n67818;
  assign n67821 = ~n68868 ^ n68867;
  assign n67820 = ~n74882 & ~n59912;
  assign n68871 = ~n67821 | ~n67820;
  assign n68876 = ~n74835 | ~P4_DATAO_REG_19__SCAN_IN;
  assign n67826 = ~n67823;
  assign n67825 = ~n67824;
  assign n67828 = ~n67827 | ~n67826;
  assign n67834 = ~n67830 | ~n67829;
  assign n67835 = ~n63005 | ~P4_DATAO_REG_18__SCAN_IN;
  assign n67838 = n67837 | n67836;
  assign n68881 = ~n74361 & ~n59984;
  assign n67839 = ~n67842;
  assign n67843 = ~n67842 | ~n67841;
  assign n67846 = ~n67845 | ~n67844;
  assign n68886 = ~n63296 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n68889 = ~n67849 | ~n67848;
  assign n67851 = ~n67848;
  assign n67850 = ~n67849;
  assign n67858 = ~n67853 | ~n67852;
  assign n67856 = ~n67854;
  assign n67857 = ~n67856 | ~n67855;
  assign n68892 = ~n76062 & ~n76012;
  assign n67863 = ~n67860 | ~n67859;
  assign n70110 = ~n67863 | ~n67862;
  assign n70113 = ~n76000 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n68920 = ~n59930 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n67873 = ~n68921 ^ n68920;
  assign n67871 = n67865 | n67864;
  assign n67869 = ~n67866;
  assign n67868 = ~n67867;
  assign n67870 = ~n67869 | ~n67868;
  assign n68826 = ~n67874 ^ n68926;
  assign n68810 = ~n67875 | ~n68799;
  assign n68809 = ~n68798 | ~n68802;
  assign n68807 = ~n63929 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n67876 = ~n68816;
  assign n67877 = ~n68807 ^ n67876;
  assign n67879 = ~n67878 ^ n67877;
  assign n67885 = ~n68821 ^ n67879;
  assign n67882 = ~n67881 | ~n67880;
  assign n67887 = n67886 & n67890;
  assign n67892 = ~n67889 | ~n67888;
  assign n67894 = ~n67892 | ~n67891;
  assign n67893 = n76067 & P4_DATAO_REG_6__SCAN_IN;
  assign n68780 = ~n67894 & ~n67893;
  assign n68783 = ~n67894 | ~n67893;
  assign n67895 = ~n68781 | ~n68783;
  assign n67910 = ~n68956;
  assign n67901 = ~n76076 | ~n76043;
  assign n67896 = ~n76076 & ~n76043;
  assign n67904 = ~n67896 & ~n74771;
  assign n67900 = ~n67899 | ~n67898;
  assign n67909 = ~n67900 | ~n68957;
  assign n67903 = ~n67902 | ~n67901;
  assign n67905 = ~n67904;
  assign n67906 = ~n60836 | ~n67905;
  assign n67908 = n67907 & n67906;
  assign n67912 = ~n71397 & ~n76044;
  assign n68973 = n67911 | n67912;
  assign n68975 = ~n67911;
  assign n67922 = ~n68973 | ~n68979;
  assign n67917 = ~n67915 ^ n67914;
  assign n67919 = ~n67916 ^ n67917;
  assign n67924 = ~n71171 & ~n76063;
  assign n67926 = ~n67923;
  assign n67925 = ~n67924;
  assign n67934 = ~n67928 | ~n67935;
  assign n67932 = ~n67929;
  assign n67931 = ~n67930;
  assign n67938 = ~n67934 | ~n67933;
  assign n69047 = ~n67943 & ~n67942;
  assign n67945 = ~P1_P1_INSTQUEUE_REG_15__1__SCAN_IN | ~n97743;
  assign n67944 = ~P1_P1_INSTQUEUE_REG_9__1__SCAN_IN | ~n98034;
  assign n67949 = ~n67945 | ~n67944;
  assign n67947 = ~P1_P1_INSTQUEUE_REG_8__1__SCAN_IN | ~n59935;
  assign n67946 = ~P1_P1_INSTQUEUE_REG_0__1__SCAN_IN | ~n97761;
  assign n67948 = ~n67947 | ~n67946;
  assign n67973 = ~n67949 & ~n67948;
  assign n67951 = ~P1_P1_INSTQUEUE_REG_11__1__SCAN_IN | ~n97185;
  assign n67950 = ~P1_P1_INSTQUEUE_REG_4__1__SCAN_IN | ~n75033;
  assign n67953 = ~n67951 | ~n67950;
  assign n67952 = n97303 & P1_P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n67955 = ~n67953 & ~n67952;
  assign n67954 = ~n97754 | ~P1_P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n67971 = ~n67955 | ~n67954;
  assign n67957 = ~P1_P1_INSTQUEUE_REG_3__1__SCAN_IN | ~n97895;
  assign n67956 = ~P1_P1_INSTQUEUE_REG_6__1__SCAN_IN | ~n59938;
  assign n67961 = ~n67957 | ~n67956;
  assign n67959 = ~P1_P1_INSTQUEUE_REG_12__1__SCAN_IN | ~n97203;
  assign n67958 = ~P1_P1_INSTQUEUE_REG_7__1__SCAN_IN | ~n97225;
  assign n67960 = ~n67959 | ~n67958;
  assign n67969 = ~n67961 & ~n67960;
  assign n67963 = ~P1_P1_INSTQUEUE_REG_2__1__SCAN_IN | ~n59936;
  assign n67962 = ~P1_P1_INSTQUEUE_REG_14__1__SCAN_IN | ~n75052;
  assign n67967 = ~n67963 | ~n67962;
  assign n67965 = ~P1_P1_INSTQUEUE_REG_10__1__SCAN_IN | ~n98037;
  assign n67964 = ~P1_P1_INSTQUEUE_REG_1__1__SCAN_IN | ~n75055;
  assign n67966 = ~n67965 | ~n67964;
  assign n67968 = ~n67967 & ~n67966;
  assign n67970 = ~n67969 | ~n67968;
  assign n67972 = ~n67971 & ~n67970;
  assign n69046 = ~n67973 | ~n67972;
  assign n68770 = ~n68769 | ~n68776;
  assign n68772 = ~n68771 & ~n68770;
  assign n68784 = ~n68782 | ~n68781;
  assign n70000 = n76043 & P4_DATAO_REG_6__SCAN_IN;
  assign n70179 = ~n70000;
  assign n70188 = n76076 & P4_DATAO_REG_5__SCAN_IN;
  assign n68785 = ~n70188;
  assign n68786 = ~n70179 ^ n68785;
  assign n68792 = ~n68790 | ~n74930;
  assign n68795 = ~n68792 | ~n68791;
  assign n68794 = ~n68793;
  assign n68796 = ~n68795 | ~n68794;
  assign n70182 = ~n68797 | ~n68796;
  assign n70005 = n76067 & P4_DATAO_REG_7__SCAN_IN;
  assign n70180 = ~n70005;
  assign n68800 = ~n68799;
  assign n68805 = ~n68804 | ~n68803;
  assign n68808 = ~n68807;
  assign n68811 = ~n68821;
  assign n68812 = ~n68815 ^ n68811;
  assign n68814 = ~n68812 | ~n67876;
  assign n68817 = ~n68815 ^ n68821;
  assign n68818 = ~n68817 | ~n68816;
  assign n70165 = ~n68819 | ~n68818;
  assign n70164 = n76051 & P4_DATAO_REG_8__SCAN_IN;
  assign n68820 = ~n70164;
  assign n68946 = ~n70165 ^ n68820;
  assign n68823 = ~n68822 | ~n68821;
  assign n70146 = ~n76045 & ~n76061;
  assign n68828 = ~n68826 | ~n68825;
  assign n68829 = ~n74846 | ~n59984;
  assign n68830 = ~n68829 | ~P4_DATAO_REG_18__SCAN_IN;
  assign n68833 = n70080 | n68830;
  assign n68831 = ~n63005 | ~n74315;
  assign n68832 = ~n70080 | ~n68831;
  assign n68834 = ~n68833 | ~n68832;
  assign n68835 = n70080 | n63005;
  assign n76007 = ~P4_DATAO_REG_25__SCAN_IN;
  assign n68839 = ~SEL | ~P4_DATAO_REG_24__SCAN_IN;
  assign n68840 = ~n76007 & ~n68839;
  assign n70038 = ~n68840 | ~n60715;
  assign n68842 = ~n74812 & ~n68841;
  assign n68844 = ~n68846;
  assign n68847 = ~n68846 | ~n68845;
  assign n70053 = ~n70035 | ~n68847;
  assign n70054 = ~n60178 & ~n74820;
  assign n70033 = ~n68848;
  assign n68850 = n68849 | n70033;
  assign n68853 = ~n68851 | ~n68850;
  assign n70057 = ~n68852 | ~n68853;
  assign n70060 = ~n70057 | ~n68854;
  assign n68855 = ~n68857 | ~n68856;
  assign n68861 = n68855 & n62954;
  assign n68859 = n68857 | n68856;
  assign n68860 = ~n68859 | ~n68858;
  assign n68862 = ~n68861 | ~n68860;
  assign n70059 = n68863 & n68862;
  assign n68865 = ~n70060 ^ n70059;
  assign n68864 = ~n59909 | ~P4_DATAO_REG_21__SCAN_IN;
  assign n68866 = ~n68865 | ~n68864;
  assign n68869 = ~n68867;
  assign n68870 = n68869 | n68868;
  assign n68872 = ~n74835 | ~P4_DATAO_REG_20__SCAN_IN;
  assign n70029 = ~n63005 | ~P4_DATAO_REG_19__SCAN_IN;
  assign n68874 = ~n68873;
  assign n70075 = ~n68878 | ~n68877;
  assign n70089 = ~n63296 | ~P4_DATAO_REG_17__SCAN_IN;
  assign n68879 = ~n70075 ^ n70089;
  assign n68885 = ~n68880 ^ n70087;
  assign n68883 = ~n68882 | ~n68881;
  assign n70099 = ~n63603 & ~n76012;
  assign n68887 = ~n68886;
  assign n68890 = ~n68889 | ~n68888;
  assign n68898 = ~n68893 | ~n68892;
  assign n68896 = ~n68894;
  assign n68897 = n68896 | n68895;
  assign n68900 = ~n76062 & ~n74881;
  assign n68902 = ~n68899;
  assign n68901 = ~n68900;
  assign n68903 = ~n68902 | ~n68901;
  assign n68906 = n70110 | n59930;
  assign n68905 = ~n59930 & ~n76000;
  assign n68908 = ~n68905 & ~n68904;
  assign n68907 = ~n68906 | ~n68908;
  assign n68914 = ~n70112 | ~n68907;
  assign n68909 = ~n68908;
  assign n68912 = n70110 | n68909;
  assign n68910 = ~n59930 | ~n76000;
  assign n68911 = ~n70110 | ~n68910;
  assign n68913 = ~n68912 | ~n68911;
  assign n68916 = n68915 & n59930;
  assign n68923 = ~n68919 | ~n68918;
  assign n68922 = ~n68921 | ~n68920;
  assign n70129 = ~n76054 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n70138 = ~n76037 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n68924 = ~n70129 ^ n70138;
  assign n68925 = ~n59866 | ~n68928;
  assign n68930 = ~n59866;
  assign n68929 = ~n68928;
  assign n68931 = ~n68930 | ~n68929;
  assign n68934 = ~n70011;
  assign n70010 = ~n64350 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n70013 = n63929 & P4_DATAO_REG_10__SCAN_IN;
  assign n68932 = ~n70013;
  assign n68933 = ~n70010 ^ n68932;
  assign n68943 = ~n68934 ^ n68933;
  assign n68937 = ~n68938 | ~n68935;
  assign n68942 = ~n68937 | ~n68936;
  assign n68940 = ~n68938;
  assign n68941 = ~n68940 | ~n68939;
  assign n70166 = ~n68945 ^ n68944;
  assign n70007 = ~n68946 ^ n70166;
  assign n70184 = ~n70007;
  assign n68951 = ~n68950;
  assign n68953 = ~n68952 | ~n68951;
  assign n68966 = ~n68955 ^ n70186;
  assign n68960 = n60835 | n68959;
  assign n68962 = ~n68961 | ~n68960;
  assign n68963 = ~n68962 | ~n76076;
  assign n68969 = ~n76046 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n68967 = ~n68969;
  assign n68971 = ~n68968 | ~n68967;
  assign n68977 = ~n68980 | ~n68976;
  assign n68981 = ~n74780 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n69999 = n68978 | n68981;
  assign n68987 = n68984 | n68983;
  assign n68986 = ~n68985 & ~n68994;
  assign n68991 = ~n68987 | ~n68986;
  assign n68988 = ~n76044 | ~n76055;
  assign n68990 = n68989 | n68988;
  assign n68999 = ~n68993 | ~n68992;
  assign n75004 = ~n76063;
  assign n69995 = ~n75004 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n69000 = ~n76038 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n98242 = ~P1_P1_EAX_REG_21__SCAN_IN;
  assign n69011 = ~P1_P1_EAX_REG_23__SCAN_IN | ~P1_P1_EAX_REG_22__SCAN_IN;
  assign n69012 = ~n98242 & ~n69011;
  assign n71457 = ~P1_P1_EAX_REG_24__SCAN_IN | ~n69012;
  assign n69017 = ~P1_P1_INSTQUEUE_REG_0__2__SCAN_IN | ~n97761;
  assign n69016 = ~P1_P1_INSTQUEUE_REG_4__2__SCAN_IN | ~n75033;
  assign n69021 = ~n69017 | ~n69016;
  assign n69019 = ~P1_P1_INSTQUEUE_REG_7__2__SCAN_IN | ~n97225;
  assign n69018 = ~P1_P1_INSTQUEUE_REG_9__2__SCAN_IN | ~n97979;
  assign n69020 = ~n69019 | ~n69018;
  assign n69029 = ~n69021 & ~n69020;
  assign n69023 = ~P1_P1_INSTQUEUE_REG_13__2__SCAN_IN | ~n97754;
  assign n69022 = ~P1_P1_INSTQUEUE_REG_3__2__SCAN_IN | ~n97895;
  assign n69027 = ~n69023 | ~n69022;
  assign n69025 = ~P1_P1_INSTQUEUE_REG_10__2__SCAN_IN | ~n97747;
  assign n69024 = ~P1_P1_INSTQUEUE_REG_2__2__SCAN_IN | ~n97746;
  assign n69026 = ~n69025 | ~n69024;
  assign n69028 = ~n69027 & ~n69026;
  assign n69045 = ~n69029 | ~n69028;
  assign n69031 = ~P1_P1_INSTQUEUE_REG_14__2__SCAN_IN | ~n75052;
  assign n69030 = ~P1_P1_INSTQUEUE_REG_11__2__SCAN_IN | ~n97185;
  assign n69035 = ~n69031 | ~n69030;
  assign n69033 = ~P1_P1_INSTQUEUE_REG_8__2__SCAN_IN | ~n59935;
  assign n69032 = ~P1_P1_INSTQUEUE_REG_15__2__SCAN_IN | ~n97743;
  assign n69034 = ~n69033 | ~n69032;
  assign n69043 = ~n69035 & ~n69034;
  assign n69037 = ~P1_P1_INSTQUEUE_REG_12__2__SCAN_IN | ~n97203;
  assign n69036 = ~P1_P1_INSTQUEUE_REG_1__2__SCAN_IN | ~n75055;
  assign n69041 = ~n69037 | ~n69036;
  assign n69039 = ~P1_P1_INSTQUEUE_REG_6__2__SCAN_IN | ~n59938;
  assign n69038 = ~P1_P1_INSTQUEUE_REG_5__2__SCAN_IN | ~n97303;
  assign n69040 = ~n69039 | ~n69038;
  assign n69042 = ~n69041 & ~n69040;
  assign n69044 = ~n69043 | ~n69042;
  assign n70205 = ~n69045 & ~n69044;
  assign n70204 = ~n69047 | ~n69046;
  assign n74457 = n76028 & DIN_26_;
  assign n71177 = ~n74457 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n71671 = ~n76038 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n71368 = ~n70003 | ~n70002;
  assign n71385 = ~n71659 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n71373 = n76046 & P4_DATAO_REG_5__SCAN_IN;
  assign n71382 = ~n71373;
  assign n70004 = ~n71385 ^ n71382;
  assign n70006 = n70007 | n70182;
  assign n70009 = ~n70006 | ~n70005;
  assign n70008 = ~n70007 | ~n70182;
  assign n70175 = n70009 & n70008;
  assign n70021 = n70011 | n70010;
  assign n70012 = ~n70011 | ~n70010;
  assign n70015 = ~n70021 | ~n70012;
  assign n70014 = ~n70015 | ~n70016;
  assign n70019 = ~n70014 | ~n70013;
  assign n70017 = ~n70016;
  assign n70018 = ~n59865 | ~n70017;
  assign n71227 = ~n70021 | ~n70020;
  assign n70024 = ~n70022;
  assign n70025 = ~n70024 | ~n70023;
  assign n71232 = ~n59930 | ~P4_DATAO_REG_15__SCAN_IN;
  assign n71329 = ~n76054 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n70026 = ~n71232 ^ n71329;
  assign n70106 = ~n71234 ^ n70026;
  assign n70027 = ~n70075;
  assign n70031 = ~n70028;
  assign n70030 = ~n70029;
  assign n70032 = ~n70031 | ~n70030;
  assign n71303 = ~n71293 & ~n60217;
  assign n70073 = ~n71295 ^ n71303;
  assign n70034 = ~n70033 | ~n70038;
  assign n71243 = ~n70035 | ~n70034;
  assign n70036 = ~n70038;
  assign n71258 = ~n70036 | ~n59870;
  assign n70037 = ~n59870 | ~P4_DATAO_REG_24__SCAN_IN;
  assign n70039 = ~n70038 | ~n70037;
  assign n70046 = n71258 & n70039;
  assign n70040 = ~n76007 | ~n74277;
  assign n70045 = ~n59991 | ~n70040;
  assign n75999 = ~P4_DATAO_REG_26__SCAN_IN;
  assign n70041 = ~SEL | ~P4_DATAO_REG_25__SCAN_IN;
  assign n70042 = ~n75999 & ~n70041;
  assign n71517 = ~n70042 | ~n60715;
  assign n70044 = ~n70043 | ~n75999;
  assign n71259 = ~n70046 | ~n70047;
  assign n70048 = ~n70046;
  assign n71242 = ~n71259 | ~n70049;
  assign n70051 = ~n71243 ^ n71242;
  assign n70050 = ~n75996 & ~n64572;
  assign n71246 = ~n70051 | ~n70050;
  assign n70055 = ~n70053;
  assign n70056 = ~n70055 | ~n70054;
  assign n70058 = ~n60178 & ~n59912;
  assign n71275 = ~n71279 & ~n63855;
  assign n70061 = n70060 | n70059;
  assign n70065 = ~n70062 | ~n70061;
  assign n71278 = ~n70066 | ~n70065;
  assign n71283 = ~n70067 | ~n71278;
  assign n70070 = n70069 | n70068;
  assign n71284 = ~n70071 | ~n70070;
  assign n70072 = ~n74882 & ~n74846;
  assign n71239 = ~n74315 | ~P4_DATAO_REG_19__SCAN_IN;
  assign n70085 = ~n70073 ^ n71294;
  assign n70076 = ~n70074;
  assign n70078 = n70076 | n70075;
  assign n70086 = n70078 & n70077;
  assign n70079 = ~n70087;
  assign n70092 = ~n70086 | ~n70079;
  assign n70081 = n59955 | n61395;
  assign n70083 = ~n70082 | ~n70081;
  assign n70084 = ~n70083 | ~n74315;
  assign n71300 = ~n70092 | ~n70084;
  assign n71308 = ~n70085 ^ n71300;
  assign n70088 = ~n70086;
  assign n70091 = ~n70088 | ~n70087;
  assign n70090 = ~n70089;
  assign n70093 = n70091 & n70090;
  assign n70094 = ~n70093 | ~n70092;
  assign n71307 = ~n70095 | ~n70094;
  assign n70100 = ~n70098;
  assign n70101 = ~n70100 | ~n70099;
  assign n70104 = ~n71315 ^ n71313;
  assign n70103 = ~n76000 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n70109 = n70108 | n59861;
  assign n70116 = n70109 & n59930;
  assign n70111 = ~n70110;
  assign n70114 = n70112 | n70111;
  assign n70115 = ~n70114 | ~n70113;
  assign n70117 = ~n70116 | ~n70115;
  assign n70120 = ~n70118 | ~n70117;
  assign n71335 = ~n70119 | ~n70120;
  assign n70121 = ~n70120;
  assign n70123 = ~n70122 | ~n70121;
  assign n71223 = ~n63929 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n70127 = ~n71349 ^ n71223;
  assign n70132 = n70128 | n70129;
  assign n71352 = ~n64350 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n71341 = ~n76037 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n70126 = ~n71352 ^ n71341;
  assign n71216 = ~n71343 ^ n70126;
  assign n70131 = ~n70128;
  assign n70130 = ~n70129;
  assign n70133 = n70131 | n70130;
  assign n70134 = n70132 & n70133;
  assign n70142 = ~n70134 | ~n70135;
  assign n70137 = ~n70134;
  assign n70136 = ~n70135;
  assign n70140 = ~n70137 | ~n70136;
  assign n70139 = ~n70138;
  assign n70141 = ~n70140 | ~n70139;
  assign n71219 = ~n70142 | ~n70141;
  assign n70155 = ~n70145 ^ n71210;
  assign n70153 = ~n70155;
  assign n70147 = n70149 | n70148;
  assign n70151 = ~n70147 | ~n70146;
  assign n70150 = ~n70149 | ~n70148;
  assign n70154 = ~n70151 | ~n70150;
  assign n70152 = ~n70154;
  assign n71206 = ~n70155 | ~n70154;
  assign n70156 = ~n71205 | ~n71206;
  assign n70157 = ~n70165 | ~n76051;
  assign n70161 = n76067 & P4_DATAO_REG_8__SCAN_IN;
  assign n70159 = ~n70158 | ~n70161;
  assign n70163 = ~n70165 | ~n70164;
  assign n70162 = ~n70161;
  assign n70168 = n70165 | n70164;
  assign n70167 = ~n70166;
  assign n70169 = ~n70168 | ~n70167;
  assign n70171 = ~n70170 | ~n70169;
  assign n70172 = ~n70174;
  assign n71196 = ~n70173 | ~n70172;
  assign n71194 = ~n70175 | ~n70174;
  assign n71191 = ~n71194 | ~n71196;
  assign n71193 = ~n76043 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n71369 = ~n71191 ^ n70176;
  assign n70177 = ~n71369;
  assign n70181 = ~n70180 ^ n70179;
  assign n70183 = ~n70182 ^ n70181;
  assign n70185 = ~n70184 ^ n70183;
  assign n70189 = ~n71371;
  assign n71377 = ~n61519 | ~n70187;
  assign n71383 = ~n71374;
  assign n70194 = ~n70196;
  assign n71189 = ~n70196 | ~n70195;
  assign n71406 = ~n75004 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n70197 = ~n71404 ^ n71406;
  assign n71455 = ~n70205 & ~n70204;
  assign n70207 = ~P1_P1_INSTQUEUE_REG_0__3__SCAN_IN | ~n97761;
  assign n70206 = ~P1_P1_INSTQUEUE_REG_6__3__SCAN_IN | ~n59938;
  assign n70211 = ~n70207 | ~n70206;
  assign n70209 = ~P1_P1_INSTQUEUE_REG_3__3__SCAN_IN | ~n97895;
  assign n70208 = ~P1_P1_INSTQUEUE_REG_1__3__SCAN_IN | ~n75055;
  assign n70210 = ~n70209 | ~n70208;
  assign n70235 = ~n70211 & ~n70210;
  assign n70213 = ~P1_P1_INSTQUEUE_REG_13__3__SCAN_IN | ~n97754;
  assign n70212 = ~P1_P1_INSTQUEUE_REG_2__3__SCAN_IN | ~n59936;
  assign n70215 = ~n70213 | ~n70212;
  assign n70214 = n97999 & P1_P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n70217 = ~n70215 & ~n70214;
  assign n70216 = ~n97747 | ~P1_P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n70233 = ~n70217 | ~n70216;
  assign n70219 = ~P1_P1_INSTQUEUE_REG_9__3__SCAN_IN | ~n97979;
  assign n70218 = ~P1_P1_INSTQUEUE_REG_4__3__SCAN_IN | ~n75033;
  assign n70223 = ~n70219 | ~n70218;
  assign n70221 = ~P1_P1_INSTQUEUE_REG_12__3__SCAN_IN | ~n97203;
  assign n70220 = ~P1_P1_INSTQUEUE_REG_11__3__SCAN_IN | ~n97185;
  assign n70222 = ~n70221 | ~n70220;
  assign n70231 = ~n70223 & ~n70222;
  assign n70225 = ~P1_P1_INSTQUEUE_REG_15__3__SCAN_IN | ~n97743;
  assign n70224 = ~P1_P1_INSTQUEUE_REG_14__3__SCAN_IN | ~n75052;
  assign n70229 = ~n70225 | ~n70224;
  assign n70227 = ~P1_P1_INSTQUEUE_REG_8__3__SCAN_IN | ~n59935;
  assign n70226 = ~P1_P1_INSTQUEUE_REG_7__3__SCAN_IN | ~n97225;
  assign n70228 = ~n70227 | ~n70226;
  assign n70230 = ~n70229 & ~n70228;
  assign n70232 = ~n70231 | ~n70230;
  assign n70234 = ~n70233 & ~n70232;
  assign n71454 = ~n70235 | ~n70234;
  assign n71456 = ~P1_P1_EAX_REG_26__SCAN_IN | ~P1_P1_EAX_REG_25__SCAN_IN;
  assign n74458 = n76028 & DIN_27_;
  assign n74762 = ~n74458;
  assign n71688 = ~n71171 & ~n74762;
  assign n71173 = ~n71172 | ~n71177;
  assign n71184 = ~n71174 | ~n71173;
  assign n71178 = ~n71177;
  assign n71179 = ~n71178 | ~n76038;
  assign n76082 = ~n74457;
  assign n74204 = ~n71188 & ~n76082;
  assign n71673 = ~n74204;
  assign n71195 = ~n71194 | ~n59969;
  assign n71654 = ~n76076 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n74238 = ~n76046 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n71201 = n76043 & P4_DATAO_REG_8__SCAN_IN;
  assign n71204 = ~n71203;
  assign n71207 = ~n71205 | ~n71204;
  assign n71640 = ~n71207 | ~n71206;
  assign n71639 = n76067 & P4_DATAO_REG_9__SCAN_IN;
  assign n71638 = ~n71640 ^ n71639;
  assign n71209 = ~n59859;
  assign n71208 = ~n71212;
  assign n71211 = ~n71209 | ~n71208;
  assign n71215 = ~n71211 | ~n71210;
  assign n71214 = ~n59860 | ~n71212;
  assign n71488 = ~n71215 | ~n71214;
  assign n71489 = ~n76051 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n71362 = ~n71488 ^ n71489;
  assign n71217 = ~n71216;
  assign n71218 = ~n71221;
  assign n71222 = n71218 | n71219;
  assign n71220 = ~n71219;
  assign n71225 = ~n71222 | ~n71358;
  assign n71226 = ~n71223;
  assign n71224 = ~n71227 | ~n71226;
  assign n71229 = ~n71225 | ~n71224;
  assign n71228 = n71227 | n71226;
  assign n71497 = ~n71230 & ~n76061;
  assign n71326 = ~n71234 ^ n71232;
  assign n71231 = ~n71327;
  assign n71332 = ~n71326 | ~n71231;
  assign n71233 = ~n71232;
  assign n71235 = ~n71234 | ~n71233;
  assign n71606 = ~n71332 | ~n71235;
  assign n71605 = ~n76062 & ~n74360;
  assign n71324 = ~n71606 ^ n71605;
  assign n71236 = n71315 | n71313;
  assign n71596 = ~n71237 | ~n71236;
  assign n71238 = ~n71295;
  assign n71241 = n71240 | n71239;
  assign n71244 = ~n71242;
  assign n71245 = ~n71244 | ~n71243;
  assign n71513 = ~n71246 | ~n71245;
  assign n71247 = ~SEL | ~P4_DATAO_REG_26__SCAN_IN;
  assign n71249 = ~n75994 & ~n71247;
  assign n71527 = ~n71249 | ~n60715;
  assign n71254 = ~n71527 ^ n71517;
  assign n71250 = n75999 & n59915;
  assign n71253 = ~n74812 & ~n71250;
  assign n71252 = ~n71251 | ~n75994;
  assign n71255 = ~n59870 | ~P4_DATAO_REG_25__SCAN_IN;
  assign n71257 = ~n71256 | ~n71255;
  assign n71534 = ~n71259 | ~n71258;
  assign n71261 = ~n71533 ^ n71534;
  assign n71260 = ~n76032 & ~n64572;
  assign n71537 = ~n71261 | ~n71260;
  assign n71262 = n71261 | n71260;
  assign n71263 = ~n75996 & ~n59912;
  assign n71508 = ~n60178 & ~n63855;
  assign n71266 = ~n71264;
  assign n71267 = ~n71266 | ~n71265;
  assign n71270 = ~n71268 | ~n71267;
  assign n71511 = ~n71269 | ~n71270;
  assign n71272 = ~n71269;
  assign n71271 = ~n71270;
  assign n71273 = ~n71272 | ~n71271;
  assign n71502 = ~n71511 | ~n71273;
  assign n71276 = ~n71274;
  assign n71277 = ~n71276 | ~n71275;
  assign n71503 = ~n71278 | ~n71277;
  assign n71281 = ~n71502 ^ n71503;
  assign n71280 = ~n71279 & ~n74846;
  assign n71548 = ~n74882 & ~n59984;
  assign n71564 = ~n63296 | ~P4_DATAO_REG_19__SCAN_IN;
  assign n71282 = ~n71548 ^ n71564;
  assign n71285 = ~n71283;
  assign n71286 = ~n71285 | ~n71284;
  assign n71549 = ~n71287 | ~n71286;
  assign n71292 = ~n71289 | ~n71288;
  assign n71291 = ~n71288;
  assign n71290 = ~n71289;
  assign n71571 = ~n71291 | ~n71290;
  assign n71580 = ~n71293 & ~n76012;
  assign n71296 = ~n71294;
  assign n71297 = n71296 | n71295;
  assign n71299 = n71298 & n71297;
  assign n71306 = ~n71299 | ~n71300;
  assign n71302 = ~n71299;
  assign n71301 = ~n71300;
  assign n71304 = ~n71302 | ~n71301;
  assign n71305 = ~n71304 | ~n71303;
  assign n71578 = ~n71306 | ~n71305;
  assign n71590 = ~n76000 | ~P4_DATAO_REG_17__SCAN_IN;
  assign n71309 = ~n71308 | ~n71307;
  assign n71587 = ~n71310 | ~n71309;
  assign n71312 = ~n71597 ^ n71596;
  assign n71311 = ~n59930 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n71322 = ~n71312 | ~n71311;
  assign n71316 = ~n71313;
  assign n71314 = ~n71316 & ~DIN_10_;
  assign n71318 = n71315 | n71314;
  assign n71317 = ~n71316 | ~DIN_10_;
  assign n71319 = ~n71318 | ~n71317;
  assign n71321 = ~n71597 ^ n71319;
  assign n71320 = ~DIN_11_ | ~P4_DATAO_REG_16__SCAN_IN;
  assign n71598 = n71321 | n71320;
  assign n71323 = ~n71322 | ~n71598;
  assign n71337 = n71325 & n71608;
  assign n71328 = ~n71326;
  assign n71331 = ~n71328 | ~n71327;
  assign n71330 = ~n71329;
  assign n71333 = n71331 & n71330;
  assign n71334 = ~n71333 | ~n71332;
  assign n71612 = ~n71335 | ~n71334;
  assign n71610 = ~n76037 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n71336 = ~n71612 ^ n71610;
  assign n71614 = ~n71337 | ~n71336;
  assign n71339 = ~n71336;
  assign n71338 = ~n71337;
  assign n71340 = ~n71339 | ~n71338;
  assign n71342 = ~n71341;
  assign n71348 = ~n71343 ^ n71342;
  assign n71355 = n71348 | n71349;
  assign n71344 = ~n71343 | ~n71342;
  assign n71620 = ~n71355 | ~n71344;
  assign n71618 = ~n64350 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n71626 = ~n63929 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n71346 = ~n71618 ^ n71626;
  assign n71347 = ~n71620 ^ n71346;
  assign n71360 = ~n71619 ^ n71347;
  assign n71351 = ~n71348;
  assign n71350 = ~n71349;
  assign n71354 = n71351 | n71350;
  assign n71353 = ~n71352;
  assign n71356 = n71354 & n71353;
  assign n71357 = ~n71356 | ~n71355;
  assign n71359 = ~n71358 | ~n71357;
  assign n71636 = ~n71362 ^ n71492;
  assign n71653 = ~n71363 ^ n71646;
  assign n71367 = ~n71365 ^ n71657;
  assign n71366 = ~n76081 & ~n76044;
  assign n71665 = n71367 | n71366;
  assign n71666 = ~n71367 | ~n71366;
  assign n71482 = ~n71665 | ~n71666;
  assign n71370 = ~n76076 & ~n76046;
  assign n71376 = ~n71372 | ~n60776;
  assign n71375 = ~n71374 | ~n71373;
  assign n71380 = ~n71376 | ~n71375;
  assign n71378 = ~n71377;
  assign n71379 = ~n71378 | ~n71382;
  assign n71386 = ~n71384 ^ n71383;
  assign n71485 = ~n71390 | ~n71389;
  assign n71393 = ~n75004 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n71476 = ~n71393;
  assign n71395 = ~n71392 | ~n71476;
  assign n71399 = ~n71401;
  assign n71396 = ~n76038;
  assign n71400 = ~n71397 & ~n71396;
  assign n71470 = ~n71399 | ~n71398;
  assign n71471 = ~n71401 | ~n71400;
  assign n71411 = ~n71470 | ~n71471;
  assign n71408 = ~n71405 ^ n71404;
  assign n71407 = ~n71406;
  assign n71409 = ~n71408 | ~n71407;
  assign n74212 = ~n71411 ^ n71469;
  assign n71425 = ~P1_P1_INSTQUEUE_REG_8__4__SCAN_IN | ~n59935;
  assign n71424 = ~P1_P1_INSTQUEUE_REG_5__4__SCAN_IN | ~n97303;
  assign n71429 = ~n71425 | ~n71424;
  assign n71427 = ~P1_P1_INSTQUEUE_REG_15__4__SCAN_IN | ~n97743;
  assign n71426 = ~P1_P1_INSTQUEUE_REG_6__4__SCAN_IN | ~n59938;
  assign n71428 = ~n71427 | ~n71426;
  assign n71437 = ~n71429 & ~n71428;
  assign n71431 = ~P1_P1_INSTQUEUE_REG_7__4__SCAN_IN | ~n97225;
  assign n71430 = ~P1_P1_INSTQUEUE_REG_9__4__SCAN_IN | ~n98034;
  assign n71435 = ~n71431 | ~n71430;
  assign n71433 = ~P1_P1_INSTQUEUE_REG_10__4__SCAN_IN | ~n97747;
  assign n71432 = ~P1_P1_INSTQUEUE_REG_2__4__SCAN_IN | ~n97746;
  assign n71434 = ~n71433 | ~n71432;
  assign n71436 = ~n71435 & ~n71434;
  assign n71453 = ~n71437 | ~n71436;
  assign n71439 = ~P1_P1_INSTQUEUE_REG_14__4__SCAN_IN | ~n75052;
  assign n71438 = ~P1_P1_INSTQUEUE_REG_1__4__SCAN_IN | ~n75055;
  assign n71443 = ~n71439 | ~n71438;
  assign n71441 = ~P1_P1_INSTQUEUE_REG_12__4__SCAN_IN | ~n97203;
  assign n71440 = ~P1_P1_INSTQUEUE_REG_3__4__SCAN_IN | ~n97895;
  assign n71442 = ~n71441 | ~n71440;
  assign n71451 = ~n71443 & ~n71442;
  assign n71445 = ~P1_P1_INSTQUEUE_REG_11__4__SCAN_IN | ~n97185;
  assign n71444 = ~P1_P1_INSTQUEUE_REG_4__4__SCAN_IN | ~n75033;
  assign n71449 = ~n71445 | ~n71444;
  assign n71447 = ~P1_P1_INSTQUEUE_REG_13__4__SCAN_IN | ~n97754;
  assign n71446 = ~P1_P1_INSTQUEUE_REG_0__4__SCAN_IN | ~n97761;
  assign n71448 = ~n71447 | ~n71446;
  assign n71450 = ~n71449 & ~n71448;
  assign n71452 = ~n71451 | ~n71450;
  assign n71705 = ~n71453 & ~n71452;
  assign n71704 = ~n71455 | ~n71454;
  assign n71741 = ~n71457 & ~n71456;
  assign n71472 = ~n71470 | ~n71469;
  assign n74460 = ~n71472 | ~n71471;
  assign n71475 = ~n59942 & ~n71476;
  assign n71477 = ~n59942 | ~n71476;
  assign n74451 = ~n76038 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n71480 = ~n71479 | ~n71478;
  assign n71484 = ~n71482 ^ n71664;
  assign n71486 = n71484 | n71483;
  assign n71493 = ~n71488;
  assign n71491 = ~n71492 | ~n71493;
  assign n71490 = ~n71489;
  assign n71495 = ~n71491 | ~n71490;
  assign n71494 = n71493 | n71492;
  assign n71498 = ~n71496;
  assign n71499 = ~n71498 | ~n71497;
  assign n74400 = ~n76051 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n74962 = ~n76067 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n71504 = ~n71502;
  assign n71505 = ~n71504 | ~n71503;
  assign n71509 = ~n71507;
  assign n71510 = ~n71509 | ~n71508;
  assign n74319 = ~n71511 | ~n71510;
  assign n71514 = ~n71512;
  assign n71515 = ~n71514 | ~n71513;
  assign n74309 = ~n71516 | ~n71515;
  assign n74307 = ~n74835 | ~P4_DATAO_REG_23__SCAN_IN;
  assign n74317 = ~n74309 ^ n74307;
  assign n71518 = ~n71517;
  assign n71519 = ~n71518 | ~n71527;
  assign n74291 = ~n71520 | ~n71519;
  assign n74290 = ~n76007 & ~n64572;
  assign n71531 = ~n74291 ^ n74290;
  assign n71522 = ~n71521 | ~P4_DATAO_REG_27__SCAN_IN;
  assign n74279 = ~P4_DATAO_REG_28__SCAN_IN;
  assign n71523 = ~n71522 | ~n74279;
  assign n74270 = n71524 | n74822;
  assign n74271 = ~n75999 & ~n63724;
  assign n71525 = ~n71527;
  assign n74274 = ~n71526 | ~n71525;
  assign n71528 = ~n71526;
  assign n71529 = ~n71528 | ~n71527;
  assign n71530 = ~n74274 | ~n71529;
  assign n71532 = ~n71531 | ~n71530;
  assign n74296 = ~n76032 & ~n59911;
  assign n71538 = ~n74295 ^ n74296;
  assign n71535 = ~n71533;
  assign n71536 = ~n71535 | ~n71534;
  assign n71539 = ~n71537 | ~n71536;
  assign n74299 = ~n71538 | ~n71539;
  assign n71541 = ~n71538;
  assign n71540 = ~n71539;
  assign n71542 = ~n71541 | ~n71540;
  assign n74316 = ~n74299 | ~n71542;
  assign n74322 = ~n63005 | ~P4_DATAO_REG_22__SCAN_IN;
  assign n71543 = ~n74316 ^ n74322;
  assign n71544 = ~n74317 ^ n71543;
  assign n74329 = ~n74315 | ~P4_DATAO_REG_21__SCAN_IN;
  assign n71551 = ~n63296 | ~P4_DATAO_REG_20__SCAN_IN;
  assign n71558 = ~n74336 ^ n71551;
  assign n71560 = ~n71549 ^ n71548;
  assign n71567 = n71560 | n71561;
  assign n71556 = n71558 | n71567;
  assign n71557 = ~n71549 | ~n71548;
  assign n74337 = ~n71551;
  assign n71550 = ~n71557 & ~n74337;
  assign n71554 = n74336 | n71550;
  assign n71552 = n71557 | n71551;
  assign n71553 = ~n74336 | ~n71552;
  assign n71555 = ~n71554 | ~n71553;
  assign n74335 = n71567 & n71557;
  assign n71563 = ~n71560;
  assign n71562 = ~n71561;
  assign n71566 = n71563 | n71562;
  assign n71565 = ~n71564;
  assign n71569 = ~n71566 | ~n71565;
  assign n71568 = ~n71567;
  assign n71570 = n71569 | n71568;
  assign n74349 = ~n71571 | ~n71570;
  assign n71573 = ~n74353 & ~n76012;
  assign n74352 = ~n71572 | ~n71573;
  assign n71574 = ~n71573;
  assign n71576 = ~n71575 | ~n71574;
  assign n74267 = ~n74352 | ~n71576;
  assign n71579 = ~n71577;
  assign n71583 = n71579 | n71578;
  assign n71581 = ~n71580;
  assign n74266 = ~n71583 | ~n71582;
  assign n71585 = ~n74267 ^ n74266;
  assign n71584 = ~n76000 | ~P4_DATAO_REG_18__SCAN_IN;
  assign n71586 = ~n71585 | ~n71584;
  assign n71594 = n71588 | n71587;
  assign n71592 = ~n71589;
  assign n71591 = ~n71590;
  assign n71593 = n71592 | n71591;
  assign n74262 = ~n71594 | ~n71593;
  assign n71595 = ~n59930 | ~P4_DATAO_REG_17__SCAN_IN;
  assign n71599 = ~n71597 | ~n71596;
  assign n74364 = ~n71599 | ~n71598;
  assign n74362 = ~n76054 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n71601 = ~n74364 ^ n74362;
  assign n74366 = ~n71600 | ~n71601;
  assign n71602 = ~n71601;
  assign n71604 = ~n71603 | ~n71602;
  assign n74373 = ~n74366 | ~n71604;
  assign n71607 = ~n71606 | ~n71605;
  assign n74374 = ~n71608 | ~n71607;
  assign n71609 = ~n76062 & ~n74367;
  assign n71611 = ~n71610;
  assign n71613 = ~n71612 | ~n71611;
  assign n74378 = ~n71614 | ~n71613;
  assign n74377 = n64350 & P4_DATAO_REG_14__SCAN_IN;
  assign n71615 = ~n74378 ^ n74377;
  assign n71617 = ~n71616 | ~n71615;
  assign n74393 = ~n74380 | ~n71617;
  assign n71625 = ~n71619 ^ n71620;
  assign n71624 = ~n71618;
  assign n71629 = ~n71625 | ~n71624;
  assign n71621 = ~n71619;
  assign n71622 = ~n71621 | ~n71620;
  assign n71623 = n63929 & P4_DATAO_REG_13__SCAN_IN;
  assign n71628 = n71625 | n71624;
  assign n71627 = ~n71626;
  assign n71630 = n71628 & n71627;
  assign n71631 = ~n71630 | ~n71629;
  assign n74256 = n60778 & n71631;
  assign n71632 = ~n74930 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n71634 = ~n71633 | ~n71632;
  assign n71637 = ~n71636;
  assign n71642 = n71638 | n71637;
  assign n71641 = ~n71640 | ~n71639;
  assign n71644 = ~n71642 | ~n71641;
  assign n71643 = n76043 & P4_DATAO_REG_9__SCAN_IN;
  assign n71645 = n71644 | n71643;
  assign n74440 = ~n71644 | ~n71643;
  assign n74432 = ~n76076 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n71649 = ~n71654;
  assign n71651 = ~n71653 | ~n71648;
  assign n74247 = ~n76046 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n71652 = ~n74250 ^ n74247;
  assign n71656 = ~n71653;
  assign n74232 = ~n71658 | ~n71657;
  assign n71661 = ~n71659 & ~n76046;
  assign n71662 = ~n71661 & ~n71660;
  assign n71663 = ~n74232 | ~n71662;
  assign n75008 = ~n74780 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n71667 = ~n75006 ^ n75008;
  assign n74454 = ~n71668 ^ n74446;
  assign n74462 = ~n71669 ^ n74454;
  assign n71670 = ~n74462 ^ n74460;
  assign n74463 = ~n74457 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n74203 = n71670 | n74463;
  assign n71674 = n71672 | n71671;
  assign n71677 = ~n71676 | ~n71675;
  assign n71679 = ~n71678 | ~n71677;
  assign n71680 = ~n74212 | ~n71679;
  assign n74211 = n71681 & n71680;
  assign n74207 = ~n74458 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n71682 = ~n74207;
  assign n71687 = ~n71694 | ~n71688;
  assign n74728 = ~n76028 | ~P4_DATAO_REG_0__SCAN_IN;
  assign n71685 = ~n74728;
  assign n71686 = ~n71685 | ~DIN_28_;
  assign n71689 = n71694 | n71688;
  assign n71690 = ~n71689 | ~n71693;
  assign n74756 = n76028 & DIN_28_;
  assign n71695 = n71693 & n74458;
  assign n74475 = ~n71705 & ~n71704;
  assign n71707 = ~P1_P1_INSTQUEUE_REG_8__5__SCAN_IN | ~n59935;
  assign n71706 = ~P1_P1_INSTQUEUE_REG_13__5__SCAN_IN | ~n97754;
  assign n71711 = ~n71707 | ~n71706;
  assign n71709 = ~P1_P1_INSTQUEUE_REG_7__5__SCAN_IN | ~n97225;
  assign n71708 = ~P1_P1_INSTQUEUE_REG_5__5__SCAN_IN | ~n97303;
  assign n71710 = ~n71709 | ~n71708;
  assign n71735 = ~n71711 & ~n71710;
  assign n71715 = n75055 & P1_P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n71713 = ~P1_P1_INSTQUEUE_REG_3__5__SCAN_IN | ~n97895;
  assign n71712 = ~P1_P1_INSTQUEUE_REG_14__5__SCAN_IN | ~n75052;
  assign n71714 = ~n71713 | ~n71712;
  assign n71717 = ~n71715 & ~n71714;
  assign n71716 = ~n59938 | ~P1_P1_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n71733 = ~n71717 | ~n71716;
  assign n71719 = ~P1_P1_INSTQUEUE_REG_15__5__SCAN_IN | ~n97743;
  assign n71718 = ~P1_P1_INSTQUEUE_REG_9__5__SCAN_IN | ~n98034;
  assign n71723 = ~n71719 | ~n71718;
  assign n71721 = ~P1_P1_INSTQUEUE_REG_0__5__SCAN_IN | ~n97761;
  assign n71720 = ~P1_P1_INSTQUEUE_REG_11__5__SCAN_IN | ~n97185;
  assign n71722 = ~n71721 | ~n71720;
  assign n71731 = ~n71723 & ~n71722;
  assign n71725 = ~P1_P1_INSTQUEUE_REG_10__5__SCAN_IN | ~n98037;
  assign n71724 = ~P1_P1_INSTQUEUE_REG_12__5__SCAN_IN | ~n97203;
  assign n71729 = ~n71725 | ~n71724;
  assign n71727 = ~P1_P1_INSTQUEUE_REG_2__5__SCAN_IN | ~n59936;
  assign n71726 = ~P1_P1_INSTQUEUE_REG_4__5__SCAN_IN | ~n75033;
  assign n71728 = ~n71727 | ~n71726;
  assign n71730 = ~n71729 & ~n71728;
  assign n71732 = ~n71731 | ~n71730;
  assign n71734 = ~n71733 & ~n71732;
  assign n74474 = ~n71735 | ~n71734;
  assign n71744 = ~n71742 | ~n71741;
  assign n71743 = ~P1_P1_EAX_REG_28__SCAN_IN | ~P1_P1_EAX_REG_27__SCAN_IN;
  assign n74508 = ~n71744 & ~n71743;
  assign n75028 = n74508 & n97930;
  assign n74205 = ~n74212 | ~n74204;
  assign n74732 = ~n74756 | ~P4_DATAO_REG_1__SCAN_IN;
  assign n74218 = ~n74209 | ~n74737;
  assign n74214 = ~n74212;
  assign n74213 = n74762 & n76082;
  assign n74215 = n74219 & n74732;
  assign n74737 = ~n74732;
  assign n74223 = ~n76055 | ~n76063;
  assign n74224 = ~n74780 | ~n75004;
  assign n74225 = ~n75006 | ~n74224;
  assign n74237 = ~n74232 | ~n60808;
  assign n74227 = ~n74247;
  assign n74230 = ~n74237 | ~n74227;
  assign n74228 = ~n74238 & ~n76064;
  assign n74229 = ~n74240 | ~n74228;
  assign n74231 = ~n74230 | ~n74229;
  assign n74235 = n74232 | n60808;
  assign n74233 = ~n74238 & ~n76044;
  assign n74234 = ~n74240 | ~n74233;
  assign n74236 = n74235 & n74234;
  assign n74244 = ~n74248;
  assign n74242 = ~n74237 | ~n74247;
  assign n74239 = ~n74238 & ~P4_DATAO_REG_7__SCAN_IN;
  assign n74241 = ~n74240 | ~n74239;
  assign n74243 = ~n74242 | ~n74241;
  assign n74783 = ~n74780 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n74252 = ~n74249;
  assign n74251 = ~n74250;
  assign n74776 = ~n74254 | ~n74253;
  assign n74766 = ~n76038 | ~P4_DATAO_REG_4__SCAN_IN;
  assign n74444 = ~n74776 ^ n74766;
  assign n74258 = ~n74255;
  assign n74257 = ~n74256;
  assign n74259 = ~n74258 | ~n74257;
  assign n74937 = ~n76051 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n74950 = ~n76067 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n74263 = ~n74261;
  assign n74264 = ~n74263 | ~n61004;
  assign n74268 = n74267 | n74266;
  assign n74897 = ~n74269 | ~n74268;
  assign n74896 = n59930 & P4_DATAO_REG_18__SCAN_IN;
  assign n74358 = ~n74897 ^ n74896;
  assign n74272 = ~n74270;
  assign n74273 = ~n74272 | ~n74271;
  assign n74800 = ~n74274 | ~n74273;
  assign n74275 = P4_DATAO_REG_28__SCAN_IN & P4_DATAO_REG_29__SCAN_IN;
  assign n74821 = ~n62948 | ~n74275;
  assign n74278 = ~n74279 | ~n74277;
  assign n74282 = ~n59991 | ~n74278;
  assign n74280 = ~n74279 & ~n63317;
  assign n74281 = ~n74280 & ~P4_DATAO_REG_29__SCAN_IN;
  assign n74283 = ~n74282 & ~n74281;
  assign n74286 = ~n74284 | ~n74283;
  assign n74285 = ~n59870 | ~P4_DATAO_REG_27__SCAN_IN;
  assign n74287 = ~n74286 | ~n74285;
  assign n74289 = ~n62954 | ~P4_DATAO_REG_26__SCAN_IN;
  assign n74802 = n74288 | n74289;
  assign n74292 = ~n74291 | ~n74290;
  assign n74293 = ~n74831 ^ n74832;
  assign n74294 = ~n59907 | ~P4_DATAO_REG_25__SCAN_IN;
  assign n74842 = ~n76032 & ~n63855;
  assign n74297 = ~n74295;
  assign n74298 = ~n74297 | ~n74296;
  assign n74301 = ~n74299 | ~n74298;
  assign n74845 = ~n74300 | ~n74301;
  assign n74303 = ~n74300;
  assign n74302 = ~n74301;
  assign n74304 = ~n74303 | ~n74302;
  assign n74856 = ~n74845 | ~n74304;
  assign n74306 = ~n74317;
  assign n74305 = ~n74316;
  assign n74311 = n74306 | n74305;
  assign n74308 = ~n74307;
  assign n74310 = n74309 | n74308;
  assign n74855 = ~n74311 | ~n74310;
  assign n74312 = ~n74856 ^ n74855;
  assign n74313 = ~n63005 | ~P4_DATAO_REG_23__SCAN_IN;
  assign n74858 = n74312 | n74313;
  assign n74862 = ~n74315 | ~P4_DATAO_REG_22__SCAN_IN;
  assign n74321 = ~n74317 ^ n74316;
  assign n74318 = ~n74322;
  assign n74320 = n74321 | n74318;
  assign n74325 = ~n74320 | ~n74319;
  assign n74323 = ~n74321;
  assign n74324 = n74323 | n74322;
  assign n74327 = n74325 & n74324;
  assign n74795 = ~n74865 | ~n74328;
  assign n74794 = ~n63296 | ~P4_DATAO_REG_21__SCAN_IN;
  assign n74333 = ~n74795 ^ n74794;
  assign n74331 = n74330 | n74329;
  assign n74334 = n74332 & n74331;
  assign n74340 = ~n74335;
  assign n74339 = ~n74336;
  assign n74338 = n74340 | n74339;
  assign n74342 = ~n74338 | ~n74337;
  assign n74341 = ~n74340 | ~n74339;
  assign n74878 = ~n74342 | ~n74341;
  assign n74876 = ~n74798 | ~P4_DATAO_REG_20__SCAN_IN;
  assign n74344 = ~n74878 ^ n74876;
  assign n74345 = ~n74344;
  assign n74347 = ~n74346 | ~n74345;
  assign n74891 = ~n74880 | ~n74347;
  assign n74350 = ~n74348;
  assign n74351 = ~n74350 | ~n74349;
  assign n74892 = ~n74352 | ~n74351;
  assign n74355 = ~n74891 ^ n74892;
  assign n74354 = ~n74353 & ~n74881;
  assign n74895 = ~n74355 | ~n74354;
  assign n74356 = n74355 | n74354;
  assign n74357 = ~n74895 | ~n74356;
  assign n74899 = n74358 | n74357;
  assign n74359 = ~n74358 | ~n74357;
  assign n74789 = ~n74899 | ~n74359;
  assign n74363 = ~n74362;
  assign n74365 = ~n74364 | ~n74363;
  assign n74904 = ~n74366 | ~n74365;
  assign n74369 = ~n63603 & ~n74367;
  assign n74907 = ~n74368 | ~n74369;
  assign n74371 = ~n74368;
  assign n74370 = ~n74369;
  assign n74372 = ~n74371 | ~n74370;
  assign n74917 = ~n74907 | ~n74372;
  assign n74375 = ~n61014 | ~n74374;
  assign n74916 = n74376 & n74375;
  assign n74379 = ~n74378 | ~n74377;
  assign n74923 = ~n74380 | ~n74379;
  assign n74919 = n64350 & P4_DATAO_REG_15__SCAN_IN;
  assign n74924 = n63929 & P4_DATAO_REG_14__SCAN_IN;
  assign n74381 = ~n74924;
  assign n74385 = ~n74919 ^ n74381;
  assign n74383 = n74923 | n74385;
  assign n74382 = ~n74923 | ~n74385;
  assign n74384 = ~n74383 | ~n74382;
  assign n74390 = ~n74915 | ~n74384;
  assign n74386 = ~n74385;
  assign n74388 = n74923 | n74386;
  assign n74387 = ~n74923 | ~n74386;
  assign n74389 = ~n74388 | ~n74387;
  assign n74392 = ~n74391;
  assign n74394 = n74393 | n74392;
  assign n74931 = ~n74395 | ~n74394;
  assign n74398 = ~n74932 ^ n74931;
  assign n74397 = ~n74396 & ~n76061;
  assign n74935 = ~n74398 | ~n74397;
  assign n74399 = ~n74411;
  assign n74413 = ~n74399 | ~n74409;
  assign n74401 = ~n74400;
  assign n74403 = ~n74402 | ~n74401;
  assign n74405 = ~n74413 | ~n74403;
  assign n74956 = ~n74404 | ~n74405;
  assign n74406 = ~n74405;
  assign n74408 = ~n74407 | ~n74406;
  assign n74958 = ~n74956 | ~n74408;
  assign n74410 = ~n74409;
  assign n74412 = ~n74411 | ~n74410;
  assign n74963 = ~n74413 | ~n74412;
  assign n74414 = n74960 | n76067;
  assign n74415 = ~n74414 | ~n76043;
  assign n74429 = ~n74963 & ~n74415;
  assign n74418 = n74960 | n76043;
  assign n74417 = ~n76067 & ~n76043;
  assign n74423 = ~n74417 & ~n74416;
  assign n74421 = n74418 & n74423;
  assign n74419 = n76067 & n76043;
  assign n74420 = ~n74960 | ~n74419;
  assign n74422 = ~n74421 | ~n74420;
  assign n74427 = ~n74963 | ~n74422;
  assign n74425 = ~n74960;
  assign n74424 = ~n74423;
  assign n74426 = ~n74425 | ~n74424;
  assign n74428 = ~n74427 | ~n74426;
  assign n74957 = ~n74429 & ~n74428;
  assign n75932 = ~n74958 ^ n74957;
  assign n74433 = ~n74432;
  assign n74435 = ~n74434 | ~n74433;
  assign n74439 = ~n74436;
  assign n74438 = ~n74437;
  assign n74441 = ~n74439 | ~n74438;
  assign n74970 = ~n76046 | ~P4_DATAO_REG_8__SCAN_IN;
  assign n75930 = ~n76076 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n74442 = ~n74970 ^ n75930;
  assign n74773 = ~n75933 ^ n74442;
  assign n74775 = ~n76064 & ~n76044;
  assign n74443 = ~n74773 ^ n74775;
  assign n74764 = ~n74774 ^ n74443;
  assign n74449 = ~n74446 | ~n74445;
  assign n74450 = ~n74449 | ~n74448;
  assign n74453 = ~n74452 | ~n74451;
  assign n74455 = ~n74454 | ~n74453;
  assign n74758 = ~n74457 | ~P4_DATAO_REG_3__SCAN_IN;
  assign n74751 = ~n74458 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n74459 = ~n74758 ^ n74751;
  assign n74750 = ~n74759 ^ n74459;
  assign n74461 = n74462 | n59988;
  assign n74464 = ~n74461 | ~n74460;
  assign n74465 = ~DIN_29_;
  assign n75064 = ~n74475 | ~n74474;
  assign n74477 = ~P1_P1_INSTQUEUE_REG_6__6__SCAN_IN | ~n59938;
  assign n74476 = ~P1_P1_INSTQUEUE_REG_11__6__SCAN_IN | ~n97185;
  assign n74481 = ~n74477 | ~n74476;
  assign n74479 = ~P1_P1_INSTQUEUE_REG_3__6__SCAN_IN | ~n97895;
  assign n74478 = ~P1_P1_INSTQUEUE_REG_5__6__SCAN_IN | ~n97303;
  assign n74480 = ~n74479 | ~n74478;
  assign n74489 = ~n74481 & ~n74480;
  assign n74483 = ~P1_P1_INSTQUEUE_REG_1__6__SCAN_IN | ~n75055;
  assign n74482 = ~P1_P1_INSTQUEUE_REG_9__6__SCAN_IN | ~n97979;
  assign n74487 = ~n74483 | ~n74482;
  assign n74485 = ~P1_P1_INSTQUEUE_REG_10__6__SCAN_IN | ~n97747;
  assign n74484 = ~P1_P1_INSTQUEUE_REG_2__6__SCAN_IN | ~n97746;
  assign n74486 = ~n74485 | ~n74484;
  assign n74488 = ~n74487 & ~n74486;
  assign n74505 = ~n74489 | ~n74488;
  assign n74491 = ~P1_P1_INSTQUEUE_REG_8__6__SCAN_IN | ~n59935;
  assign n74490 = ~P1_P1_INSTQUEUE_REG_13__6__SCAN_IN | ~n97754;
  assign n74495 = ~n74491 | ~n74490;
  assign n74493 = ~P1_P1_INSTQUEUE_REG_15__6__SCAN_IN | ~n97743;
  assign n74492 = ~P1_P1_INSTQUEUE_REG_7__6__SCAN_IN | ~n97225;
  assign n74494 = ~n74493 | ~n74492;
  assign n74503 = ~n74495 & ~n74494;
  assign n74497 = ~P1_P1_INSTQUEUE_REG_12__6__SCAN_IN | ~n97203;
  assign n74496 = ~P1_P1_INSTQUEUE_REG_4__6__SCAN_IN | ~n75033;
  assign n74501 = ~n74497 | ~n74496;
  assign n74499 = ~P1_P1_INSTQUEUE_REG_0__6__SCAN_IN | ~n97761;
  assign n74498 = ~P1_P1_INSTQUEUE_REG_14__6__SCAN_IN | ~n75052;
  assign n74500 = ~n74499 | ~n74498;
  assign n74502 = ~n74501 & ~n74500;
  assign n74504 = ~n74503 | ~n74502;
  assign n75065 = ~n74505 & ~n74504;
  assign n97721 = ~n97928;
  assign n74509 = ~n74508 & ~n97620;
  assign n74510 = ~n97721 & ~n74509;
  assign n75026 = ~n74510 | ~P1_P1_EAX_REG_29__SCAN_IN;
  assign n74729 = ~DIN_30_;
  assign n75020 = ~n75900 | ~n75899;
  assign n74731 = ~n74749 & ~n74737;
  assign n74740 = n74750 & n74731;
  assign n74734 = n74750 | n74733;
  assign n74736 = n76028 & P4_DATAO_REG_1__SCAN_IN;
  assign n74746 = ~n74736 | ~DIN_29_;
  assign n74745 = ~n74739 | ~n61577;
  assign n74741 = ~n74740;
  assign n76220 = ~n74746;
  assign n74742 = ~n74741 | ~n76220;
  assign n74744 = ~n60452 | ~n74743;
  assign n74748 = n74745 & n74744;
  assign n76217 = ~n74748 | ~n74747;
  assign n74755 = n74750 | n74749;
  assign n74753 = ~n74759 ^ n59986;
  assign n74752 = ~n74751;
  assign n74757 = ~n74756 | ~P4_DATAO_REG_2__SCAN_IN;
  assign n75019 = ~n76210 | ~n76213;
  assign n76205 = ~n74763 & ~n74762;
  assign n75018 = ~n76206 ^ n76205;
  assign n74765 = ~n74782;
  assign n74768 = ~n75002 ^ n75001;
  assign n74767 = ~n74766;
  assign n75910 = ~n74770 | ~n74769;
  assign n75906 = ~n74771 & ~n76082;
  assign n75901 = ~n76038 | ~P4_DATAO_REG_5__SCAN_IN;
  assign n74772 = ~n75906 ^ n75901;
  assign n75017 = ~n75910 ^ n74772;
  assign n74777 = ~n74774 ^ n74773;
  assign n74779 = ~n60759 | ~n74775;
  assign n74778 = ~n74777 | ~n74776;
  assign n75921 = ~n74779 | ~n74778;
  assign n75918 = ~n74780 | ~P4_DATAO_REG_7__SCAN_IN;
  assign n76194 = ~n75004 | ~P4_DATAO_REG_6__SCAN_IN;
  assign n74781 = ~n75918 ^ n76194;
  assign n74784 = ~n74783;
  assign n74786 = ~n74785 | ~n74784;
  assign n76197 = ~n74787 | ~n74786;
  assign n74791 = ~n74789;
  assign n74792 = ~n74791 | ~n74790;
  assign n76160 = ~n74793 | ~n74792;
  assign n76161 = ~n76037 | ~P4_DATAO_REG_17__SCAN_IN;
  assign n76159 = ~n76160 ^ n76161;
  assign n74796 = n74795 | n74794;
  assign n76114 = ~n74797 | ~n74796;
  assign n76112 = ~n74798 | ~P4_DATAO_REG_21__SCAN_IN;
  assign n74871 = ~n76114 ^ n76112;
  assign n74801 = ~n74800 | ~n74799;
  assign n76096 = ~n74802 | ~n74801;
  assign n74803 = ~DIN_0_ | ~P4_DATAO_REG_29__SCAN_IN;
  assign n76019 = ~n63317 & ~n74803;
  assign n74805 = ~n76019;
  assign n74809 = ~n74805 | ~P4_DATAO_REG_30__SCAN_IN;
  assign n74810 = ~P4_DATAO_REG_29__SCAN_IN;
  assign n74807 = ~n74810 & ~P4_DATAO_REG_30__SCAN_IN;
  assign n74808 = ~n74807 | ~n60375;
  assign n74814 = ~n74809 | ~n74808;
  assign n74811 = n74810 & n74277;
  assign n74813 = ~n74812 & ~n74811;
  assign n74816 = ~n74814 | ~n74813;
  assign n74815 = ~n60722 | ~P4_DATAO_REG_28__SCAN_IN;
  assign n75992 = n74816 | n74815;
  assign n74817 = ~n74816 | ~n74815;
  assign n74818 = ~n75992 | ~n74817;
  assign n75993 = n74818 | n74821;
  assign n74819 = ~n74818 | ~n74821;
  assign n76105 = ~n75993 | ~n74819;
  assign n76106 = ~n75994 & ~n74820;
  assign n74825 = ~n76105 ^ n76106;
  assign n74823 = ~n74822 | ~n74821;
  assign n74826 = ~n74824 | ~n74823;
  assign n76109 = ~n74825 | ~n74826;
  assign n74828 = ~n74825;
  assign n74827 = ~n74826;
  assign n74829 = ~n74828 | ~n74827;
  assign n76097 = ~n76109 | ~n74829;
  assign n76095 = ~n76096 ^ n76097;
  assign n76094 = ~n59908 | ~P4_DATAO_REG_26__SCAN_IN;
  assign n76127 = ~n76095 ^ n76094;
  assign n74833 = n74832 | n74831;
  assign n76126 = ~n74834 | ~n74833;
  assign n74836 = ~n76127 ^ n76126;
  assign n74837 = ~n74835 | ~P4_DATAO_REG_25__SCAN_IN;
  assign n76129 = n74836 | n74837;
  assign n74839 = ~n74836;
  assign n74838 = ~n74837;
  assign n74840 = n74839 | n74838;
  assign n76089 = ~n76129 | ~n74840;
  assign n74843 = ~n74841;
  assign n74844 = ~n74843 | ~n74842;
  assign n76090 = ~n74845 | ~n74844;
  assign n74848 = ~n76089 ^ n76090;
  assign n74847 = ~n76032 & ~n74846;
  assign n76093 = ~n74848 | ~n74847;
  assign n74849 = n74848 | n74847;
  assign n74850 = n76093 & n74849;
  assign n74851 = ~n75996 & ~n59984;
  assign n76147 = ~n74850 | ~n74851;
  assign n74853 = ~n74850;
  assign n74852 = ~n74851;
  assign n74854 = ~n74853 | ~n74852;
  assign n74860 = ~n76147 | ~n74854;
  assign n74857 = n74856 | n74855;
  assign n74859 = n74858 & n74857;
  assign n76146 = n74860 | n74859;
  assign n74861 = ~n74860 | ~n74859;
  assign n76117 = ~n76146 | ~n74861;
  assign n74864 = n74863 | n74862;
  assign n76118 = ~n74865 | ~n74864;
  assign n74866 = ~n76117 ^ n76118;
  assign n74867 = ~n60178 & ~n60217;
  assign n76121 = ~n74866 | ~n74867;
  assign n74869 = ~n74866;
  assign n74868 = ~n74867;
  assign n74870 = ~n74869 | ~n74868;
  assign n74872 = n76121 & n74870;
  assign n76116 = ~n74871 | ~n74872;
  assign n74874 = ~n74871;
  assign n74873 = ~n74872;
  assign n74875 = ~n74874 | ~n74873;
  assign n74887 = n76116 & n74875;
  assign n74877 = ~n74876;
  assign n74879 = ~n74878 | ~n74877;
  assign n74884 = ~n74880 | ~n74879;
  assign n74883 = ~n74882 & ~n74881;
  assign n76151 = ~n74884 | ~n74883;
  assign n74888 = ~n74885 | ~n76151;
  assign n74886 = ~n74888;
  assign n76150 = ~n74887 | ~n74886;
  assign n74889 = ~n74887;
  assign n74890 = ~n74889 | ~n74888;
  assign n76139 = ~n76150 | ~n74890;
  assign n76138 = ~n59930 | ~P4_DATAO_REG_19__SCAN_IN;
  assign n74893 = ~n74891;
  assign n74894 = ~n74893 | ~n74892;
  assign n76136 = ~n74895 | ~n74894;
  assign n76133 = ~n76137 ^ n76136;
  assign n74898 = ~n74897 | ~n74896;
  assign n76132 = ~n74899 | ~n74898;
  assign n74900 = ~n76133 ^ n76132;
  assign n74901 = ~n76054 | ~P4_DATAO_REG_18__SCAN_IN;
  assign n76135 = n74900 | n74901;
  assign n76158 = ~n76135 | ~n74902;
  assign n74909 = ~n76159 ^ n76158;
  assign n74905 = ~n74903;
  assign n74906 = ~n74905 | ~n74904;
  assign n74908 = ~n74907 | ~n74906;
  assign n75990 = ~n74909 | ~n74908;
  assign n74910 = n74909 | n74908;
  assign n74912 = ~n75990 | ~n74910;
  assign n74911 = ~n64350 | ~P4_DATAO_REG_16__SCAN_IN;
  assign n74913 = ~n74912 | ~n74911;
  assign n75985 = n63929 & P4_DATAO_REG_15__SCAN_IN;
  assign n74914 = ~n74919;
  assign n74922 = n74915 | n74914;
  assign n74918 = n74917 | n74916;
  assign n75982 = ~n74922 | ~n74918;
  assign n75979 = ~n75984 ^ n75982;
  assign n74921 = n74920 | n74919;
  assign n74927 = ~n74922 | ~n74921;
  assign n74926 = ~n74923;
  assign n74925 = ~n74927 | ~n74926;
  assign n74929 = ~n74925 | ~n74924;
  assign n74928 = n74927 | n74926;
  assign n75977 = ~n74929 | ~n74928;
  assign n75976 = ~n75979 ^ n75977;
  assign n75975 = ~n74930 | ~P4_DATAO_REG_14__SCAN_IN;
  assign n75967 = ~n75976 ^ n75975;
  assign n74933 = ~n74931;
  assign n74934 = n74933 | n74932;
  assign n75970 = ~n74935 | ~n74934;
  assign n75971 = ~n76051 | ~P4_DATAO_REG_13__SCAN_IN;
  assign n75968 = ~n75970 ^ n75971;
  assign n74941 = ~n75967 ^ n75968;
  assign n74947 = ~n74939 ^ n74937;
  assign n74936 = ~n74948;
  assign n74953 = ~n74947 | ~n74936;
  assign n74938 = ~n74937;
  assign n74940 = ~n74939 | ~n74938;
  assign n74942 = n74953 & n74940;
  assign n75965 = n74941 | n74942;
  assign n74944 = ~n74941;
  assign n74943 = ~n74942;
  assign n75925 = ~n74945 | ~n75965;
  assign n75961 = ~n76043 | ~P4_DATAO_REG_11__SCAN_IN;
  assign n75924 = ~n76067 | ~P4_DATAO_REG_12__SCAN_IN;
  assign n74946 = ~n75961 ^ n75924;
  assign n74949 = ~n74947;
  assign n74952 = ~n74949 | ~n74948;
  assign n74951 = ~n74950;
  assign n74954 = n74952 & n74951;
  assign n74955 = ~n74954 | ~n74953;
  assign n75950 = ~n74956 | ~n74955;
  assign n75954 = ~n76076 | ~P4_DATAO_REG_10__SCAN_IN;
  assign n74969 = ~n75950 ^ n75954;
  assign n74959 = ~n74957;
  assign n74968 = n74959 | n74958;
  assign n74961 = ~n74963 | ~n74962;
  assign n74965 = ~n74961 | ~n74960;
  assign n74964 = n74963 | n74962;
  assign n74966 = ~n74965 | ~n74964;
  assign n74967 = ~n74966 | ~n76043;
  assign n75953 = ~n74968 | ~n74967;
  assign n75928 = ~n74969 ^ n75953;
  assign n75931 = ~n75932 ^ n75933;
  assign n74983 = ~n75930;
  assign n74972 = ~n74976 | ~n74983;
  assign n74977 = ~n74970;
  assign n74971 = ~n74977 | ~n74983;
  assign n74973 = ~n74972 | ~n74971;
  assign n74975 = ~n75931 | ~n74973;
  assign n74974 = ~n74976 | ~n74977;
  assign n74981 = ~n75931;
  assign n74979 = ~n74976 | ~n75930;
  assign n74978 = ~n74977 | ~n75930;
  assign n74980 = ~n74979 | ~n74978;
  assign n74984 = ~n75933 | ~n74983;
  assign n75938 = ~n76056 & ~n76044;
  assign n76181 = ~n76046 | ~P4_DATAO_REG_9__SCAN_IN;
  assign n74991 = ~n75938 ^ n76181;
  assign n74985 = ~n74984 | ~n74991;
  assign n74990 = n75932 | n74985;
  assign n74986 = n74991 & n75930;
  assign n74988 = n75933 | n74986;
  assign n74993 = n74991 | n75930;
  assign n74987 = ~n75933 | ~n74993;
  assign n74989 = ~n74988 | ~n74987;
  assign n74997 = ~n74990 | ~n74989;
  assign n74992 = ~n74991;
  assign n74994 = ~n75933 | ~n74992;
  assign n74995 = ~n74994 | ~n74993;
  assign n74996 = n75932 & n74995;
  assign n74998 = ~n74997 & ~n74996;
  assign n74999 = ~n75941 ^ n74998;
  assign n76192 = ~n76182 ^ n74999;
  assign n75015 = ~n75000 ^ n76192;
  assign n75003 = ~n75001;
  assign n75013 = n75003 | n75002;
  assign n75011 = n75005 & n75004;
  assign n75009 = n75007 | n60640;
  assign n75010 = ~n75009 | ~n75008;
  assign n75012 = ~n75011 | ~n75010;
  assign n75014 = ~n75013 | ~n75012;
  assign n75916 = n75015 | n75014;
  assign n75016 = ~n75015 | ~n75014;
  assign n75915 = ~n75916 | ~n75016;
  assign n76204 = ~n75017 ^ n75915;
  assign n75075 = ~n77917 | ~n76224;
  assign n75023 = n75022 ^ n75021;
  assign n75025 = ~n75023 | ~n97648;
  assign n75024 = ~n97645 | ~P1_BUF1_REG_14__SCAN_IN;
  assign n97668 = ~n75025 | ~n75024;
  assign n98286 = ~n97668;
  assign n75073 = ~n98286 & ~n97630;
  assign n75071 = ~n97564 | ~P1_BUF1_REG_30__SCAN_IN;
  assign n75027 = ~n97929 | ~n75026;
  assign n76225 = ~n75027 | ~P1_P1_EAX_REG_30__SCAN_IN;
  assign n98287 = ~P1_P1_EAX_REG_30__SCAN_IN;
  assign n75029 = ~P1_P1_EAX_REG_29__SCAN_IN | ~n75028;
  assign n75030 = ~n98287 | ~n75029;
  assign n75069 = n76225 & n75030;
  assign n75032 = ~n97743 | ~P1_P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n75031 = ~P1_P1_INSTQUEUE_REG_6__7__SCAN_IN | ~n59938;
  assign n75037 = ~n75032 | ~n75031;
  assign n75035 = ~P1_P1_INSTQUEUE_REG_5__7__SCAN_IN | ~n97303;
  assign n75034 = ~P1_P1_INSTQUEUE_REG_4__7__SCAN_IN | ~n75033;
  assign n75036 = ~n75035 | ~n75034;
  assign n75045 = ~n75037 & ~n75036;
  assign n75039 = ~n97747 | ~P1_P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n75038 = ~n97225 | ~P1_P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n75043 = ~n75039 | ~n75038;
  assign n75041 = ~n97895 | ~P1_P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n75040 = ~n97746 | ~P1_P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n75042 = ~n75041 | ~n75040;
  assign n75044 = ~n75043 & ~n75042;
  assign n75063 = ~n75045 | ~n75044;
  assign n75047 = ~P1_P1_INSTQUEUE_REG_11__7__SCAN_IN | ~n97185;
  assign n75046 = ~n97761 | ~P1_P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n75051 = ~n75047 | ~n75046;
  assign n75049 = ~n59935 | ~P1_P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n75048 = ~P1_P1_INSTQUEUE_REG_9__7__SCAN_IN | ~n98034;
  assign n75050 = ~n75049 | ~n75048;
  assign n75061 = ~n75051 & ~n75050;
  assign n75054 = ~P1_P1_INSTQUEUE_REG_14__7__SCAN_IN | ~n75052;
  assign n75053 = ~n97754 | ~P1_P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n75059 = ~n75054 | ~n75053;
  assign n75057 = ~n97203 | ~P1_P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n75056 = ~n75055 | ~P1_P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n75058 = ~n75057 | ~n75056;
  assign n75060 = ~n75059 & ~n75058;
  assign n75062 = ~n75061 | ~n75060;
  assign n75067 = ~n75063 & ~n75062;
  assign n75066 = n75065 | n75064;
  assign n96922 = ~n75067 ^ n75066;
  assign n75068 = ~n98061 & ~n96922;
  assign n75070 = ~n75069 & ~n75068;
  assign n75072 = ~n75071 | ~n75070;
  assign n75074 = ~n75073 & ~n75072;
  assign P1_P1_U2721_Lock = ~n75075 | ~n75074;
  assign input_0 = keyinput_0 ^ SEL;
  assign input_1 = keyinput_1 ^ DIN_30_;
  assign AND_1 = input_0 & input_1;
  assign input_2 = keyinput_2 ^ DIN_29_;
  assign OR_2 = input_2 | AND_1;
  assign input_3 = keyinput_3 ^ DIN_28_;
  assign AND_3 = input_3 & OR_2;
  assign input_4 = keyinput_4 ^ DIN_27_;
  assign OR_4 = input_4 | AND_3;
  assign input_5 = keyinput_5 ^ DIN_26_;
  assign OR_5 = input_5 | OR_4;
  assign input_6 = keyinput_6 ^ DIN_25_;
  assign OR_6 = input_6 | OR_5;
  assign input_7 = ~keyinput_7 ^ DIN_24_;
  assign OR_7 = input_7 | OR_6;
  assign input_8 = keyinput_8 ^ DIN_23_;
  assign AND_8 = input_8 & OR_7;
  assign input_9 = ~keyinput_9 ^ DIN_22_;
  assign OR_9 = input_9 | AND_8;
  assign input_10 = keyinput_10 ^ DIN_21_;
  assign AND_10 = input_10 & OR_9;
  assign input_11 = ~keyinput_11 ^ DIN_20_;
  assign OR_11 = input_11 | AND_10;
  assign input_12 = keyinput_12 ^ DIN_19_;
  assign OR_12 = input_12 | OR_11;
  assign input_13 = ~keyinput_13 ^ DIN_18_;
  assign AND_13 = input_13 & OR_12;
  assign input_14 = ~keyinput_14 ^ DIN_17_;
  assign OR_14 = input_14 | AND_13;
  assign input_15 = ~keyinput_15 ^ DIN_16_;
  assign AND_15 = input_15 & OR_14;
  assign input_16 = keyinput_16 ^ DIN_15_;
  assign AND_16 = input_16 & AND_15;
  assign input_17 = ~keyinput_17 ^ DIN_14_;
  assign AND_17 = input_17 & AND_16;
  assign input_18 = keyinput_18 ^ DIN_13_;
  assign AND_18 = input_18 & AND_17;
  assign input_19 = keyinput_19 ^ DIN_12_;
  assign OR_19 = input_19 | AND_18;
  assign input_20 = keyinput_20 ^ DIN_11_;
  assign AND_20 = input_20 & OR_19;
  assign input_21 = ~keyinput_21 ^ DIN_10_;
  assign AND_21 = input_21 & AND_20;
  assign input_22 = ~keyinput_22 ^ DIN_9_;
  assign AND_22 = input_22 & AND_21;
  assign input_23 = keyinput_23 ^ DIN_8_;
  assign AND_23 = input_23 & AND_22;
  assign input_24 = ~keyinput_24 ^ DIN_7_;
  assign AND_24 = input_24 & AND_23;
  assign input_25 = keyinput_25 ^ DIN_6_;
  assign OR_25 = input_25 | AND_24;
  assign input_26 = ~keyinput_26 ^ DIN_5_;
  assign OR_26 = input_26 | OR_25;
  assign input_27 = keyinput_27 ^ DIN_4_;
  assign AND_27 = input_27 & OR_26;
  assign input_28 = ~keyinput_28 ^ DIN_3_;
  assign AND_28 = input_28 & AND_27;
  assign input_29 = keyinput_29 ^ DIN_2_;
  assign AND_29 = input_29 & AND_28;
  assign input_30 = ~keyinput_30 ^ DIN_1_;
  assign AND_30 = input_30 & AND_29;
  assign input_31 = ~keyinput_31 ^ DIN_0_;
  assign AND_31 = input_31 & AND_30;
  assign input_32 = keyinput_32 ^ P2_P1_ADS_N_REG_SCAN_IN;
  assign OR_32 = input_32 | AND_31;
  assign input_33 = ~keyinput_33 ^ P1_BUF1_REG_14__SCAN_IN;
  assign AND_33 = input_33 & OR_32;
  assign input_34 = keyinput_34 ^ P1_BUF1_REG_30__SCAN_IN;
  assign AND_34 = input_34 & AND_33;
  assign input_35 = ~keyinput_35 ^ P1_READY11_REG_SCAN_IN;
  assign OR_35 = input_35 | AND_34;
  assign input_36 = ~keyinput_36 ^ P4_DATAO_REG_0__SCAN_IN;
  assign OR_36 = input_36 | OR_35;
  assign input_37 = keyinput_37 ^ P4_DATAO_REG_1__SCAN_IN;
  assign AND_37 = input_37 & OR_36;
  assign input_38 = ~keyinput_38 ^ P4_DATAO_REG_2__SCAN_IN;
  assign AND_38 = input_38 & AND_37;
  assign input_39 = keyinput_39 ^ P4_DATAO_REG_3__SCAN_IN;
  assign AND_39 = input_39 & AND_38;
  assign input_40 = keyinput_40 ^ P4_DATAO_REG_4__SCAN_IN;
  assign AND_40 = input_40 & AND_39;
  assign input_41 = ~keyinput_41 ^ P4_DATAO_REG_5__SCAN_IN;
  assign AND_41 = input_41 & AND_40;
  assign input_42 = keyinput_42 ^ P4_DATAO_REG_6__SCAN_IN;
  assign AND_42 = input_42 & AND_41;
  assign input_43 = ~keyinput_43 ^ P4_DATAO_REG_7__SCAN_IN;
  assign AND_43 = input_43 & AND_42;
  assign input_44 = ~keyinput_44 ^ P4_DATAO_REG_8__SCAN_IN;
  assign AND_44 = input_44 & AND_43;
  assign input_45 = keyinput_45 ^ P4_DATAO_REG_9__SCAN_IN;
  assign AND_45 = input_45 & AND_44;
  assign input_46 = ~keyinput_46 ^ P4_DATAO_REG_10__SCAN_IN;
  assign AND_46 = input_46 & AND_45;
  assign input_47 = keyinput_47 ^ P4_DATAO_REG_11__SCAN_IN;
  assign AND_47 = input_47 & AND_46;
  assign input_48 = ~keyinput_48 ^ P4_DATAO_REG_12__SCAN_IN;
  assign OR_48 = input_48 | AND_47;
  assign input_49 = ~keyinput_49 ^ P4_DATAO_REG_13__SCAN_IN;
  assign AND_49 = input_49 & OR_48;
  assign input_50 = ~keyinput_50 ^ P4_DATAO_REG_14__SCAN_IN;
  assign AND_50 = input_50 & AND_49;
  assign input_51 = keyinput_51 ^ P4_DATAO_REG_15__SCAN_IN;
  assign AND_51 = input_51 & AND_50;
  assign input_52 = keyinput_52 ^ P4_DATAO_REG_16__SCAN_IN;
  assign AND_52 = input_52 & AND_51;
  assign input_53 = ~keyinput_53 ^ P4_DATAO_REG_17__SCAN_IN;
  assign AND_53 = input_53 & AND_52;
  assign input_54 = keyinput_54 ^ P4_DATAO_REG_18__SCAN_IN;
  assign OR_54 = input_54 | AND_53;
  assign input_55 = ~keyinput_55 ^ P4_DATAO_REG_19__SCAN_IN;
  assign OR_55 = input_55 | OR_54;
  assign input_56 = ~keyinput_56 ^ P4_DATAO_REG_20__SCAN_IN;
  assign OR_56 = input_56 | OR_55;
  assign input_57 = ~keyinput_57 ^ P4_DATAO_REG_21__SCAN_IN;
  assign OR_57 = input_57 | OR_56;
  assign input_58 = keyinput_58 ^ P4_DATAO_REG_22__SCAN_IN;
  assign AND_58 = input_58 & OR_57;
  assign input_59 = keyinput_59 ^ P4_DATAO_REG_23__SCAN_IN;
  assign OR_59 = input_59 | AND_58;
  assign input_60 = ~keyinput_60 ^ P4_DATAO_REG_24__SCAN_IN;
  assign OR_60 = input_60 | OR_59;
  assign input_61 = keyinput_61 ^ P4_DATAO_REG_25__SCAN_IN;
  assign OR_61 = input_61 | OR_60;
  assign input_62 = ~keyinput_62 ^ P4_DATAO_REG_26__SCAN_IN;
  assign OR_62 = input_62 | OR_61;
  assign input_63 = ~keyinput_63 ^ P4_DATAO_REG_27__SCAN_IN;
  assign OR_63 = input_63 | OR_62;
  assign input_64 = ~keyinput_64 ^ P4_DATAO_REG_28__SCAN_IN;
  assign AND_64 = input_64 & OR_63;
  assign input_65 = keyinput_65 ^ P4_DATAO_REG_29__SCAN_IN;
  assign OR_65 = input_65 | AND_64;
  assign input_66 = keyinput_66 ^ P4_DATAO_REG_30__SCAN_IN;
  assign AND_66 = input_66 & OR_65;
  assign input_67 = ~keyinput_67 ^ P1_P1_ADDRESS_REG_29__SCAN_IN;
  assign AND_67 = input_67 & AND_66;
  assign input_68 = keyinput_68 ^ P1_P1_ADDRESS_REG_28__SCAN_IN;
  assign OR_68 = input_68 | AND_67;
  assign input_69 = keyinput_69 ^ P1_P1_ADDRESS_REG_27__SCAN_IN;
  assign OR_69 = input_69 | OR_68;
  assign input_70 = keyinput_70 ^ P1_P1_ADDRESS_REG_26__SCAN_IN;
  assign OR_70 = input_70 | OR_69;
  assign input_71 = ~keyinput_71 ^ P1_P1_ADDRESS_REG_25__SCAN_IN;
  assign AND_71 = input_71 & OR_70;
  assign input_72 = ~keyinput_72 ^ P1_P1_ADDRESS_REG_24__SCAN_IN;
  assign OR_72 = input_72 | AND_71;
  assign input_73 = ~keyinput_73 ^ P1_P1_ADDRESS_REG_23__SCAN_IN;
  assign OR_73 = input_73 | OR_72;
  assign input_74 = keyinput_74 ^ P1_P1_ADDRESS_REG_22__SCAN_IN;
  assign AND_74 = input_74 & OR_73;
  assign input_75 = keyinput_75 ^ P1_P1_ADDRESS_REG_21__SCAN_IN;
  assign OR_75 = input_75 | AND_74;
  assign input_76 = keyinput_76 ^ P1_P1_ADDRESS_REG_20__SCAN_IN;
  assign AND_76 = input_76 & OR_75;
  assign input_77 = ~keyinput_77 ^ P1_P1_ADDRESS_REG_19__SCAN_IN;
  assign OR_77 = input_77 | AND_76;
  assign input_78 = keyinput_78 ^ P1_P1_ADDRESS_REG_18__SCAN_IN;
  assign OR_78 = input_78 | OR_77;
  assign input_79 = keyinput_79 ^ P1_P1_ADDRESS_REG_17__SCAN_IN;
  assign AND_79 = input_79 & OR_78;
  assign input_80 = keyinput_80 ^ SEL;
  assign input_81 = keyinput_81 ^ DIN_30_;
  assign AND_81 = input_80 & input_81;
  assign input_82 = keyinput_82 ^ DIN_29_;
  assign OR_82 = input_82 | AND_81;
  assign input_83 = keyinput_83 ^ DIN_28_;
  assign AND_83 = input_83 & OR_82;
  assign input_84 = keyinput_84 ^ DIN_27_;
  assign OR_84 = input_84 | AND_83;
  assign input_85 = ~keyinput_85 ^ DIN_26_;
  assign OR_85 = input_85 | OR_84;
  assign input_86 = ~keyinput_86 ^ DIN_25_;
  assign OR_86 = input_86 | OR_85;
  assign input_87 = ~keyinput_87 ^ DIN_24_;
  assign OR_87 = input_87 | OR_86;
  assign input_88 = keyinput_88 ^ DIN_23_;
  assign AND_88 = input_88 & OR_87;
  assign input_89 = ~keyinput_89 ^ DIN_22_;
  assign OR_89 = input_89 | AND_88;
  assign input_90 = keyinput_90 ^ DIN_21_;
  assign AND_90 = input_90 & OR_89;
  assign input_91 = keyinput_91 ^ DIN_20_;
  assign OR_91 = input_91 | AND_90;
  assign input_92 = ~keyinput_92 ^ DIN_19_;
  assign OR_92 = input_92 | OR_91;
  assign input_93 = keyinput_93 ^ DIN_18_;
  assign AND_93 = input_93 & OR_92;
  assign input_94 = keyinput_94 ^ DIN_17_;
  assign OR_94 = input_94 | AND_93;
  assign input_95 = ~keyinput_95 ^ DIN_16_;
  assign AND_95 = input_95 & OR_94;
  assign input_96 = ~keyinput_96 ^ DIN_15_;
  assign AND_96 = input_96 & AND_95;
  assign input_97 = ~keyinput_97 ^ DIN_14_;
  assign AND_97 = input_97 & AND_96;
  assign input_98 = ~keyinput_98 ^ DIN_13_;
  assign AND_98 = input_98 & AND_97;
  assign input_99 = ~keyinput_99 ^ DIN_12_;
  assign OR_99 = input_99 | AND_98;
  assign input_100 = keyinput_100 ^ DIN_11_;
  assign AND_100 = input_100 & OR_99;
  assign input_101 = keyinput_101 ^ DIN_10_;
  assign AND_101 = input_101 & AND_100;
  assign input_102 = ~keyinput_102 ^ DIN_9_;
  assign AND_102 = input_102 & AND_101;
  assign input_103 = keyinput_103 ^ DIN_8_;
  assign AND_103 = input_103 & AND_102;
  assign input_104 = keyinput_104 ^ DIN_7_;
  assign AND_104 = input_104 & AND_103;
  assign input_105 = ~keyinput_105 ^ DIN_6_;
  assign OR_105 = input_105 | AND_104;
  assign input_106 = ~keyinput_106 ^ DIN_5_;
  assign OR_106 = input_106 | OR_105;
  assign input_107 = ~keyinput_107 ^ DIN_4_;
  assign AND_107 = input_107 & OR_106;
  assign input_108 = ~keyinput_108 ^ DIN_3_;
  assign AND_108 = input_108 & AND_107;
  assign input_109 = keyinput_109 ^ DIN_2_;
  assign AND_109 = input_109 & AND_108;
  assign input_110 = keyinput_110 ^ DIN_1_;
  assign AND_110 = input_110 & AND_109;
  assign input_111 = keyinput_111 ^ DIN_0_;
  assign AND_111 = input_111 & AND_110;
  assign input_112 = keyinput_112 ^ P2_P1_ADS_N_REG_SCAN_IN;
  assign OR_112 = input_112 | AND_111;
  assign input_113 = ~keyinput_113 ^ P1_BUF1_REG_14__SCAN_IN;
  assign AND_113 = input_113 & OR_112;
  assign input_114 = keyinput_114 ^ P1_BUF1_REG_30__SCAN_IN;
  assign AND_114 = input_114 & AND_113;
  assign input_115 = ~keyinput_115 ^ P1_READY11_REG_SCAN_IN;
  assign OR_115 = input_115 | AND_114;
  assign input_116 = keyinput_116 ^ P4_DATAO_REG_0__SCAN_IN;
  assign OR_116 = input_116 | OR_115;
  assign input_117 = ~keyinput_117 ^ P4_DATAO_REG_1__SCAN_IN;
  assign AND_117 = input_117 & OR_116;
  assign input_118 = ~keyinput_118 ^ P4_DATAO_REG_2__SCAN_IN;
  assign AND_118 = input_118 & AND_117;
  assign input_119 = keyinput_119 ^ P4_DATAO_REG_3__SCAN_IN;
  assign AND_119 = input_119 & AND_118;
  assign input_120 = keyinput_120 ^ P4_DATAO_REG_4__SCAN_IN;
  assign AND_120 = input_120 & AND_119;
  assign input_121 = ~keyinput_121 ^ P4_DATAO_REG_5__SCAN_IN;
  assign AND_121 = input_121 & AND_120;
  assign input_122 = ~keyinput_122 ^ P4_DATAO_REG_6__SCAN_IN;
  assign AND_122 = input_122 & AND_121;
  assign input_123 = keyinput_123 ^ P4_DATAO_REG_7__SCAN_IN;
  assign AND_123 = input_123 & AND_122;
  assign input_124 = keyinput_124 ^ P4_DATAO_REG_8__SCAN_IN;
  assign AND_124 = input_124 & AND_123;
  assign input_125 = ~keyinput_125 ^ P4_DATAO_REG_9__SCAN_IN;
  assign AND_125 = input_125 & AND_124;
  assign input_126 = keyinput_126 ^ P4_DATAO_REG_10__SCAN_IN;
  assign AND_126 = input_126 & AND_125;
  assign input_127 = ~keyinput_127 ^ P4_DATAO_REG_11__SCAN_IN;
  assign AND_127 = input_127 & AND_126;
  assign input_128 = ~keyinput_128 ^ P4_DATAO_REG_12__SCAN_IN;
  assign OR_128 = input_128 | AND_127;
  assign input_129 = keyinput_129 ^ P4_DATAO_REG_13__SCAN_IN;
  assign AND_129 = input_129 & OR_128;
  assign input_130 = keyinput_130 ^ P4_DATAO_REG_14__SCAN_IN;
  assign AND_130 = input_130 & AND_129;
  assign input_131 = keyinput_131 ^ P4_DATAO_REG_15__SCAN_IN;
  assign AND_131 = input_131 & AND_130;
  assign input_132 = ~keyinput_132 ^ P4_DATAO_REG_16__SCAN_IN;
  assign AND_132 = input_132 & AND_131;
  assign input_133 = keyinput_133 ^ P4_DATAO_REG_17__SCAN_IN;
  assign AND_133 = input_133 & AND_132;
  assign input_134 = keyinput_134 ^ P4_DATAO_REG_18__SCAN_IN;
  assign OR_134 = input_134 | AND_133;
  assign input_135 = ~keyinput_135 ^ P4_DATAO_REG_19__SCAN_IN;
  assign OR_135 = input_135 | OR_134;
  assign input_136 = keyinput_136 ^ P4_DATAO_REG_20__SCAN_IN;
  assign OR_136 = input_136 | OR_135;
  assign input_137 = ~keyinput_137 ^ P4_DATAO_REG_21__SCAN_IN;
  assign OR_137 = input_137 | OR_136;
  assign input_138 = keyinput_138 ^ P4_DATAO_REG_22__SCAN_IN;
  assign AND_138 = input_138 & OR_137;
  assign input_139 = ~keyinput_139 ^ P4_DATAO_REG_23__SCAN_IN;
  assign OR_139 = input_139 | AND_138;
  assign input_140 = ~keyinput_140 ^ P4_DATAO_REG_24__SCAN_IN;
  assign OR_140 = input_140 | OR_139;
  assign input_141 = ~keyinput_141 ^ P4_DATAO_REG_25__SCAN_IN;
  assign OR_141 = input_141 | OR_140;
  assign input_142 = keyinput_142 ^ P4_DATAO_REG_26__SCAN_IN;
  assign OR_142 = input_142 | OR_141;
  assign input_143 = keyinput_143 ^ P4_DATAO_REG_27__SCAN_IN;
  assign OR_143 = input_143 | OR_142;
  assign input_144 = keyinput_144 ^ P4_DATAO_REG_28__SCAN_IN;
  assign AND_144 = input_144 & OR_143;
  assign input_145 = ~keyinput_145 ^ P4_DATAO_REG_29__SCAN_IN;
  assign OR_145 = input_145 | AND_144;
  assign input_146 = keyinput_146 ^ P4_DATAO_REG_30__SCAN_IN;
  assign AND_146 = input_146 & OR_145;
  assign input_147 = keyinput_147 ^ P1_P1_ADDRESS_REG_29__SCAN_IN;
  assign AND_147 = input_147 & AND_146;
  assign input_148 = keyinput_148 ^ P1_P1_ADDRESS_REG_28__SCAN_IN;
  assign OR_148 = input_148 | AND_147;
  assign input_149 = keyinput_149 ^ P1_P1_ADDRESS_REG_27__SCAN_IN;
  assign OR_149 = input_149 | OR_148;
  assign input_150 = keyinput_150 ^ P1_P1_ADDRESS_REG_26__SCAN_IN;
  assign OR_150 = input_150 | OR_149;
  assign input_151 = ~keyinput_151 ^ P1_P1_ADDRESS_REG_25__SCAN_IN;
  assign AND_151 = input_151 & OR_150;
  assign input_152 = keyinput_152 ^ P1_P1_ADDRESS_REG_24__SCAN_IN;
  assign OR_152 = input_152 | AND_151;
  assign input_153 = ~keyinput_153 ^ P1_P1_ADDRESS_REG_23__SCAN_IN;
  assign OR_153 = input_153 | OR_152;
  assign input_154 = ~keyinput_154 ^ P1_P1_ADDRESS_REG_22__SCAN_IN;
  assign AND_154 = input_154 & OR_153;
  assign input_155 = ~keyinput_155 ^ P1_P1_ADDRESS_REG_21__SCAN_IN;
  assign OR_155 = input_155 | AND_154;
  assign input_156 = ~keyinput_156 ^ P1_P1_ADDRESS_REG_20__SCAN_IN;
  assign AND_156 = input_156 & OR_155;
  assign input_157 = ~keyinput_157 ^ P1_P1_ADDRESS_REG_19__SCAN_IN;
  assign OR_157 = input_157 | AND_156;
  assign input_158 = keyinput_158 ^ P1_P1_ADDRESS_REG_18__SCAN_IN;
  assign OR_158 = input_158 | OR_157;
  assign input_159 = keyinput_159 ^ P1_P1_ADDRESS_REG_17__SCAN_IN;
  assign AND_159 = input_159 & OR_158;
  assign AND_159_INV = ~AND_159;
  assign CASOP = AND_79 & AND_159_INV;
  assign P1_P1_U2721 = P1_P1_U2721_Lock ^ CASOP;
endmodule


