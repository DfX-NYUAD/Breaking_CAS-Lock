// Benchmark "c432" written by ABC on Tue Feb  4 01:12:58 2020

module c432_10 ( 
    G1GAT, G4GAT, G8GAT, G11GAT, G14GAT, G17GAT, G21GAT, G24GAT, G27GAT,
    G30GAT, G34GAT, G37GAT, G40GAT, G43GAT, G47GAT, G50GAT, G53GAT, G56GAT,
    G60GAT, G63GAT, G66GAT, G69GAT, G73GAT, G76GAT, G79GAT, G82GAT, G86GAT,
    G89GAT, G92GAT, G95GAT, G99GAT, G102GAT, G105GAT, G108GAT, G112GAT,
    G115GAT,
    G223GAT, G329GAT, G370GAT, G421GAT, G430GAT, G431GAT, G432GAT  );
  input  G1GAT, G4GAT, G8GAT, G11GAT, G14GAT, G17GAT, G21GAT, G24GAT,
    G27GAT, G30GAT, G34GAT, G37GAT, G40GAT, G43GAT, G47GAT, G50GAT, G53GAT,
    G56GAT, G60GAT, G63GAT, G66GAT, G69GAT, G73GAT, G76GAT, G79GAT, G82GAT,
    G86GAT, G89GAT, G92GAT, G95GAT, G99GAT, G102GAT, G105GAT, G108GAT,
    G112GAT, G115GAT;
  output G223GAT, G329GAT, G370GAT, G421GAT, G430GAT, G431GAT, G432GAT;
  wire G118GAT, G119GAT, G122GAT, G123GAT, G126GAT, G127GAT, G130GAT,
    G131GAT, G134GAT, G135GAT, G138GAT, G139GAT, G142GAT, G143GAT, G146GAT,
    G147GAT, G150GAT, G151GAT, G154GAT, G157GAT, G158GAT, G159GAT, G162GAT,
    G165GAT, G168GAT, G171GAT, G174GAT, G177GAT, G180GAT, G183GAT, G184GAT,
    G185GAT, G186GAT, G187GAT, G188GAT, G189GAT, G190GAT, G191GAT, G192GAT,
    G193GAT, G194GAT, G195GAT, G196GAT, G197GAT, G198GAT, G199GAT, G203GAT,
    G213GAT, G224GAT, G227GAT, G230GAT, G233GAT, G236GAT, G239GAT, G242GAT,
    G243GAT, G246GAT, G247GAT, G250GAT, G251GAT, G254GAT, G255GAT, G256GAT,
    G257GAT, G258GAT, G259GAT, G260GAT, G263GAT, G264GAT, G267GAT, G270GAT,
    G273GAT, G276GAT, G279GAT, G282GAT, G285GAT, G288GAT, G289GAT, G290GAT,
    G291GAT, G292GAT, G293GAT, G294GAT, G295GAT, G296GAT, G300GAT, G301GAT,
    G302GAT, G303GAT, G304GAT, G305GAT, G306GAT, G307GAT, G308GAT, G309GAT,
    G319GAT, G330GAT, G331GAT, G332GAT, G333GAT, G334GAT, G335GAT, G336GAT,
    G337GAT, G338GAT, G339GAT, G340GAT, G341GAT, G342GAT, G343GAT, G344GAT,
    G345GAT, G346GAT, G347GAT, G348GAT, G349GAT, G350GAT, G351GAT, G352GAT,
    G353GAT, G354GAT, G355GAT, G356GAT, G357GAT, G360GAT, G371GAT, G372GAT,
    G373GAT, G374GAT, G375GAT, G376GAT, G377GAT, G378GAT, G379GAT, G380GAT,
    G381GAT, G386GAT, G393GAT, G399GAT, G404GAT, G407GAT, G411GAT, G414GAT,
    G415GAT, G416GAT, G417GAT, G418GAT, G419GAT, G420GAT, G422GAT, G425GAT,
    G428GAT, G429GAT;
  assign G118GAT = ~G1GAT;
  assign G119GAT = ~G4GAT;
  assign G122GAT = ~G11GAT;
  assign G123GAT = ~G17GAT;
  assign G126GAT = ~G24GAT;
  assign G127GAT = ~G30GAT;
  assign G130GAT = ~G37GAT;
  assign G131GAT = ~G43GAT;
  assign G134GAT = ~G50GAT;
  assign G135GAT = ~G56GAT;
  assign G138GAT = ~G63GAT;
  assign G139GAT = ~G69GAT;
  assign G142GAT = ~G76GAT;
  assign G143GAT = ~G82GAT;
  assign G146GAT = ~G89GAT;
  assign G147GAT = ~G95GAT;
  assign G150GAT = ~G102GAT;
  assign G151GAT = ~G108GAT;
  assign G154GAT = ~G118GAT | ~G4GAT;
  assign G157GAT = ~G8GAT & ~G119GAT;
  assign G158GAT = ~G14GAT & ~G119GAT;
  assign G159GAT = ~G122GAT | ~G17GAT;
  assign G162GAT = ~G126GAT | ~G30GAT;
  assign G165GAT = ~G130GAT | ~G43GAT;
  assign G168GAT = ~G134GAT | ~G56GAT;
  assign G171GAT = ~G138GAT | ~G69GAT;
  assign G174GAT = ~G142GAT | ~G82GAT;
  assign G177GAT = ~G146GAT | ~G95GAT;
  assign G180GAT = ~G150GAT | ~G108GAT;
  assign G183GAT = ~G21GAT & ~G123GAT;
  assign G184GAT = ~G27GAT & ~G123GAT;
  assign G185GAT = ~G34GAT & ~G127GAT;
  assign G186GAT = ~G40GAT & ~G127GAT;
  assign G187GAT = ~G47GAT & ~G131GAT;
  assign G188GAT = ~G53GAT & ~G131GAT;
  assign G189GAT = ~G60GAT & ~G135GAT;
  assign G190GAT = ~G66GAT & ~G135GAT;
  assign G191GAT = ~G73GAT & ~G139GAT;
  assign G192GAT = ~G79GAT & ~G139GAT;
  assign G193GAT = ~G86GAT & ~G143GAT;
  assign G194GAT = ~G92GAT & ~G143GAT;
  assign G195GAT = ~G99GAT & ~G147GAT;
  assign G196GAT = ~G105GAT & ~G147GAT;
  assign G197GAT = ~G112GAT & ~G151GAT;
  assign G198GAT = ~G115GAT & ~G151GAT;
  assign G199GAT = G180GAT & G177GAT & G174GAT & G171GAT & G168GAT & G165GAT & G162GAT & G154GAT & G159GAT;
  assign G203GAT = ~G199GAT;
  assign G213GAT = ~G199GAT;
  assign G223GAT = ~G199GAT;
  assign G224GAT = G203GAT ^ G154GAT;
  assign G227GAT = G203GAT ^ G159GAT;
  assign G230GAT = G203GAT ^ G162GAT;
  assign G233GAT = G203GAT ^ G165GAT;
  assign G236GAT = G203GAT ^ G168GAT;
  assign G239GAT = G203GAT ^ G171GAT;
  assign G242GAT = ~G1GAT | ~G213GAT;
  assign G243GAT = G203GAT ^ G174GAT;
  assign G246GAT = ~G213GAT | ~G11GAT;
  assign G247GAT = G203GAT ^ G177GAT;
  assign G250GAT = ~G213GAT | ~G24GAT;
  assign G251GAT = G203GAT ^ G180GAT;
  assign G254GAT = ~G213GAT | ~G37GAT;
  assign G255GAT = ~G213GAT | ~G50GAT;
  assign G256GAT = ~G213GAT | ~G63GAT;
  assign G257GAT = ~G213GAT | ~G76GAT;
  assign G258GAT = ~G213GAT | ~G89GAT;
  assign G259GAT = ~G213GAT | ~G102GAT;
  assign G260GAT = ~G224GAT | ~G157GAT;
  assign G263GAT = ~G224GAT | ~G158GAT;
  assign G264GAT = ~G227GAT | ~G183GAT;
  assign G267GAT = ~G230GAT | ~G185GAT;
  assign G270GAT = ~G233GAT | ~G187GAT;
  assign G273GAT = ~G236GAT | ~G189GAT;
  assign G276GAT = ~G239GAT | ~G191GAT;
  assign G279GAT = ~G243GAT | ~G193GAT;
  assign G282GAT = ~G247GAT | ~G195GAT;
  assign G285GAT = ~G251GAT | ~G197GAT;
  assign G288GAT = ~G227GAT | ~G184GAT;
  assign G289GAT = ~G230GAT | ~G186GAT;
  assign G290GAT = ~G233GAT | ~G188GAT;
  assign G291GAT = ~G236GAT | ~G190GAT;
  assign G292GAT = ~G239GAT | ~G192GAT;
  assign G293GAT = ~G243GAT | ~G194GAT;
  assign G294GAT = ~G247GAT | ~G196GAT;
  assign G295GAT = ~G251GAT | ~G198GAT;
  assign G296GAT = G285GAT & G282GAT & G279GAT & G276GAT & G273GAT & G270GAT & G267GAT & G260GAT & G264GAT;
  assign G300GAT = ~G263GAT;
  assign G301GAT = ~G288GAT;
  assign G302GAT = ~G289GAT;
  assign G303GAT = ~G290GAT;
  assign G304GAT = ~G291GAT;
  assign G305GAT = ~G292GAT;
  assign G306GAT = ~G293GAT;
  assign G307GAT = ~G294GAT;
  assign G308GAT = ~G295GAT;
  assign G309GAT = ~G296GAT;
  assign G319GAT = ~G296GAT;
  assign G329GAT = ~G296GAT;
  assign G330GAT = G309GAT ^ G260GAT;
  assign G331GAT = G309GAT ^ G264GAT;
  assign G332GAT = G309GAT ^ G267GAT;
  assign G333GAT = G309GAT ^ G270GAT;
  assign G334GAT = ~G8GAT | ~G319GAT;
  assign G335GAT = G309GAT ^ G273GAT;
  assign G336GAT = ~G319GAT | ~G21GAT;
  assign G337GAT = G309GAT ^ G276GAT;
  assign G338GAT = ~G319GAT | ~G34GAT;
  assign G339GAT = G309GAT ^ G279GAT;
  assign G340GAT = ~G319GAT | ~G47GAT;
  assign G341GAT = G309GAT ^ G282GAT;
  assign G342GAT = ~G319GAT | ~G60GAT;
  assign G343GAT = G309GAT ^ G285GAT;
  assign G344GAT = ~G319GAT | ~G73GAT;
  assign G345GAT = ~G319GAT | ~G86GAT;
  assign G346GAT = ~G319GAT | ~G99GAT;
  assign G347GAT = ~G319GAT | ~G112GAT;
  assign G348GAT = ~G330GAT | ~G300GAT;
  assign G349GAT = ~G331GAT | ~G301GAT;
  assign G350GAT = ~G332GAT | ~G302GAT;
  assign G351GAT = ~G333GAT | ~G303GAT;
  assign G352GAT = ~G335GAT | ~G304GAT;
  assign G353GAT = ~G337GAT | ~G305GAT;
  assign G354GAT = ~G339GAT | ~G306GAT;
  assign G355GAT = ~G341GAT | ~G307GAT;
  assign G356GAT = ~G343GAT | ~G308GAT;
  assign G357GAT = G356GAT & G355GAT & G354GAT & G353GAT & G352GAT & G351GAT & G350GAT & G348GAT & G349GAT;
  assign G360GAT = ~G357GAT;
  assign G370GAT = ~G357GAT;
  assign G371GAT = ~G14GAT | ~G360GAT;
  assign G372GAT = ~G360GAT | ~G27GAT;
  assign G373GAT = ~G360GAT | ~G40GAT;
  assign G374GAT = ~G360GAT | ~G53GAT;
  assign G375GAT = ~G360GAT | ~G66GAT;
  assign G376GAT = ~G360GAT | ~G79GAT;
  assign G377GAT = ~G360GAT | ~G92GAT;
  assign G378GAT = ~G360GAT | ~G105GAT;
  assign G379GAT = ~G360GAT | ~G115GAT;
  assign G380GAT = ~G371GAT | ~G334GAT | ~G4GAT | ~G242GAT;
  assign G381GAT = ~G17GAT | ~G372GAT | ~G246GAT | ~G336GAT;
  assign G386GAT = ~G30GAT | ~G373GAT | ~G250GAT | ~G338GAT;
  assign G393GAT = ~G43GAT | ~G374GAT | ~G254GAT | ~G340GAT;
  assign G399GAT = ~G56GAT | ~G375GAT | ~G255GAT | ~G342GAT;
  assign G404GAT = ~G69GAT | ~G376GAT | ~G256GAT | ~G344GAT;
  assign G407GAT = ~G82GAT | ~G377GAT | ~G257GAT | ~G345GAT;
  assign G411GAT = ~G95GAT | ~G378GAT | ~G258GAT | ~G346GAT;
  assign G414GAT = ~G108GAT | ~G379GAT | ~G259GAT | ~G347GAT;
  assign G415GAT = ~G380GAT;
  assign G416GAT = G414GAT & G411GAT & G407GAT & G404GAT & G399GAT & G393GAT & G381GAT & G386GAT;
  assign G417GAT = ~G393GAT;
  assign G418GAT = ~G404GAT;
  assign G419GAT = ~G407GAT;
  assign G420GAT = ~G411GAT;
  assign G421GAT = ~G415GAT & ~G416GAT;
  assign G422GAT = ~G386GAT | ~G417GAT;
  assign G425GAT = ~G399GAT | ~G418GAT | ~G386GAT | ~G393GAT;
  assign G428GAT = ~G419GAT | ~G399GAT | ~G393GAT;
  assign G429GAT = ~G420GAT | ~G407GAT | ~G386GAT | ~G393GAT;
  assign G430GAT = ~G399GAT | ~G422GAT | ~G381GAT | ~G386GAT;
  assign G431GAT = ~G428GAT | ~G425GAT | ~G381GAT | ~G386GAT;
  assign G432GAT = ~G429GAT | ~G425GAT | ~G381GAT | ~G422GAT;
endmodule


