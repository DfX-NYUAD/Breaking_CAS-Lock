// Benchmark "c1908" written by ABC on Thu Mar  5 01:06:14 2020

module c1908 ( 
    G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
    G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237,
    G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire G149, G153, G156, G160, G165, G168, G171, G175, G179, G184, G188,
    G191, G194, G198, G202, G206, G231, G233, G241, G244, G245, G248, G517,
    G529, G541, G553, G859, G862, G907, G909, G911, G918, G919, G922, G926,
    G930, G932, G934, G938, G943, G947, G949, G1506, G1514, G1522, G1530,
    G1538, G1546, G1554, G1562, G1570, G1578, G1586, G1594, G1602, G1610,
    G1618, G1626, G1512, G1520, G1528, G1536, G1544, G1552, G1560, G1568,
    G1576, G1584, G1592, G1600, G1608, G1616, G1624, G1632, G50, G52, G56,
    G58, G62, G64, G251, G254, G288, G291, G299, G302, G318, G321, G327,
    G330, G352, G355, G369, G382, G385, G853, G856, G893, G954, G955,
    G1050, G1053, G1176, G1179, G1197, G1207, G1222, G1244, G1278, G1290,
    G1300, G1312, G1332, G1335, G1442, G1450, G1458, G1466, G1474, G1482,
    G1490, G1498, G1634, G1644, G1657, G1665, G1697, G1705, G1713, G1721,
    G1745, G1753, G1785, G1793, G1814, G1817, G1830, G1833, G1841, G1849,
    G1854, G1857, G1870, G1873, G1878, G1881, G1642, G1652, G1056, G1057,
    G1182, G1183, G1211, G1298, G1320, G1338, G1339, G457, G459, G482,
    G487, G492, G505, G1456, G1448, G1472, G1464, G1488, G1480, G1504,
    G1496, G956, G967, G978, G979, G980, G1661, G990, G1669, G1030, G1701,
    G1040, G1709, G1058, G1717, G1068, G1725, G1078, G1090, G1100, G1749,
    G1112, G1757, G1154, G1789, G1166, G1797, G1194, G1201, G1204, G1820,
    G1821, G1230, G1836, G1837, G1252, G1256, G1845, G1268, G1853, G1860,
    G1861, G1286, G1876, G1877, G1308, G1884, G1885, G1654, G1662, G1694,
    G1702, G1710, G1718, G1726, G1734, G1742, G1750, G1782, G1790, G1838,
    G1846, G297, G298, G361, G362, G404, G405, G1225, G1226, G1247, G1248,
    G1281, G1282, G1303, G1304, G1315, G1316, G998, G988, G268, G1038,
    G1048, G1076, G1066, G1098, G1120, G1174, G363, G1210, G373, G1276,
    G406, G565, G566, G614, G615, G958, G969, G1660, G984, G1668, G994,
    G1700, G1034, G1708, G1044, G1716, G1062, G1724, G1072, G1732, G1086,
    G1740, G1748, G1104, G1108, G1756, G1116, G1788, G1158, G1162, G1796,
    G1170, G1200, G1203, G1227, G1249, G1844, G1260, G1264, G1852, G1272,
    G1283, G1305, G1317, G1410, G1418, G1426, G1434, G269, G372, G983,
    G993, G1033, G1043, G1061, G1071, G1103, G1115, G1157, G1169, G1184,
    G1202, G1259, G1271, G1322, G374, G396, G1321, G1424, G1416, G1440,
    G1432, G985, G995, G1035, G1045, G1063, G1073, G1105, G1117, G1159,
    G1171, G1212, G1231, G1232, G1253, G1254, G1261, G1273, G1287, G1288,
    G1309, G1310, G1192, G397, G1330, G1000, G1010, G1233, G1255, G1289,
    G1311, G1381, G257, G999, G260, G989, G272, G1039, G294, G1049, G305,
    G1077, G308, G1067, G333, G1121, G358, G1175, G1220, G388, G1277, G398,
    G1109, G1110, G1163, G1164, G1234, G1265, G1266, G1822, G1862, G1865,
    G258, G261, G273, G1018, G1008, G295, G306, G309, G334, G359, G389,
    G1385, G1111, G1165, G1267, G1886, G259, G262, G274, G296, G307, G310,
    G335, G360, G1242, G390, G1828, G1868, G1869, G1373, G1798, G1825,
    G265, G314, G336, G407, G1293, G1294, G1892, G1777, G1889, G410, G1377,
    G1804, G1237, G1829, G1295, G1670, G1678, G1729, G1737, G1761, G1769,
    G340, G343, G1781, G1238, G1325, G1893, G1340, G1352, G1673, G1681,
    G1801, G1897, G1905, G391, G1299, G1676, G1684, G1081, G1733, G1093,
    G1741, G1765, G1773, G1239, G1326, G1894, G1902, G392, G1360, G1003,
    G1677, G1013, G1685, G1082, G1094, G1122, G1134, G1187, G1805, G1327,
    G1901, G1348, G1909, G1758, G1766, G377, G1243, G393, G1004, G1014,
    G1083, G1095, G1188, G1900, G1344, G1908, G1356, G1142, G378, G399,
    G1331, G1005, G1015, G1764, G1126, G1130, G1772, G1138, G1189, G1343,
    G1355, G324, G1099, G379, G400, G449, G1087, G1088, G1125, G1137,
    G1345, G1357, G1397, G277, G1019, G280, G1009, G325, G364, G1193, G401,
    G1089, G1127, G1139, G278, G281, G326, G365, G413, G1361, G1401, G445,
    G1349, G1350, G1389, G1493, G1501, G1689, G279, G282, G346, G1143,
    G366, G414, G453, G1131, G1132, G1351, G1365, G1405, G285, G347, G367,
    G415, G1393, G556, G1505, G559, G1497, G1693, G1133, G1477, G1485,
    G1809, G348, G1369, G1409, G557, G560, G1362, G1378, G1429, G1437,
    G1686, G1774, G1910, G1918, G544, G1489, G547, G1481, G558, G561,
    G1813, G1370, G1368, G417, G1384, G424, G508, G1441, G511, G1433, G545,
    G548, G564, G1692, G1024, G1780, G1148, G1916, G1924, G416, G1376,
    G421, G423, G509, G512, G546, G549, G719, G722, G1023, G1147, G418,
    G420, G425, G510, G513, G552, G1025, G1149, G419, G422, G441, G516,
    G725, G728, G1029, G1153, G433, G437, G663, G666, G731, G746, G756,
    G770, G1461, G1469, G1413, G1421, G1445, G1453, G532, G1473, G535,
    G1465, G495, G1425, G498, G1417, G520, G1457, G523, G1449, G533, G536,
    G496, G499, G521, G524, G534, G537, G497, G500, G522, G525, G540, G503,
    G528, G669, G672, G569, G588, G618, G639, G867, G588A, G588B, G639A,
    G639B, G675, G688, G696, G710, G73, G572, G573, G621, G622, G776, G780,
    G784, G788, G812, G832, G836, G1509, G1517, G1525, G1533, G1581, G1621,
    G1629, G792, G796, G800, G804, G808, G816, G820, G824, G828, G871,
    G873, G875, G877, G879, G881, G883, G885, G1541, G1549, G1557, G1565,
    G1573, G1589, G1597, G1605, G1613, G1, G1513, G4, G1521, G7, G1529,
    G10, G1537, G28, G1585, G43, G1625, G46, G1633, G886, G2, G5, G8, G11,
    G13, G1545, G16, G1553, G19, G1561, G22, G1569, G25, G1577, G29, G31,
    G1593, G34, G1601, G37, G1609, G40, G1617, G44, G47, G857, G860, G863,
    G865, G14, G17, G20, G23, G26, G32, G35, G38, G41, G1913, G1921, G887,
    G462, G74, G1637, G1917, G1647, G1925, G1020, G1144, G1386, G1394,
    G1402, G1638, G1648, G1806, G1639, G1649, G287, G350, G427, G429, G431,
    G1028, G1152, G1392, G1400, G1408, G1812, G1216, G286, G349, G426,
    G428, G430, G67, G1643, G70, G1653, G1215, G49, G53, G59, G61, G65,
    G68, G71, G1217, G375, G1221, G376, G55;
  assign G149 = ~G101;
  assign G153 = ~G104;
  assign G156 = ~G107;
  assign G160 = ~G110;
  assign G165 = ~G113;
  assign G168 = ~G116;
  assign G171 = ~G119;
  assign G175 = ~G122;
  assign G179 = ~G125;
  assign G184 = ~G128;
  assign G188 = ~G131;
  assign G191 = ~G134;
  assign G194 = ~G137;
  assign G198 = ~G140;
  assign G202 = ~G143;
  assign G206 = ~G146;
  assign G231 = ~G224 | ~G898;
  assign G233 = ~G227 | ~G900;
  assign G241 = ~G237;
  assign G244 = ~G237;
  assign G245 = G234;
  assign G248 = G234;
  assign G517 = ~G469;
  assign G529 = ~G472;
  assign G541 = ~G475;
  assign G553 = ~G478;
  assign G859 = ~G953;
  assign G862 = ~G953;
  assign G907 = ~G898;
  assign G909 = ~G900;
  assign G911 = G902;
  assign G918 = ~G902;
  assign G919 = G902;
  assign G922 = ~G902;
  assign G926 = G952;
  assign G930 = ~G952;
  assign G932 = ~G952;
  assign G934 = G953;
  assign G938 = ~G953;
  assign G943 = G953;
  assign G947 = G953;
  assign G949 = ~G953;
  assign G1506 = G101;
  assign G1514 = G104;
  assign G1522 = G107;
  assign G1530 = G110;
  assign G1538 = G113;
  assign G1546 = G116;
  assign G1554 = G119;
  assign G1562 = G122;
  assign G1570 = G125;
  assign G1578 = G128;
  assign G1586 = G131;
  assign G1594 = G134;
  assign G1602 = G137;
  assign G1610 = G140;
  assign G1618 = G143;
  assign G1626 = G146;
  assign G1512 = ~G1506;
  assign G1520 = ~G1514;
  assign G1528 = ~G1522;
  assign G1536 = ~G1530;
  assign G1544 = ~G1538;
  assign G1552 = ~G1546;
  assign G1560 = ~G1554;
  assign G1568 = ~G1562;
  assign G1576 = ~G1570;
  assign G1584 = ~G1578;
  assign G1592 = ~G1586;
  assign G1600 = ~G1594;
  assign G1608 = ~G1602;
  assign G1616 = ~G1610;
  assign G1624 = ~G1618;
  assign G1632 = ~G1626;
  assign G50 = ~G930 | ~G947;
  assign G52 = ~G930 | ~G947;
  assign G56 = ~G930 | ~G947;
  assign G58 = ~G930 | ~G947;
  assign G62 = ~G930 | ~G947;
  assign G64 = ~G930 | ~G947;
  assign G251 = G149;
  assign G254 = G153;
  assign G288 = G165;
  assign G291 = G168;
  assign G299 = G184;
  assign G302 = G202;
  assign G318 = G224 & G938;
  assign G321 = G179;
  assign G327 = G188;
  assign G330 = G191;
  assign G352 = G227 & G938;
  assign G355 = G198;
  assign G369 = G938 & G210 & G241;
  assign G382 = G206;
  assign G385 = G198;
  assign G853 = ~G943 | ~G907;
  assign G856 = ~G943 | ~G909;
  assign G893 = ~G248 | ~G237;
  assign G954 = ~G248 | ~G922;
  assign G955 = ~G244 | ~G922;
  assign G1050 = G160;
  assign G1053 = G175;
  assign G1176 = G179;
  assign G1179 = G198;
  assign G1197 = G149;
  assign G1207 = G149;
  assign G1222 = G153;
  assign G1244 = G188;
  assign G1278 = G156;
  assign G1290 = G938 & G217 & G245;
  assign G1300 = G191;
  assign G1312 = G160;
  assign G1332 = G194;
  assign G1335 = G938 & G221 & G245;
  assign G1442 = G517;
  assign G1450 = G517;
  assign G1458 = G529;
  assign G1466 = G529;
  assign G1474 = G541;
  assign G1482 = G541;
  assign G1490 = G553;
  assign G1498 = G553;
  assign G1634 = G231 & G934;
  assign G1644 = G233 & G934;
  assign G1657 = G156;
  assign G1665 = G156;
  assign G1697 = G171;
  assign G1705 = G171;
  assign G1713 = G206;
  assign G1721 = G206;
  assign G1745 = G194;
  assign G1753 = G194;
  assign G1785 = G160;
  assign G1793 = G160;
  assign G1814 = G165;
  assign G1817 = G175;
  assign G1830 = G938 & G214 & G241;
  assign G1833 = G202;
  assign G1841 = G179;
  assign G1849 = G179;
  assign G1854 = G168;
  assign G1857 = G175;
  assign G1870 = G184;
  assign G1873 = G202;
  assign G1878 = G171;
  assign G1881 = G184;
  assign G1642 = ~G1634;
  assign G1652 = ~G1644;
  assign G1056 = ~G1050;
  assign G1057 = ~G1053;
  assign G1182 = ~G1176;
  assign G1183 = ~G1179;
  assign G1211 = ~G1207;
  assign G1298 = ~G1290;
  assign G1320 = ~G1312;
  assign G1338 = ~G1332;
  assign G1339 = ~G1335;
  assign G457 = G210 & G955;
  assign G459 = G217 & G954;
  assign G482 = ~G214 | ~G955;
  assign G487 = ~G221 | ~G954;
  assign G492 = ~G210 | ~G955;
  assign G505 = ~G217 | ~G954;
  assign G1456 = ~G1450;
  assign G1448 = ~G1442;
  assign G1472 = ~G1466;
  assign G1464 = ~G1458;
  assign G1488 = ~G1482;
  assign G1480 = ~G1474;
  assign G1504 = ~G1498;
  assign G1496 = ~G1490;
  assign G956 = ~G893 | ~G943 | ~G907 | ~G919;
  assign G967 = ~G893 | ~G943 | ~G909 | ~G919;
  assign G978 = ~G893 | ~G926 | ~G949;
  assign G979 = G893 & G926 & G949;
  assign G980 = G251;
  assign G1661 = ~G1657;
  assign G990 = G251;
  assign G1669 = ~G1665;
  assign G1030 = G288;
  assign G1701 = ~G1697;
  assign G1040 = G288;
  assign G1709 = ~G1705;
  assign G1058 = G299;
  assign G1717 = ~G1713;
  assign G1068 = G299;
  assign G1725 = ~G1721;
  assign G1078 = G318;
  assign G1090 = G318;
  assign G1100 = G327;
  assign G1749 = ~G1745;
  assign G1112 = G327;
  assign G1757 = ~G1753;
  assign G1154 = G352;
  assign G1789 = ~G1785;
  assign G1166 = G352;
  assign G1797 = ~G1793;
  assign G1194 = G369;
  assign G1201 = ~G1197;
  assign G1204 = G369;
  assign G1820 = ~G1814;
  assign G1821 = ~G1817;
  assign G1230 = ~G1222;
  assign G1836 = ~G1830;
  assign G1837 = ~G1833;
  assign G1252 = ~G1244;
  assign G1256 = G382;
  assign G1845 = ~G1841;
  assign G1268 = G382;
  assign G1853 = ~G1849;
  assign G1860 = ~G1854;
  assign G1861 = ~G1857;
  assign G1286 = ~G1278;
  assign G1876 = ~G1870;
  assign G1877 = ~G1873;
  assign G1308 = ~G1300;
  assign G1884 = ~G1878;
  assign G1885 = ~G1881;
  assign G1654 = G254;
  assign G1662 = G254;
  assign G1694 = G291;
  assign G1702 = G291;
  assign G1710 = G302;
  assign G1718 = G302;
  assign G1726 = G321;
  assign G1734 = G321;
  assign G1742 = G330;
  assign G1750 = G330;
  assign G1782 = G355;
  assign G1790 = G355;
  assign G1838 = G385;
  assign G1846 = G385;
  assign G297 = ~G1053 | ~G1056;
  assign G298 = ~G1050 | ~G1057;
  assign G361 = ~G1179 | ~G1182;
  assign G362 = ~G1176 | ~G1183;
  assign G404 = ~G1335 | ~G1338;
  assign G405 = ~G1332 | ~G1339;
  assign G1225 = ~G1817 | ~G1820;
  assign G1226 = ~G1814 | ~G1821;
  assign G1247 = ~G1833 | ~G1836;
  assign G1248 = ~G1830 | ~G1837;
  assign G1281 = ~G1857 | ~G1860;
  assign G1282 = ~G1854 | ~G1861;
  assign G1303 = ~G1873 | ~G1876;
  assign G1304 = ~G1870 | ~G1877;
  assign G1315 = ~G1881 | ~G1884;
  assign G1316 = ~G1878 | ~G1885;
  assign G998 = ~G990;
  assign G988 = ~G980;
  assign G268 = ~G297 | ~G298;
  assign G1038 = ~G1030;
  assign G1048 = ~G1040;
  assign G1076 = ~G1068;
  assign G1066 = ~G1058;
  assign G1098 = ~G1090;
  assign G1120 = ~G1112;
  assign G1174 = ~G1166;
  assign G363 = ~G361 | ~G362;
  assign G1210 = ~G1204;
  assign G373 = ~G1204 | ~G1211;
  assign G1276 = ~G1268;
  assign G406 = ~G404 | ~G405;
  assign G565 = ~G482;
  assign G566 = G482;
  assign G614 = ~G487;
  assign G615 = G487;
  assign G958 = ~G956 | ~G978;
  assign G969 = ~G967 | ~G978;
  assign G1660 = ~G1654;
  assign G984 = ~G1654 | ~G1661;
  assign G1668 = ~G1662;
  assign G994 = ~G1662 | ~G1669;
  assign G1700 = ~G1694;
  assign G1034 = ~G1694 | ~G1701;
  assign G1708 = ~G1702;
  assign G1044 = ~G1702 | ~G1709;
  assign G1716 = ~G1710;
  assign G1062 = ~G1710 | ~G1717;
  assign G1724 = ~G1718;
  assign G1072 = ~G1718 | ~G1725;
  assign G1732 = ~G1726;
  assign G1086 = ~G1078;
  assign G1740 = ~G1734;
  assign G1748 = ~G1742;
  assign G1104 = ~G1742 | ~G1749;
  assign G1108 = ~G1100;
  assign G1756 = ~G1750;
  assign G1116 = ~G1750 | ~G1757;
  assign G1788 = ~G1782;
  assign G1158 = ~G1782 | ~G1789;
  assign G1162 = ~G1154;
  assign G1796 = ~G1790;
  assign G1170 = ~G1790 | ~G1797;
  assign G1200 = ~G1194;
  assign G1203 = ~G1194 | ~G1201;
  assign G1227 = ~G1225 | ~G1226;
  assign G1249 = ~G1247 | ~G1248;
  assign G1844 = ~G1838;
  assign G1260 = ~G1838 | ~G1845;
  assign G1264 = ~G1256;
  assign G1852 = ~G1846;
  assign G1272 = ~G1846 | ~G1853;
  assign G1283 = ~G1281 | ~G1282;
  assign G1305 = ~G1303 | ~G1304;
  assign G1317 = ~G1315 | ~G1316;
  assign G1410 = G492;
  assign G1418 = G492;
  assign G1426 = G505;
  assign G1434 = G505;
  assign G269 = ~G268;
  assign G372 = ~G1207 | ~G1210;
  assign G983 = ~G1657 | ~G1660;
  assign G993 = ~G1665 | ~G1668;
  assign G1033 = ~G1697 | ~G1700;
  assign G1043 = ~G1705 | ~G1708;
  assign G1061 = ~G1713 | ~G1716;
  assign G1071 = ~G1721 | ~G1724;
  assign G1103 = ~G1745 | ~G1748;
  assign G1115 = ~G1753 | ~G1756;
  assign G1157 = ~G1785 | ~G1788;
  assign G1169 = ~G1793 | ~G1796;
  assign G1184 = ~G363;
  assign G1202 = ~G1197 | ~G1200;
  assign G1259 = ~G1841 | ~G1844;
  assign G1271 = ~G1849 | ~G1852;
  assign G1322 = ~G406;
  assign G374 = ~G372 | ~G373;
  assign G396 = ~G1317 | ~G1320;
  assign G1321 = ~G1317;
  assign G1424 = ~G1418;
  assign G1416 = ~G1410;
  assign G1440 = ~G1434;
  assign G1432 = ~G1426;
  assign G985 = ~G983 | ~G984;
  assign G995 = ~G993 | ~G994;
  assign G1035 = ~G1033 | ~G1034;
  assign G1045 = ~G1043 | ~G1044;
  assign G1063 = ~G1061 | ~G1062;
  assign G1073 = ~G1071 | ~G1072;
  assign G1105 = ~G1103 | ~G1104;
  assign G1117 = ~G1115 | ~G1116;
  assign G1159 = ~G1157 | ~G1158;
  assign G1171 = ~G1169 | ~G1170;
  assign G1212 = ~G1202 | ~G1203;
  assign G1231 = ~G1227;
  assign G1232 = ~G1227 | ~G1230;
  assign G1253 = ~G1249;
  assign G1254 = ~G1249 | ~G1252;
  assign G1261 = ~G1259 | ~G1260;
  assign G1273 = ~G1271 | ~G1272;
  assign G1287 = ~G1283;
  assign G1288 = ~G1283 | ~G1286;
  assign G1309 = ~G1305;
  assign G1310 = ~G1305 | ~G1308;
  assign G1192 = ~G1184;
  assign G397 = ~G1312 | ~G1321;
  assign G1330 = ~G1322;
  assign G1000 = G269;
  assign G1010 = G269;
  assign G1233 = ~G1222 | ~G1231;
  assign G1255 = ~G1244 | ~G1253;
  assign G1289 = ~G1278 | ~G1287;
  assign G1311 = ~G1300 | ~G1309;
  assign G1381 = ~G374;
  assign G257 = ~G995 | ~G998;
  assign G999 = ~G995;
  assign G260 = ~G985 | ~G988;
  assign G989 = ~G985;
  assign G272 = ~G1035 | ~G1038;
  assign G1039 = ~G1035;
  assign G294 = ~G1045 | ~G1048;
  assign G1049 = ~G1045;
  assign G305 = ~G1073 | ~G1076;
  assign G1077 = ~G1073;
  assign G308 = ~G1063 | ~G1066;
  assign G1067 = ~G1063;
  assign G333 = ~G1117 | ~G1120;
  assign G1121 = ~G1117;
  assign G358 = ~G1171 | ~G1174;
  assign G1175 = ~G1171;
  assign G1220 = ~G1212;
  assign G388 = ~G1273 | ~G1276;
  assign G1277 = ~G1273;
  assign G398 = ~G396 | ~G397;
  assign G1109 = ~G1105;
  assign G1110 = ~G1105 | ~G1108;
  assign G1163 = ~G1159;
  assign G1164 = ~G1159 | ~G1162;
  assign G1234 = ~G1232 | ~G1233;
  assign G1265 = ~G1261;
  assign G1266 = ~G1261 | ~G1264;
  assign G1822 = ~G1254 | ~G1255;
  assign G1862 = ~G1310 | ~G1311;
  assign G1865 = ~G1288 | ~G1289;
  assign G258 = ~G990 | ~G999;
  assign G261 = ~G980 | ~G989;
  assign G273 = ~G1030 | ~G1039;
  assign G1018 = ~G1010;
  assign G1008 = ~G1000;
  assign G295 = ~G1040 | ~G1049;
  assign G306 = ~G1068 | ~G1077;
  assign G309 = ~G1058 | ~G1067;
  assign G334 = ~G1112 | ~G1121;
  assign G359 = ~G1166 | ~G1175;
  assign G389 = ~G1268 | ~G1277;
  assign G1385 = ~G1381;
  assign G1111 = ~G1100 | ~G1109;
  assign G1165 = ~G1154 | ~G1163;
  assign G1267 = ~G1256 | ~G1265;
  assign G1886 = ~G398;
  assign G259 = ~G257 | ~G258;
  assign G262 = ~G260 | ~G261;
  assign G274 = ~G272 | ~G273;
  assign G296 = ~G294 | ~G295;
  assign G307 = ~G305 | ~G306;
  assign G310 = ~G308 | ~G309;
  assign G335 = ~G333 | ~G334;
  assign G360 = ~G358 | ~G359;
  assign G1242 = ~G1234;
  assign G390 = ~G388 | ~G389;
  assign G1828 = ~G1822;
  assign G1868 = ~G1862;
  assign G1869 = ~G1865;
  assign G1373 = ~G1164 | ~G1165;
  assign G1798 = ~G1110 | ~G1111;
  assign G1825 = ~G1266 | ~G1267;
  assign G265 = ~G259;
  assign G314 = ~G307;
  assign G336 = ~G335;
  assign G407 = ~G296;
  assign G1293 = ~G1865 | ~G1868;
  assign G1294 = ~G1862 | ~G1869;
  assign G1892 = ~G1886;
  assign G1777 = ~G360;
  assign G1889 = ~G390;
  assign G410 = G310;
  assign G1377 = ~G1373;
  assign G1804 = ~G1798;
  assign G1237 = ~G1825 | ~G1828;
  assign G1829 = ~G1825;
  assign G1295 = ~G1293 | ~G1294;
  assign G1670 = G274;
  assign G1678 = G274;
  assign G1729 = G310;
  assign G1737 = G310;
  assign G1761 = G262;
  assign G1769 = G262;
  assign G340 = G336;
  assign G343 = G314;
  assign G1781 = ~G1777;
  assign G1238 = ~G1822 | ~G1829;
  assign G1325 = ~G1889 | ~G1892;
  assign G1893 = ~G1889;
  assign G1340 = G407;
  assign G1352 = G407;
  assign G1673 = G265;
  assign G1681 = G265;
  assign G1801 = G314;
  assign G1897 = G336;
  assign G1905 = G336;
  assign G391 = ~G1295 | ~G1298;
  assign G1299 = ~G1295;
  assign G1676 = ~G1670;
  assign G1684 = ~G1678;
  assign G1081 = ~G1729 | ~G1732;
  assign G1733 = ~G1729;
  assign G1093 = ~G1737 | ~G1740;
  assign G1741 = ~G1737;
  assign G1765 = ~G1761;
  assign G1773 = ~G1769;
  assign G1239 = ~G1237 | ~G1238;
  assign G1326 = ~G1886 | ~G1893;
  assign G1894 = G410;
  assign G1902 = G410;
  assign G392 = ~G1290 | ~G1299;
  assign G1360 = ~G1352;
  assign G1003 = ~G1673 | ~G1676;
  assign G1677 = ~G1673;
  assign G1013 = ~G1681 | ~G1684;
  assign G1685 = ~G1681;
  assign G1082 = ~G1726 | ~G1733;
  assign G1094 = ~G1734 | ~G1741;
  assign G1122 = G340;
  assign G1134 = G340;
  assign G1187 = ~G1801 | ~G1804;
  assign G1805 = ~G1801;
  assign G1327 = ~G1325 | ~G1326;
  assign G1901 = ~G1897;
  assign G1348 = ~G1340;
  assign G1909 = ~G1905;
  assign G1758 = G343;
  assign G1766 = G343;
  assign G377 = ~G1239 | ~G1242;
  assign G1243 = ~G1239;
  assign G393 = ~G391 | ~G392;
  assign G1004 = ~G1670 | ~G1677;
  assign G1014 = ~G1678 | ~G1685;
  assign G1083 = ~G1081 | ~G1082;
  assign G1095 = ~G1093 | ~G1094;
  assign G1188 = ~G1798 | ~G1805;
  assign G1900 = ~G1894;
  assign G1344 = ~G1894 | ~G1901;
  assign G1908 = ~G1902;
  assign G1356 = ~G1902 | ~G1909;
  assign G1142 = ~G1134;
  assign G378 = ~G1234 | ~G1243;
  assign G399 = ~G1327 | ~G1330;
  assign G1331 = ~G1327;
  assign G1005 = ~G1003 | ~G1004;
  assign G1015 = ~G1013 | ~G1014;
  assign G1764 = ~G1758;
  assign G1126 = ~G1758 | ~G1765;
  assign G1130 = ~G1122;
  assign G1772 = ~G1766;
  assign G1138 = ~G1766 | ~G1773;
  assign G1189 = ~G1187 | ~G1188;
  assign G1343 = ~G1897 | ~G1900;
  assign G1355 = ~G1905 | ~G1908;
  assign G324 = ~G1095 | ~G1098;
  assign G1099 = ~G1095;
  assign G379 = ~G377 | ~G378;
  assign G400 = ~G1322 | ~G1331;
  assign G449 = ~G393 | ~G918;
  assign G1087 = ~G1083;
  assign G1088 = ~G1083 | ~G1086;
  assign G1125 = ~G1761 | ~G1764;
  assign G1137 = ~G1769 | ~G1772;
  assign G1345 = ~G1343 | ~G1344;
  assign G1357 = ~G1355 | ~G1356;
  assign G1397 = G393;
  assign G277 = ~G1015 | ~G1018;
  assign G1019 = ~G1015;
  assign G280 = ~G1005 | ~G1008;
  assign G1009 = ~G1005;
  assign G325 = ~G1090 | ~G1099;
  assign G364 = ~G1189 | ~G1192;
  assign G1193 = ~G1189;
  assign G401 = ~G399 | ~G400;
  assign G1089 = ~G1078 | ~G1087;
  assign G1127 = ~G1125 | ~G1126;
  assign G1139 = ~G1137 | ~G1138;
  assign G278 = ~G1010 | ~G1019;
  assign G281 = ~G1000 | ~G1009;
  assign G326 = ~G324 | ~G325;
  assign G365 = ~G1184 | ~G1193;
  assign G413 = ~G1357 | ~G1360;
  assign G1361 = ~G1357;
  assign G1401 = ~G1397;
  assign G445 = ~G379 | ~G918;
  assign G1349 = ~G1345;
  assign G1350 = ~G1345 | ~G1348;
  assign G1389 = G379;
  assign G1493 = G449;
  assign G1501 = G449;
  assign G1689 = ~G1088 | ~G1089;
  assign G279 = ~G277 | ~G278;
  assign G282 = ~G280 | ~G281;
  assign G346 = ~G1139 | ~G1142;
  assign G1143 = ~G1139;
  assign G366 = ~G364 | ~G365;
  assign G414 = ~G1352 | ~G1361;
  assign G453 = ~G401 | ~G918;
  assign G1131 = ~G1127;
  assign G1132 = ~G1127 | ~G1130;
  assign G1351 = ~G1340 | ~G1349;
  assign G1365 = ~G326;
  assign G1405 = G401;
  assign G285 = ~G279;
  assign G347 = ~G1134 | ~G1143;
  assign G367 = ~G366;
  assign G415 = ~G413 | ~G414;
  assign G1393 = ~G1389;
  assign G556 = ~G1501 | ~G1504;
  assign G1505 = ~G1501;
  assign G559 = ~G1493 | ~G1496;
  assign G1497 = ~G1493;
  assign G1693 = ~G1689;
  assign G1133 = ~G1122 | ~G1131;
  assign G1477 = G445;
  assign G1485 = G445;
  assign G1809 = ~G1350 | ~G1351;
  assign G348 = ~G346 | ~G347;
  assign G1369 = ~G1365;
  assign G1409 = ~G1405;
  assign G557 = ~G1498 | ~G1505;
  assign G560 = ~G1490 | ~G1497;
  assign G1362 = G282;
  assign G1378 = ~G415;
  assign G1429 = G453;
  assign G1437 = G453;
  assign G1686 = G282;
  assign G1774 = ~G1132 | ~G1133;
  assign G1910 = G285 & G853;
  assign G1918 = G856 & G367;
  assign G544 = ~G1485 | ~G1488;
  assign G1489 = ~G1485;
  assign G547 = ~G1477 | ~G1480;
  assign G1481 = ~G1477;
  assign G558 = ~G556 | ~G557;
  assign G561 = ~G559 | ~G560;
  assign G1813 = ~G1809;
  assign G1370 = ~G348;
  assign G1368 = ~G1362;
  assign G417 = ~G1362 | ~G1369;
  assign G1384 = ~G1378;
  assign G424 = ~G1378 | ~G1385;
  assign G508 = ~G1437 | ~G1440;
  assign G1441 = ~G1437;
  assign G511 = ~G1429 | ~G1432;
  assign G1433 = ~G1429;
  assign G545 = ~G1482 | ~G1489;
  assign G548 = ~G1474 | ~G1481;
  assign G564 = ~G558;
  assign G1692 = ~G1686;
  assign G1024 = ~G1686 | ~G1693;
  assign G1780 = ~G1774;
  assign G1148 = ~G1774 | ~G1781;
  assign G1916 = ~G1910;
  assign G1924 = ~G1918;
  assign G416 = ~G1365 | ~G1368;
  assign G1376 = ~G1370;
  assign G421 = ~G1370 | ~G1377;
  assign G423 = ~G1381 | ~G1384;
  assign G509 = ~G1434 | ~G1441;
  assign G512 = ~G1426 | ~G1433;
  assign G546 = ~G544 | ~G545;
  assign G549 = ~G547 | ~G548;
  assign G719 = ~G561;
  assign G722 = G561;
  assign G1023 = ~G1689 | ~G1692;
  assign G1147 = ~G1777 | ~G1780;
  assign G418 = ~G416 | ~G417;
  assign G420 = ~G1373 | ~G1376;
  assign G425 = ~G423 | ~G424;
  assign G510 = ~G508 | ~G509;
  assign G513 = ~G511 | ~G512;
  assign G552 = ~G546;
  assign G1025 = ~G1023 | ~G1024;
  assign G1149 = ~G1147 | ~G1148;
  assign G419 = ~G418;
  assign G422 = ~G420 | ~G421;
  assign G441 = ~G425 | ~G918;
  assign G516 = ~G510;
  assign G725 = ~G549;
  assign G728 = G549;
  assign G1029 = ~G1025;
  assign G1153 = ~G1149;
  assign G433 = ~G419 | ~G918;
  assign G437 = ~G422 | ~G918;
  assign G663 = ~G513;
  assign G666 = G513;
  assign G731 = G719 & G725;
  assign G746 = G722 & G725;
  assign G756 = G719 & G728;
  assign G770 = G722 & G728;
  assign G1461 = G441;
  assign G1469 = G441;
  assign G1413 = G433;
  assign G1421 = G433;
  assign G1445 = G437;
  assign G1453 = G437;
  assign G532 = ~G1469 | ~G1472;
  assign G1473 = ~G1469;
  assign G535 = ~G1461 | ~G1464;
  assign G1465 = ~G1461;
  assign G495 = ~G1421 | ~G1424;
  assign G1425 = ~G1421;
  assign G498 = ~G1413 | ~G1416;
  assign G1417 = ~G1413;
  assign G520 = ~G1453 | ~G1456;
  assign G1457 = ~G1453;
  assign G523 = ~G1445 | ~G1448;
  assign G1449 = ~G1445;
  assign G533 = ~G1466 | ~G1473;
  assign G536 = ~G1458 | ~G1465;
  assign G496 = ~G1418 | ~G1425;
  assign G499 = ~G1410 | ~G1417;
  assign G521 = ~G1450 | ~G1457;
  assign G524 = ~G1442 | ~G1449;
  assign G534 = ~G532 | ~G533;
  assign G537 = ~G535 | ~G536;
  assign G497 = ~G495 | ~G496;
  assign G500 = ~G498 | ~G499;
  assign G522 = ~G520 | ~G521;
  assign G525 = ~G523 | ~G524;
  assign G540 = ~G534;
  assign G503 = ~G497;
  assign G528 = ~G522;
  assign G669 = ~G537;
  assign G672 = G537;
  assign G569 = ~G500;
  assign G588 = G566 & G500;
  assign G618 = ~G525;
  assign G639 = G615 & G525;
  assign G867 = ~G487 | ~G503 | ~G528 | ~G482 | ~G540 | ~G552 | ~G516 | ~G564;
  assign G588A = G588;
  assign G588B = G588;
  assign G639A = G639;
  assign G639B = G639;
  assign G675 = G663 & G669;
  assign G688 = G666 & G669;
  assign G696 = G663 & G672;
  assign G710 = G666 & G672;
  assign G73 = G932 & G932 & G949 & G867;
  assign G572 = G565 & G569;
  assign G573 = G566 & G569;
  assign G621 = G614 & G618;
  assign G622 = G615 & G618;
  assign G776 = ~G958 | ~G731 | ~G696 | ~G588A | ~G639A;
  assign G780 = ~G958 | ~G756 | ~G675 | ~G588A | ~G639A;
  assign G784 = ~G958 | ~G746 | ~G675 | ~G588A | ~G639A;
  assign G788 = ~G958 | ~G731 | ~G688 | ~G588A | ~G639A;
  assign G812 = ~G969 | ~G746 | ~G710 | ~G588B | ~G639A;
  assign G832 = ~G969 | ~G770 | ~G696 | ~G588B | ~G639B;
  assign G836 = ~G969 | ~G756 | ~G710 | ~G588B | ~G639B;
  assign G1509 = G958 & G731 & G696 & G588A & G639A;
  assign G1517 = G958 & G756 & G675 & G588A & G639A;
  assign G1525 = G958 & G746 & G675 & G588A & G639A;
  assign G1533 = G958 & G731 & G688 & G588A & G639A;
  assign G1581 = G969 & G746 & G710 & G588B & G639A;
  assign G1621 = G969 & G770 & G696 & G588B & G639B;
  assign G1629 = G969 & G756 & G710 & G588B & G639B;
  assign G792 = ~G958 | ~G756 | ~G696 | ~G588A | ~G622;
  assign G796 = ~G958 | ~G746 | ~G696 | ~G588B | ~G622;
  assign G800 = ~G958 | ~G731 | ~G710 | ~G588B | ~G622;
  assign G804 = ~G958 | ~G770 | ~G675 | ~G588B | ~G622;
  assign G808 = ~G969 | ~G756 | ~G688 | ~G588B | ~G622;
  assign G816 = ~G969 | ~G756 | ~G696 | ~G573 | ~G639B;
  assign G820 = ~G969 | ~G746 | ~G696 | ~G573 | ~G639B;
  assign G824 = ~G969 | ~G731 | ~G710 | ~G573 | ~G639B;
  assign G828 = ~G969 | ~G756 | ~G688 | ~G573 | ~G639B;
  assign G871 = ~G979 | ~G731 | ~G675 | ~G588B | ~G622;
  assign G873 = ~G979 | ~G731 | ~G675 | ~G573 | ~G639B;
  assign G875 = ~G979 | ~G731 | ~G696 | ~G573 | ~G622;
  assign G877 = ~G979 | ~G756 | ~G675 | ~G573 | ~G622;
  assign G879 = ~G979 | ~G746 | ~G675 | ~G573 | ~G622;
  assign G881 = ~G979 | ~G731 | ~G688 | ~G573 | ~G622;
  assign G883 = ~G979 | ~G731 | ~G675 | ~G573 | ~G621;
  assign G885 = ~G979 | ~G731 | ~G675 | ~G572 | ~G622;
  assign G1541 = G958 & G756 & G696 & G588A & G622;
  assign G1549 = G958 & G746 & G696 & G588B & G622;
  assign G1557 = G958 & G731 & G710 & G588B & G622;
  assign G1565 = G958 & G770 & G675 & G588B & G622;
  assign G1573 = G969 & G756 & G688 & G588B & G622;
  assign G1589 = G969 & G756 & G696 & G573 & G639B;
  assign G1597 = G969 & G746 & G696 & G573 & G639B;
  assign G1605 = G969 & G731 & G710 & G573 & G639B;
  assign G1613 = G969 & G756 & G688 & G573 & G639B;
  assign G1 = ~G1509 | ~G1512;
  assign G1513 = ~G1509;
  assign G4 = ~G1517 | ~G1520;
  assign G1521 = ~G1517;
  assign G7 = ~G1525 | ~G1528;
  assign G1529 = ~G1525;
  assign G10 = ~G1533 | ~G1536;
  assign G1537 = ~G1533;
  assign G28 = ~G1581 | ~G1584;
  assign G1585 = ~G1581;
  assign G43 = ~G1621 | ~G1624;
  assign G1625 = ~G1621;
  assign G46 = ~G1629 | ~G1632;
  assign G1633 = ~G1629;
  assign G886 = G885 & G883 & G881 & G879 & G877 & G875 & G871 & G873;
  assign G2 = ~G1506 | ~G1513;
  assign G5 = ~G1514 | ~G1521;
  assign G8 = ~G1522 | ~G1529;
  assign G11 = ~G1530 | ~G1537;
  assign G13 = ~G1541 | ~G1544;
  assign G1545 = ~G1541;
  assign G16 = ~G1549 | ~G1552;
  assign G1553 = ~G1549;
  assign G19 = ~G1557 | ~G1560;
  assign G1561 = ~G1557;
  assign G22 = ~G1565 | ~G1568;
  assign G1569 = ~G1565;
  assign G25 = ~G1573 | ~G1576;
  assign G1577 = ~G1573;
  assign G29 = ~G1578 | ~G1585;
  assign G31 = ~G1589 | ~G1592;
  assign G1593 = ~G1589;
  assign G34 = ~G1597 | ~G1600;
  assign G1601 = ~G1597;
  assign G37 = ~G1605 | ~G1608;
  assign G1609 = ~G1605;
  assign G40 = ~G1613 | ~G1616;
  assign G1617 = ~G1613;
  assign G44 = ~G1618 | ~G1625;
  assign G47 = ~G1626 | ~G1633;
  assign G857 = ~G804 | ~G800 | ~G796 | ~G792 | ~G788 | ~G784 | ~G776 | ~G780;
  assign G860 = ~G836 | ~G832 | ~G828 | ~G824 | ~G820 | ~G816 | ~G808 | ~G812;
  assign G863 = G804 & G800 & G796 & G792 & G788 & G784 & G776 & G780;
  assign G865 = G836 & G832 & G828 & G824 & G820 & G816 & G808 & G812;
  assign G3 = ~G1 | ~G2;
  assign G6 = ~G4 | ~G5;
  assign G9 = ~G7 | ~G8;
  assign G12 = ~G10 | ~G11;
  assign G14 = ~G1538 | ~G1545;
  assign G17 = ~G1546 | ~G1553;
  assign G20 = ~G1554 | ~G1561;
  assign G23 = ~G1562 | ~G1569;
  assign G26 = ~G1570 | ~G1577;
  assign G30 = ~G28 | ~G29;
  assign G32 = ~G1586 | ~G1593;
  assign G35 = ~G1594 | ~G1601;
  assign G38 = ~G1602 | ~G1609;
  assign G41 = ~G1610 | ~G1617;
  assign G45 = ~G43 | ~G44;
  assign G48 = ~G46 | ~G47;
  assign G1913 = G857 & G859;
  assign G1921 = G860 & G862;
  assign G15 = ~G13 | ~G14;
  assign G18 = ~G16 | ~G17;
  assign G21 = ~G19 | ~G20;
  assign G24 = ~G22 | ~G23;
  assign G27 = ~G25 | ~G26;
  assign G33 = ~G31 | ~G32;
  assign G36 = ~G34 | ~G35;
  assign G39 = ~G37 | ~G38;
  assign G42 = ~G40 | ~G41;
  assign G887 = G886 & G863 & G865;
  assign G462 = ~G863 | ~G865;
  assign G74 = G887 & G952 & G949 & G867;
  assign G1637 = ~G1913 | ~G1916;
  assign G1917 = ~G1913;
  assign G1647 = ~G1921 | ~G1924;
  assign G1925 = ~G1921;
  assign G75 = ~G73 & ~G74;
  assign G1020 = G462 & G457 & G911;
  assign G1144 = G462 & G469 & G911;
  assign G1386 = G462 & G475 & G911;
  assign G1394 = G462 & G478 & G911;
  assign G1402 = G462 & G459 & G911;
  assign G1638 = ~G1910 | ~G1917;
  assign G1648 = ~G1918 | ~G1925;
  assign G1806 = G462 & G472 & G911;
  assign G1639 = ~G1637 | ~G1638;
  assign G1649 = ~G1647 | ~G1648;
  assign G287 = ~G1020 | ~G1029;
  assign G350 = ~G1144 | ~G1153;
  assign G427 = ~G1386 | ~G1393;
  assign G429 = ~G1394 | ~G1401;
  assign G431 = ~G1402 | ~G1409;
  assign G1028 = ~G1020;
  assign G1152 = ~G1144;
  assign G1392 = ~G1386;
  assign G1400 = ~G1394;
  assign G1408 = ~G1402;
  assign G1812 = ~G1806;
  assign G1216 = ~G1806 | ~G1813;
  assign G286 = ~G1025 | ~G1028;
  assign G349 = ~G1149 | ~G1152;
  assign G426 = ~G1389 | ~G1392;
  assign G428 = ~G1397 | ~G1400;
  assign G430 = ~G1405 | ~G1408;
  assign G67 = ~G1639 | ~G1642;
  assign G1643 = ~G1639;
  assign G70 = ~G1649 | ~G1652;
  assign G1653 = ~G1649;
  assign G1215 = ~G1809 | ~G1812;
  assign G49 = ~G286 | ~G287;
  assign G53 = ~G349 | ~G350;
  assign G59 = ~G426 | ~G427;
  assign G61 = ~G428 | ~G429;
  assign G65 = ~G430 | ~G431;
  assign G68 = ~G1634 | ~G1643;
  assign G71 = ~G1644 | ~G1653;
  assign G1217 = ~G1215 | ~G1216;
  assign G51 = G49 & G50;
  assign G54 = G52 & G53;
  assign G60 = G58 & G59;
  assign G63 = G61 & G62;
  assign G66 = G64 & G65;
  assign G69 = ~G67 | ~G68;
  assign G72 = ~G70 | ~G71;
  assign G375 = ~G1217 | ~G1220;
  assign G1221 = ~G1217;
  assign G376 = ~G1212 | ~G1221;
  assign G55 = ~G375 | ~G376;
  assign G57 = G55 & G56;
endmodule


