// Benchmark "c1355" written by ABC on Thu Mar  5 01:05:54 2020

module c1355 ( 
    G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
    G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
    G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT,
    G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT,
    G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT,
    G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
    G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
    G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
    G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
    G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT,
    G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT,
    G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
    G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT,
    G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT,
    G233GAT;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
    G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
    G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
    G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
    G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire G242GAT, G245GAT, G248GAT, G251GAT, G254GAT, G257GAT, G260GAT,
    G263GAT, G266GAT, G269GAT, G272GAT, G275GAT, G278GAT, G281GAT, G284GAT,
    G287GAT, G290GAT, G293GAT, G296GAT, G299GAT, G302GAT, G305GAT, G308GAT,
    G311GAT, G314GAT, G317GAT, G320GAT, G323GAT, G326GAT, G329GAT, G332GAT,
    G335GAT, G338GAT, G341GAT, G344GAT, G347GAT, G350GAT, G353GAT, G356GAT,
    G359GAT, G362GAT, G363GAT, G364GAT, G365GAT, G366GAT, G367GAT, G368GAT,
    G369GAT, G370GAT, G371GAT, G372GAT, G373GAT, G374GAT, G375GAT, G376GAT,
    G377GAT, G378GAT, G379GAT, G380GAT, G381GAT, G382GAT, G383GAT, G384GAT,
    G385GAT, G386GAT, G387GAT, G388GAT, G389GAT, G390GAT, G391GAT, G392GAT,
    G393GAT, G394GAT, G395GAT, G396GAT, G397GAT, G398GAT, G399GAT, G400GAT,
    G401GAT, G402GAT, G403GAT, G404GAT, G405GAT, G406GAT, G407GAT, G408GAT,
    G409GAT, G410GAT, G411GAT, G412GAT, G413GAT, G414GAT, G415GAT, G416GAT,
    G417GAT, G418GAT, G419GAT, G420GAT, G421GAT, G422GAT, G423GAT, G424GAT,
    G425GAT, G426GAT, G429GAT, G432GAT, G435GAT, G438GAT, G441GAT, G444GAT,
    G447GAT, G450GAT, G453GAT, G456GAT, G459GAT, G462GAT, G465GAT, G468GAT,
    G471GAT, G474GAT, G477GAT, G480GAT, G483GAT, G486GAT, G489GAT, G492GAT,
    G495GAT, G498GAT, G501GAT, G504GAT, G507GAT, G510GAT, G513GAT, G516GAT,
    G519GAT, G522GAT, G525GAT, G528GAT, G531GAT, G534GAT, G537GAT, G540GAT,
    G543GAT, G546GAT, G549GAT, G552GAT, G555GAT, G558GAT, G561GAT, G564GAT,
    G567GAT, G570GAT, G571GAT, G572GAT, G573GAT, G574GAT, G575GAT, G576GAT,
    G577GAT, G578GAT, G579GAT, G580GAT, G581GAT, G582GAT, G583GAT, G584GAT,
    G585GAT, G586GAT, G587GAT, G588GAT, G589GAT, G590GAT, G591GAT, G592GAT,
    G593GAT, G594GAT, G595GAT, G596GAT, G597GAT, G598GAT, G599GAT, G600GAT,
    G601GAT, G602GAT, G607GAT, G612GAT, G617GAT, G622GAT, G627GAT, G632GAT,
    G637GAT, G642GAT, G645GAT, G648GAT, G651GAT, G654GAT, G657GAT, G660GAT,
    G663GAT, G666GAT, G669GAT, G672GAT, G675GAT, G678GAT, G681GAT, G684GAT,
    G687GAT, G690GAT, G691GAT, G692GAT, G693GAT, G694GAT, G695GAT, G696GAT,
    G697GAT, G698GAT, G699GAT, G700GAT, G701GAT, G702GAT, G703GAT, G704GAT,
    G705GAT, G706GAT, G709GAT, G712GAT, G715GAT, G718GAT, G721GAT, G724GAT,
    G727GAT, G730GAT, G733GAT, G736GAT, G739GAT, G742GAT, G745GAT, G748GAT,
    G751GAT, G754GAT, G755GAT, G756GAT, G757GAT, G758GAT, G759GAT, G760GAT,
    G761GAT, G762GAT, G763GAT, G764GAT, G765GAT, G766GAT, G767GAT, G768GAT,
    G769GAT, G770GAT, G773GAT, G776GAT, G779GAT, G782GAT, G785GAT, G788GAT,
    G791GAT, G794GAT, G797GAT, G800GAT, G803GAT, G806GAT, G809GAT, G812GAT,
    G815GAT, G818GAT, G819GAT, G820GAT, G821GAT, G822GAT, G823GAT, G824GAT,
    G825GAT, G826GAT, G827GAT, G828GAT, G829GAT, G830GAT, G831GAT, G832GAT,
    G833GAT, G834GAT, G847GAT, G860GAT, G873GAT, G886GAT, G899GAT, G912GAT,
    G925GAT, G938GAT, G939GAT, G940GAT, G941GAT, G942GAT, G943GAT, G944GAT,
    G945GAT, G946GAT, G947GAT, G948GAT, G949GAT, G950GAT, G951GAT, G952GAT,
    G953GAT, G954GAT, G955GAT, G956GAT, G957GAT, G958GAT, G959GAT, G960GAT,
    G961GAT, G962GAT, G963GAT, G964GAT, G965GAT, G966GAT, G967GAT, G968GAT,
    G969GAT, G970GAT, G971GAT, G972GAT, G973GAT, G974GAT, G975GAT, G976GAT,
    G977GAT, G978GAT, G979GAT, G980GAT, G981GAT, G982GAT, G983GAT, G984GAT,
    G985GAT, G986GAT, G991GAT, G996GAT, G1001GAT, G1006GAT, G1011GAT,
    G1016GAT, G1021GAT, G1026GAT, G1031GAT, G1036GAT, G1039GAT, G1042GAT,
    G1045GAT, G1048GAT, G1051GAT, G1054GAT, G1057GAT, G1060GAT, G1063GAT,
    G1066GAT, G1069GAT, G1072GAT, G1075GAT, G1078GAT, G1081GAT, G1084GAT,
    G1087GAT, G1090GAT, G1093GAT, G1096GAT, G1099GAT, G1102GAT, G1105GAT,
    G1108GAT, G1111GAT, G1114GAT, G1117GAT, G1120GAT, G1123GAT, G1126GAT,
    G1129GAT, G1132GAT, G1135GAT, G1138GAT, G1141GAT, G1144GAT, G1147GAT,
    G1150GAT, G1153GAT, G1156GAT, G1159GAT, G1162GAT, G1165GAT, G1168GAT,
    G1171GAT, G1174GAT, G1177GAT, G1180GAT, G1183GAT, G1186GAT, G1189GAT,
    G1192GAT, G1195GAT, G1198GAT, G1201GAT, G1204GAT, G1207GAT, G1210GAT,
    G1213GAT, G1216GAT, G1219GAT, G1222GAT, G1225GAT, G1228GAT, G1229GAT,
    G1230GAT, G1231GAT, G1232GAT, G1233GAT, G1234GAT, G1235GAT, G1236GAT,
    G1237GAT, G1238GAT, G1239GAT, G1240GAT, G1241GAT, G1242GAT, G1243GAT,
    G1244GAT, G1245GAT, G1246GAT, G1247GAT, G1248GAT, G1249GAT, G1250GAT,
    G1251GAT, G1252GAT, G1253GAT, G1254GAT, G1255GAT, G1256GAT, G1257GAT,
    G1258GAT, G1259GAT, G1260GAT, G1261GAT, G1262GAT, G1263GAT, G1264GAT,
    G1265GAT, G1266GAT, G1267GAT, G1268GAT, G1269GAT, G1270GAT, G1271GAT,
    G1272GAT, G1273GAT, G1274GAT, G1275GAT, G1276GAT, G1277GAT, G1278GAT,
    G1279GAT, G1280GAT, G1281GAT, G1282GAT, G1283GAT, G1284GAT, G1285GAT,
    G1286GAT, G1287GAT, G1288GAT, G1289GAT, G1290GAT, G1291GAT, G1292GAT,
    G1293GAT, G1294GAT, G1295GAT, G1296GAT, G1297GAT, G1298GAT, G1299GAT,
    G1300GAT, G1301GAT, G1302GAT, G1303GAT, G1304GAT, G1305GAT, G1306GAT,
    G1307GAT, G1308GAT, G1309GAT, G1310GAT, G1311GAT, G1312GAT, G1313GAT,
    G1314GAT, G1315GAT, G1316GAT, G1317GAT, G1318GAT, G1319GAT, G1320GAT,
    G1321GAT, G1322GAT, G1323GAT;
  assign G242GAT = G225GAT & G233GAT;
  assign G245GAT = G226GAT & G233GAT;
  assign G248GAT = G227GAT & G233GAT;
  assign G251GAT = G228GAT & G233GAT;
  assign G254GAT = G229GAT & G233GAT;
  assign G257GAT = G230GAT & G233GAT;
  assign G260GAT = G231GAT & G233GAT;
  assign G263GAT = G232GAT & G233GAT;
  assign G266GAT = ~G1GAT | ~G8GAT;
  assign G269GAT = ~G15GAT | ~G22GAT;
  assign G272GAT = ~G29GAT | ~G36GAT;
  assign G275GAT = ~G43GAT | ~G50GAT;
  assign G278GAT = ~G57GAT | ~G64GAT;
  assign G281GAT = ~G71GAT | ~G78GAT;
  assign G284GAT = ~G85GAT | ~G92GAT;
  assign G287GAT = ~G99GAT | ~G106GAT;
  assign G290GAT = ~G113GAT | ~G120GAT;
  assign G293GAT = ~G127GAT | ~G134GAT;
  assign G296GAT = ~G141GAT | ~G148GAT;
  assign G299GAT = ~G155GAT | ~G162GAT;
  assign G302GAT = ~G169GAT | ~G176GAT;
  assign G305GAT = ~G183GAT | ~G190GAT;
  assign G308GAT = ~G197GAT | ~G204GAT;
  assign G311GAT = ~G211GAT | ~G218GAT;
  assign G314GAT = ~G1GAT | ~G29GAT;
  assign G317GAT = ~G57GAT | ~G85GAT;
  assign G320GAT = ~G8GAT | ~G36GAT;
  assign G323GAT = ~G64GAT | ~G92GAT;
  assign G326GAT = ~G15GAT | ~G43GAT;
  assign G329GAT = ~G71GAT | ~G99GAT;
  assign G332GAT = ~G22GAT | ~G50GAT;
  assign G335GAT = ~G78GAT | ~G106GAT;
  assign G338GAT = ~G113GAT | ~G141GAT;
  assign G341GAT = ~G169GAT | ~G197GAT;
  assign G344GAT = ~G120GAT | ~G148GAT;
  assign G347GAT = ~G176GAT | ~G204GAT;
  assign G350GAT = ~G127GAT | ~G155GAT;
  assign G353GAT = ~G183GAT | ~G211GAT;
  assign G356GAT = ~G134GAT | ~G162GAT;
  assign G359GAT = ~G190GAT | ~G218GAT;
  assign G362GAT = ~G1GAT | ~G266GAT;
  assign G363GAT = ~G8GAT | ~G266GAT;
  assign G364GAT = ~G15GAT | ~G269GAT;
  assign G365GAT = ~G22GAT | ~G269GAT;
  assign G366GAT = ~G29GAT | ~G272GAT;
  assign G367GAT = ~G36GAT | ~G272GAT;
  assign G368GAT = ~G43GAT | ~G275GAT;
  assign G369GAT = ~G50GAT | ~G275GAT;
  assign G370GAT = ~G57GAT | ~G278GAT;
  assign G371GAT = ~G64GAT | ~G278GAT;
  assign G372GAT = ~G71GAT | ~G281GAT;
  assign G373GAT = ~G78GAT | ~G281GAT;
  assign G374GAT = ~G85GAT | ~G284GAT;
  assign G375GAT = ~G92GAT | ~G284GAT;
  assign G376GAT = ~G99GAT | ~G287GAT;
  assign G377GAT = ~G106GAT | ~G287GAT;
  assign G378GAT = ~G113GAT | ~G290GAT;
  assign G379GAT = ~G120GAT | ~G290GAT;
  assign G380GAT = ~G127GAT | ~G293GAT;
  assign G381GAT = ~G134GAT | ~G293GAT;
  assign G382GAT = ~G141GAT | ~G296GAT;
  assign G383GAT = ~G148GAT | ~G296GAT;
  assign G384GAT = ~G155GAT | ~G299GAT;
  assign G385GAT = ~G162GAT | ~G299GAT;
  assign G386GAT = ~G169GAT | ~G302GAT;
  assign G387GAT = ~G176GAT | ~G302GAT;
  assign G388GAT = ~G183GAT | ~G305GAT;
  assign G389GAT = ~G190GAT | ~G305GAT;
  assign G390GAT = ~G197GAT | ~G308GAT;
  assign G391GAT = ~G204GAT | ~G308GAT;
  assign G392GAT = ~G211GAT | ~G311GAT;
  assign G393GAT = ~G218GAT | ~G311GAT;
  assign G394GAT = ~G1GAT | ~G314GAT;
  assign G395GAT = ~G29GAT | ~G314GAT;
  assign G396GAT = ~G57GAT | ~G317GAT;
  assign G397GAT = ~G85GAT | ~G317GAT;
  assign G398GAT = ~G8GAT | ~G320GAT;
  assign G399GAT = ~G36GAT | ~G320GAT;
  assign G400GAT = ~G64GAT | ~G323GAT;
  assign G401GAT = ~G92GAT | ~G323GAT;
  assign G402GAT = ~G15GAT | ~G326GAT;
  assign G403GAT = ~G43GAT | ~G326GAT;
  assign G404GAT = ~G71GAT | ~G329GAT;
  assign G405GAT = ~G99GAT | ~G329GAT;
  assign G406GAT = ~G22GAT | ~G332GAT;
  assign G407GAT = ~G50GAT | ~G332GAT;
  assign G408GAT = ~G78GAT | ~G335GAT;
  assign G409GAT = ~G106GAT | ~G335GAT;
  assign G410GAT = ~G113GAT | ~G338GAT;
  assign G411GAT = ~G141GAT | ~G338GAT;
  assign G412GAT = ~G169GAT | ~G341GAT;
  assign G413GAT = ~G197GAT | ~G341GAT;
  assign G414GAT = ~G120GAT | ~G344GAT;
  assign G415GAT = ~G148GAT | ~G344GAT;
  assign G416GAT = ~G176GAT | ~G347GAT;
  assign G417GAT = ~G204GAT | ~G347GAT;
  assign G418GAT = ~G127GAT | ~G350GAT;
  assign G419GAT = ~G155GAT | ~G350GAT;
  assign G420GAT = ~G183GAT | ~G353GAT;
  assign G421GAT = ~G211GAT | ~G353GAT;
  assign G422GAT = ~G134GAT | ~G356GAT;
  assign G423GAT = ~G162GAT | ~G356GAT;
  assign G424GAT = ~G190GAT | ~G359GAT;
  assign G425GAT = ~G218GAT | ~G359GAT;
  assign G426GAT = ~G362GAT | ~G363GAT;
  assign G429GAT = ~G364GAT | ~G365GAT;
  assign G432GAT = ~G366GAT | ~G367GAT;
  assign G435GAT = ~G368GAT | ~G369GAT;
  assign G438GAT = ~G370GAT | ~G371GAT;
  assign G441GAT = ~G372GAT | ~G373GAT;
  assign G444GAT = ~G374GAT | ~G375GAT;
  assign G447GAT = ~G376GAT | ~G377GAT;
  assign G450GAT = ~G378GAT | ~G379GAT;
  assign G453GAT = ~G380GAT | ~G381GAT;
  assign G456GAT = ~G382GAT | ~G383GAT;
  assign G459GAT = ~G384GAT | ~G385GAT;
  assign G462GAT = ~G386GAT | ~G387GAT;
  assign G465GAT = ~G388GAT | ~G389GAT;
  assign G468GAT = ~G390GAT | ~G391GAT;
  assign G471GAT = ~G392GAT | ~G393GAT;
  assign G474GAT = ~G394GAT | ~G395GAT;
  assign G477GAT = ~G396GAT | ~G397GAT;
  assign G480GAT = ~G398GAT | ~G399GAT;
  assign G483GAT = ~G400GAT | ~G401GAT;
  assign G486GAT = ~G402GAT | ~G403GAT;
  assign G489GAT = ~G404GAT | ~G405GAT;
  assign G492GAT = ~G406GAT | ~G407GAT;
  assign G495GAT = ~G408GAT | ~G409GAT;
  assign G498GAT = ~G410GAT | ~G411GAT;
  assign G501GAT = ~G412GAT | ~G413GAT;
  assign G504GAT = ~G414GAT | ~G415GAT;
  assign G507GAT = ~G416GAT | ~G417GAT;
  assign G510GAT = ~G418GAT | ~G419GAT;
  assign G513GAT = ~G420GAT | ~G421GAT;
  assign G516GAT = ~G422GAT | ~G423GAT;
  assign G519GAT = ~G424GAT | ~G425GAT;
  assign G522GAT = ~G426GAT | ~G429GAT;
  assign G525GAT = ~G432GAT | ~G435GAT;
  assign G528GAT = ~G438GAT | ~G441GAT;
  assign G531GAT = ~G444GAT | ~G447GAT;
  assign G534GAT = ~G450GAT | ~G453GAT;
  assign G537GAT = ~G456GAT | ~G459GAT;
  assign G540GAT = ~G462GAT | ~G465GAT;
  assign G543GAT = ~G468GAT | ~G471GAT;
  assign G546GAT = ~G474GAT | ~G477GAT;
  assign G549GAT = ~G480GAT | ~G483GAT;
  assign G552GAT = ~G486GAT | ~G489GAT;
  assign G555GAT = ~G492GAT | ~G495GAT;
  assign G558GAT = ~G498GAT | ~G501GAT;
  assign G561GAT = ~G504GAT | ~G507GAT;
  assign G564GAT = ~G510GAT | ~G513GAT;
  assign G567GAT = ~G516GAT | ~G519GAT;
  assign G570GAT = ~G426GAT | ~G522GAT;
  assign G571GAT = ~G429GAT | ~G522GAT;
  assign G572GAT = ~G432GAT | ~G525GAT;
  assign G573GAT = ~G435GAT | ~G525GAT;
  assign G574GAT = ~G438GAT | ~G528GAT;
  assign G575GAT = ~G441GAT | ~G528GAT;
  assign G576GAT = ~G444GAT | ~G531GAT;
  assign G577GAT = ~G447GAT | ~G531GAT;
  assign G578GAT = ~G450GAT | ~G534GAT;
  assign G579GAT = ~G453GAT | ~G534GAT;
  assign G580GAT = ~G456GAT | ~G537GAT;
  assign G581GAT = ~G459GAT | ~G537GAT;
  assign G582GAT = ~G462GAT | ~G540GAT;
  assign G583GAT = ~G465GAT | ~G540GAT;
  assign G584GAT = ~G468GAT | ~G543GAT;
  assign G585GAT = ~G471GAT | ~G543GAT;
  assign G586GAT = ~G474GAT | ~G546GAT;
  assign G587GAT = ~G477GAT | ~G546GAT;
  assign G588GAT = ~G480GAT | ~G549GAT;
  assign G589GAT = ~G483GAT | ~G549GAT;
  assign G590GAT = ~G486GAT | ~G552GAT;
  assign G591GAT = ~G489GAT | ~G552GAT;
  assign G592GAT = ~G492GAT | ~G555GAT;
  assign G593GAT = ~G495GAT | ~G555GAT;
  assign G594GAT = ~G498GAT | ~G558GAT;
  assign G595GAT = ~G501GAT | ~G558GAT;
  assign G596GAT = ~G504GAT | ~G561GAT;
  assign G597GAT = ~G507GAT | ~G561GAT;
  assign G598GAT = ~G510GAT | ~G564GAT;
  assign G599GAT = ~G513GAT | ~G564GAT;
  assign G600GAT = ~G516GAT | ~G567GAT;
  assign G601GAT = ~G519GAT | ~G567GAT;
  assign G602GAT = ~G570GAT | ~G571GAT;
  assign G607GAT = ~G572GAT | ~G573GAT;
  assign G612GAT = ~G574GAT | ~G575GAT;
  assign G617GAT = ~G576GAT | ~G577GAT;
  assign G622GAT = ~G578GAT | ~G579GAT;
  assign G627GAT = ~G580GAT | ~G581GAT;
  assign G632GAT = ~G582GAT | ~G583GAT;
  assign G637GAT = ~G584GAT | ~G585GAT;
  assign G642GAT = ~G586GAT | ~G587GAT;
  assign G645GAT = ~G588GAT | ~G589GAT;
  assign G648GAT = ~G590GAT | ~G591GAT;
  assign G651GAT = ~G592GAT | ~G593GAT;
  assign G654GAT = ~G594GAT | ~G595GAT;
  assign G657GAT = ~G596GAT | ~G597GAT;
  assign G660GAT = ~G598GAT | ~G599GAT;
  assign G663GAT = ~G600GAT | ~G601GAT;
  assign G666GAT = ~G602GAT | ~G607GAT;
  assign G669GAT = ~G612GAT | ~G617GAT;
  assign G672GAT = ~G602GAT | ~G612GAT;
  assign G675GAT = ~G607GAT | ~G617GAT;
  assign G678GAT = ~G622GAT | ~G627GAT;
  assign G681GAT = ~G632GAT | ~G637GAT;
  assign G684GAT = ~G622GAT | ~G632GAT;
  assign G687GAT = ~G627GAT | ~G637GAT;
  assign G690GAT = ~G602GAT | ~G666GAT;
  assign G691GAT = ~G607GAT | ~G666GAT;
  assign G692GAT = ~G612GAT | ~G669GAT;
  assign G693GAT = ~G617GAT | ~G669GAT;
  assign G694GAT = ~G602GAT | ~G672GAT;
  assign G695GAT = ~G612GAT | ~G672GAT;
  assign G696GAT = ~G607GAT | ~G675GAT;
  assign G697GAT = ~G617GAT | ~G675GAT;
  assign G698GAT = ~G622GAT | ~G678GAT;
  assign G699GAT = ~G627GAT | ~G678GAT;
  assign G700GAT = ~G632GAT | ~G681GAT;
  assign G701GAT = ~G637GAT | ~G681GAT;
  assign G702GAT = ~G622GAT | ~G684GAT;
  assign G703GAT = ~G632GAT | ~G684GAT;
  assign G704GAT = ~G627GAT | ~G687GAT;
  assign G705GAT = ~G637GAT | ~G687GAT;
  assign G706GAT = ~G690GAT | ~G691GAT;
  assign G709GAT = ~G692GAT | ~G693GAT;
  assign G712GAT = ~G694GAT | ~G695GAT;
  assign G715GAT = ~G696GAT | ~G697GAT;
  assign G718GAT = ~G698GAT | ~G699GAT;
  assign G721GAT = ~G700GAT | ~G701GAT;
  assign G724GAT = ~G702GAT | ~G703GAT;
  assign G727GAT = ~G704GAT | ~G705GAT;
  assign G730GAT = ~G242GAT | ~G718GAT;
  assign G733GAT = ~G245GAT | ~G721GAT;
  assign G736GAT = ~G248GAT | ~G724GAT;
  assign G739GAT = ~G251GAT | ~G727GAT;
  assign G742GAT = ~G254GAT | ~G706GAT;
  assign G745GAT = ~G257GAT | ~G709GAT;
  assign G748GAT = ~G260GAT | ~G712GAT;
  assign G751GAT = ~G263GAT | ~G715GAT;
  assign G754GAT = ~G242GAT | ~G730GAT;
  assign G755GAT = ~G718GAT | ~G730GAT;
  assign G756GAT = ~G245GAT | ~G733GAT;
  assign G757GAT = ~G721GAT | ~G733GAT;
  assign G758GAT = ~G248GAT | ~G736GAT;
  assign G759GAT = ~G724GAT | ~G736GAT;
  assign G760GAT = ~G251GAT | ~G739GAT;
  assign G761GAT = ~G727GAT | ~G739GAT;
  assign G762GAT = ~G254GAT | ~G742GAT;
  assign G763GAT = ~G706GAT | ~G742GAT;
  assign G764GAT = ~G257GAT | ~G745GAT;
  assign G765GAT = ~G709GAT | ~G745GAT;
  assign G766GAT = ~G260GAT | ~G748GAT;
  assign G767GAT = ~G712GAT | ~G748GAT;
  assign G768GAT = ~G263GAT | ~G751GAT;
  assign G769GAT = ~G715GAT | ~G751GAT;
  assign G770GAT = ~G754GAT | ~G755GAT;
  assign G773GAT = ~G756GAT | ~G757GAT;
  assign G776GAT = ~G758GAT | ~G759GAT;
  assign G779GAT = ~G760GAT | ~G761GAT;
  assign G782GAT = ~G762GAT | ~G763GAT;
  assign G785GAT = ~G764GAT | ~G765GAT;
  assign G788GAT = ~G766GAT | ~G767GAT;
  assign G791GAT = ~G768GAT | ~G769GAT;
  assign G794GAT = ~G642GAT | ~G770GAT;
  assign G797GAT = ~G645GAT | ~G773GAT;
  assign G800GAT = ~G648GAT | ~G776GAT;
  assign G803GAT = ~G651GAT | ~G779GAT;
  assign G806GAT = ~G654GAT | ~G782GAT;
  assign G809GAT = ~G657GAT | ~G785GAT;
  assign G812GAT = ~G660GAT | ~G788GAT;
  assign G815GAT = ~G663GAT | ~G791GAT;
  assign G818GAT = ~G642GAT | ~G794GAT;
  assign G819GAT = ~G770GAT | ~G794GAT;
  assign G820GAT = ~G645GAT | ~G797GAT;
  assign G821GAT = ~G773GAT | ~G797GAT;
  assign G822GAT = ~G648GAT | ~G800GAT;
  assign G823GAT = ~G776GAT | ~G800GAT;
  assign G824GAT = ~G651GAT | ~G803GAT;
  assign G825GAT = ~G779GAT | ~G803GAT;
  assign G826GAT = ~G654GAT | ~G806GAT;
  assign G827GAT = ~G782GAT | ~G806GAT;
  assign G828GAT = ~G657GAT | ~G809GAT;
  assign G829GAT = ~G785GAT | ~G809GAT;
  assign G830GAT = ~G660GAT | ~G812GAT;
  assign G831GAT = ~G788GAT | ~G812GAT;
  assign G832GAT = ~G663GAT | ~G815GAT;
  assign G833GAT = ~G791GAT | ~G815GAT;
  assign G834GAT = ~G818GAT | ~G819GAT;
  assign G847GAT = ~G820GAT | ~G821GAT;
  assign G860GAT = ~G822GAT | ~G823GAT;
  assign G873GAT = ~G824GAT | ~G825GAT;
  assign G886GAT = ~G828GAT | ~G829GAT;
  assign G899GAT = ~G832GAT | ~G833GAT;
  assign G912GAT = ~G830GAT | ~G831GAT;
  assign G925GAT = ~G826GAT | ~G827GAT;
  assign G938GAT = ~G834GAT;
  assign G939GAT = ~G847GAT;
  assign G940GAT = ~G860GAT;
  assign G941GAT = ~G834GAT;
  assign G942GAT = ~G847GAT;
  assign G943GAT = ~G873GAT;
  assign G944GAT = ~G834GAT;
  assign G945GAT = ~G860GAT;
  assign G946GAT = ~G873GAT;
  assign G947GAT = ~G847GAT;
  assign G948GAT = ~G860GAT;
  assign G949GAT = ~G873GAT;
  assign G950GAT = ~G886GAT;
  assign G951GAT = ~G899GAT;
  assign G952GAT = ~G886GAT;
  assign G953GAT = ~G912GAT;
  assign G954GAT = ~G925GAT;
  assign G955GAT = ~G899GAT;
  assign G956GAT = ~G925GAT;
  assign G957GAT = ~G912GAT;
  assign G958GAT = ~G925GAT;
  assign G959GAT = ~G886GAT;
  assign G960GAT = ~G912GAT;
  assign G961GAT = ~G925GAT;
  assign G962GAT = ~G886GAT;
  assign G963GAT = ~G899GAT;
  assign G964GAT = ~G925GAT;
  assign G965GAT = ~G912GAT;
  assign G966GAT = ~G899GAT;
  assign G967GAT = ~G886GAT;
  assign G968GAT = ~G912GAT;
  assign G969GAT = ~G899GAT;
  assign G970GAT = ~G847GAT;
  assign G971GAT = ~G873GAT;
  assign G972GAT = ~G847GAT;
  assign G973GAT = ~G860GAT;
  assign G974GAT = ~G834GAT;
  assign G975GAT = ~G873GAT;
  assign G976GAT = ~G834GAT;
  assign G977GAT = ~G860GAT;
  assign G978GAT = G873GAT & G940GAT & G938GAT & G939GAT;
  assign G979GAT = G943GAT & G860GAT & G941GAT & G942GAT;
  assign G980GAT = G946GAT & G945GAT & G944GAT & G847GAT;
  assign G981GAT = G949GAT & G948GAT & G834GAT & G947GAT;
  assign G982GAT = G899GAT & G960GAT & G958GAT & G959GAT;
  assign G983GAT = G963GAT & G912GAT & G961GAT & G962GAT;
  assign G984GAT = G966GAT & G965GAT & G964GAT & G886GAT;
  assign G985GAT = G969GAT & G968GAT & G925GAT & G967GAT;
  assign G986GAT = G981GAT | G980GAT | G978GAT | G979GAT;
  assign G991GAT = G985GAT | G984GAT | G982GAT | G983GAT;
  assign G996GAT = G986GAT & G951GAT & G912GAT & G925GAT & G950GAT;
  assign G1001GAT = G986GAT & G899GAT & G953GAT & G925GAT & G952GAT;
  assign G1006GAT = G986GAT & G955GAT & G912GAT & G954GAT & G886GAT;
  assign G1011GAT = G986GAT & G899GAT & G957GAT & G956GAT & G886GAT;
  assign G1016GAT = G991GAT & G971GAT & G860GAT & G834GAT & G970GAT;
  assign G1021GAT = G991GAT & G873GAT & G973GAT & G834GAT & G972GAT;
  assign G1026GAT = G991GAT & G975GAT & G860GAT & G974GAT & G847GAT;
  assign G1031GAT = G991GAT & G873GAT & G977GAT & G976GAT & G847GAT;
  assign G1036GAT = G834GAT & G996GAT;
  assign G1039GAT = G847GAT & G996GAT;
  assign G1042GAT = G860GAT & G996GAT;
  assign G1045GAT = G873GAT & G996GAT;
  assign G1048GAT = G834GAT & G1001GAT;
  assign G1051GAT = G847GAT & G1001GAT;
  assign G1054GAT = G860GAT & G1001GAT;
  assign G1057GAT = G873GAT & G1001GAT;
  assign G1060GAT = G834GAT & G1006GAT;
  assign G1063GAT = G847GAT & G1006GAT;
  assign G1066GAT = G860GAT & G1006GAT;
  assign G1069GAT = G873GAT & G1006GAT;
  assign G1072GAT = G834GAT & G1011GAT;
  assign G1075GAT = G847GAT & G1011GAT;
  assign G1078GAT = G860GAT & G1011GAT;
  assign G1081GAT = G873GAT & G1011GAT;
  assign G1084GAT = G925GAT & G1016GAT;
  assign G1087GAT = G886GAT & G1016GAT;
  assign G1090GAT = G912GAT & G1016GAT;
  assign G1093GAT = G899GAT & G1016GAT;
  assign G1096GAT = G925GAT & G1021GAT;
  assign G1099GAT = G886GAT & G1021GAT;
  assign G1102GAT = G912GAT & G1021GAT;
  assign G1105GAT = G899GAT & G1021GAT;
  assign G1108GAT = G925GAT & G1026GAT;
  assign G1111GAT = G886GAT & G1026GAT;
  assign G1114GAT = G912GAT & G1026GAT;
  assign G1117GAT = G899GAT & G1026GAT;
  assign G1120GAT = G925GAT & G1031GAT;
  assign G1123GAT = G886GAT & G1031GAT;
  assign G1126GAT = G912GAT & G1031GAT;
  assign G1129GAT = G899GAT & G1031GAT;
  assign G1132GAT = ~G1GAT | ~G1036GAT;
  assign G1135GAT = ~G8GAT | ~G1039GAT;
  assign G1138GAT = ~G15GAT | ~G1042GAT;
  assign G1141GAT = ~G22GAT | ~G1045GAT;
  assign G1144GAT = ~G29GAT | ~G1048GAT;
  assign G1147GAT = ~G36GAT | ~G1051GAT;
  assign G1150GAT = ~G43GAT | ~G1054GAT;
  assign G1153GAT = ~G50GAT | ~G1057GAT;
  assign G1156GAT = ~G57GAT | ~G1060GAT;
  assign G1159GAT = ~G64GAT | ~G1063GAT;
  assign G1162GAT = ~G71GAT | ~G1066GAT;
  assign G1165GAT = ~G78GAT | ~G1069GAT;
  assign G1168GAT = ~G85GAT | ~G1072GAT;
  assign G1171GAT = ~G92GAT | ~G1075GAT;
  assign G1174GAT = ~G99GAT | ~G1078GAT;
  assign G1177GAT = ~G106GAT | ~G1081GAT;
  assign G1180GAT = ~G113GAT | ~G1084GAT;
  assign G1183GAT = ~G120GAT | ~G1087GAT;
  assign G1186GAT = ~G127GAT | ~G1090GAT;
  assign G1189GAT = ~G134GAT | ~G1093GAT;
  assign G1192GAT = ~G141GAT | ~G1096GAT;
  assign G1195GAT = ~G148GAT | ~G1099GAT;
  assign G1198GAT = ~G155GAT | ~G1102GAT;
  assign G1201GAT = ~G162GAT | ~G1105GAT;
  assign G1204GAT = ~G169GAT | ~G1108GAT;
  assign G1207GAT = ~G176GAT | ~G1111GAT;
  assign G1210GAT = ~G183GAT | ~G1114GAT;
  assign G1213GAT = ~G190GAT | ~G1117GAT;
  assign G1216GAT = ~G197GAT | ~G1120GAT;
  assign G1219GAT = ~G204GAT | ~G1123GAT;
  assign G1222GAT = ~G211GAT | ~G1126GAT;
  assign G1225GAT = ~G218GAT | ~G1129GAT;
  assign G1228GAT = ~G1GAT | ~G1132GAT;
  assign G1229GAT = ~G1036GAT | ~G1132GAT;
  assign G1230GAT = ~G8GAT | ~G1135GAT;
  assign G1231GAT = ~G1039GAT | ~G1135GAT;
  assign G1232GAT = ~G15GAT | ~G1138GAT;
  assign G1233GAT = ~G1042GAT | ~G1138GAT;
  assign G1234GAT = ~G22GAT | ~G1141GAT;
  assign G1235GAT = ~G1045GAT | ~G1141GAT;
  assign G1236GAT = ~G29GAT | ~G1144GAT;
  assign G1237GAT = ~G1048GAT | ~G1144GAT;
  assign G1238GAT = ~G36GAT | ~G1147GAT;
  assign G1239GAT = ~G1051GAT | ~G1147GAT;
  assign G1240GAT = ~G43GAT | ~G1150GAT;
  assign G1241GAT = ~G1054GAT | ~G1150GAT;
  assign G1242GAT = ~G50GAT | ~G1153GAT;
  assign G1243GAT = ~G1057GAT | ~G1153GAT;
  assign G1244GAT = ~G57GAT | ~G1156GAT;
  assign G1245GAT = ~G1060GAT | ~G1156GAT;
  assign G1246GAT = ~G64GAT | ~G1159GAT;
  assign G1247GAT = ~G1063GAT | ~G1159GAT;
  assign G1248GAT = ~G71GAT | ~G1162GAT;
  assign G1249GAT = ~G1066GAT | ~G1162GAT;
  assign G1250GAT = ~G78GAT | ~G1165GAT;
  assign G1251GAT = ~G1069GAT | ~G1165GAT;
  assign G1252GAT = ~G85GAT | ~G1168GAT;
  assign G1253GAT = ~G1072GAT | ~G1168GAT;
  assign G1254GAT = ~G92GAT | ~G1171GAT;
  assign G1255GAT = ~G1075GAT | ~G1171GAT;
  assign G1256GAT = ~G99GAT | ~G1174GAT;
  assign G1257GAT = ~G1078GAT | ~G1174GAT;
  assign G1258GAT = ~G106GAT | ~G1177GAT;
  assign G1259GAT = ~G1081GAT | ~G1177GAT;
  assign G1260GAT = ~G113GAT | ~G1180GAT;
  assign G1261GAT = ~G1084GAT | ~G1180GAT;
  assign G1262GAT = ~G120GAT | ~G1183GAT;
  assign G1263GAT = ~G1087GAT | ~G1183GAT;
  assign G1264GAT = ~G127GAT | ~G1186GAT;
  assign G1265GAT = ~G1090GAT | ~G1186GAT;
  assign G1266GAT = ~G134GAT | ~G1189GAT;
  assign G1267GAT = ~G1093GAT | ~G1189GAT;
  assign G1268GAT = ~G141GAT | ~G1192GAT;
  assign G1269GAT = ~G1096GAT | ~G1192GAT;
  assign G1270GAT = ~G148GAT | ~G1195GAT;
  assign G1271GAT = ~G1099GAT | ~G1195GAT;
  assign G1272GAT = ~G155GAT | ~G1198GAT;
  assign G1273GAT = ~G1102GAT | ~G1198GAT;
  assign G1274GAT = ~G162GAT | ~G1201GAT;
  assign G1275GAT = ~G1105GAT | ~G1201GAT;
  assign G1276GAT = ~G169GAT | ~G1204GAT;
  assign G1277GAT = ~G1108GAT | ~G1204GAT;
  assign G1278GAT = ~G176GAT | ~G1207GAT;
  assign G1279GAT = ~G1111GAT | ~G1207GAT;
  assign G1280GAT = ~G183GAT | ~G1210GAT;
  assign G1281GAT = ~G1114GAT | ~G1210GAT;
  assign G1282GAT = ~G190GAT | ~G1213GAT;
  assign G1283GAT = ~G1117GAT | ~G1213GAT;
  assign G1284GAT = ~G197GAT | ~G1216GAT;
  assign G1285GAT = ~G1120GAT | ~G1216GAT;
  assign G1286GAT = ~G204GAT | ~G1219GAT;
  assign G1287GAT = ~G1123GAT | ~G1219GAT;
  assign G1288GAT = ~G211GAT | ~G1222GAT;
  assign G1289GAT = ~G1126GAT | ~G1222GAT;
  assign G1290GAT = ~G218GAT | ~G1225GAT;
  assign G1291GAT = ~G1129GAT | ~G1225GAT;
  assign G1292GAT = ~G1228GAT | ~G1229GAT;
  assign G1293GAT = ~G1230GAT | ~G1231GAT;
  assign G1294GAT = ~G1232GAT | ~G1233GAT;
  assign G1295GAT = ~G1234GAT | ~G1235GAT;
  assign G1296GAT = ~G1236GAT | ~G1237GAT;
  assign G1297GAT = ~G1238GAT | ~G1239GAT;
  assign G1298GAT = ~G1240GAT | ~G1241GAT;
  assign G1299GAT = ~G1242GAT | ~G1243GAT;
  assign G1300GAT = ~G1244GAT | ~G1245GAT;
  assign G1301GAT = ~G1246GAT | ~G1247GAT;
  assign G1302GAT = ~G1248GAT | ~G1249GAT;
  assign G1303GAT = ~G1250GAT | ~G1251GAT;
  assign G1304GAT = ~G1252GAT | ~G1253GAT;
  assign G1305GAT = ~G1254GAT | ~G1255GAT;
  assign G1306GAT = ~G1256GAT | ~G1257GAT;
  assign G1307GAT = ~G1258GAT | ~G1259GAT;
  assign G1308GAT = ~G1260GAT | ~G1261GAT;
  assign G1309GAT = ~G1262GAT | ~G1263GAT;
  assign G1310GAT = ~G1264GAT | ~G1265GAT;
  assign G1311GAT = ~G1266GAT | ~G1267GAT;
  assign G1312GAT = ~G1268GAT | ~G1269GAT;
  assign G1313GAT = ~G1270GAT | ~G1271GAT;
  assign G1314GAT = ~G1272GAT | ~G1273GAT;
  assign G1315GAT = ~G1274GAT | ~G1275GAT;
  assign G1316GAT = ~G1276GAT | ~G1277GAT;
  assign G1317GAT = ~G1278GAT | ~G1279GAT;
  assign G1318GAT = ~G1280GAT | ~G1281GAT;
  assign G1319GAT = ~G1282GAT | ~G1283GAT;
  assign G1320GAT = ~G1284GAT | ~G1285GAT;
  assign G1321GAT = ~G1286GAT | ~G1287GAT;
  assign G1322GAT = ~G1288GAT | ~G1289GAT;
  assign G1323GAT = ~G1290GAT | ~G1291GAT;
  assign G1324GAT = G1292GAT;
  assign G1325GAT = G1293GAT;
  assign G1326GAT = G1294GAT;
  assign G1327GAT = G1295GAT;
  assign G1328GAT = G1296GAT;
  assign G1329GAT = G1297GAT;
  assign G1330GAT = G1298GAT;
  assign G1331GAT = G1299GAT;
  assign G1332GAT = G1300GAT;
  assign G1333GAT = G1301GAT;
  assign G1334GAT = G1302GAT;
  assign G1335GAT = G1303GAT;
  assign G1336GAT = G1304GAT;
  assign G1337GAT = G1305GAT;
  assign G1338GAT = G1306GAT;
  assign G1339GAT = G1307GAT;
  assign G1340GAT = G1308GAT;
  assign G1341GAT = G1309GAT;
  assign G1342GAT = G1310GAT;
  assign G1343GAT = G1311GAT;
  assign G1344GAT = G1312GAT;
  assign G1345GAT = G1313GAT;
  assign G1346GAT = G1314GAT;
  assign G1347GAT = G1315GAT;
  assign G1348GAT = G1316GAT;
  assign G1349GAT = G1317GAT;
  assign G1350GAT = G1318GAT;
  assign G1351GAT = G1319GAT;
  assign G1352GAT = G1320GAT;
  assign G1353GAT = G1321GAT;
  assign G1354GAT = G1322GAT;
  assign G1355GAT = G1323GAT;
endmodule


