// Benchmark "b22_C_lock" written by ABC on Thu May 13 23:43:20 2021

module b22_C_lock ( 
    SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_,
    SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_,
    SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_,
    SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P1_ADDR_REG_19__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_RD_REG_SCAN_IN,
    P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN,
    P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN,
    P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN,
    P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN,
    P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN,
    P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN,
    P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN,
    P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN,
    P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN,
    P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN,
    P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
    P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
    P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
    P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
    P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
    P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
    P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
    P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
    P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
    P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
    P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
    P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
    P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
    P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
    P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
    P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
    P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
    P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
    P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
    P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
    P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
    P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
    P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
    P3_ADDR_REG_19__SCAN_IN,
    P2_U3328  );
  input  SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_,
    SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_,
    SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_,
    SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P1_ADDR_REG_19__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_RD_REG_SCAN_IN,
    P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN,
    P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN,
    P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN,
    P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN,
    P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN,
    P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN,
    P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN,
    P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN,
    P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN,
    P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN,
    P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
    P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
    P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
    P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
    P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
    P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
    P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
    P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
    P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
    P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
    P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
    P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
    P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
    P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
    P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
    P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
    P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
    P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
    P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
    P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
    P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
    P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
    P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
    P3_ADDR_REG_19__SCAN_IN;
  output P2_U3328;
  wire n13293, n13257, n11682, n16904, n21822, n11667, n11671, n22473,
    n22268, n22115, n22334, n22135, n21536, n21716, n12577, n12713, n12732,
    n19373, n12329, n19100, n18880, n18900, n18756, n12841, n15740, n13114,
    n11677, n11680, n22834, n12636, n12789, n13493, n12609, n13037, n18814,
    n13579, n12406, n12418, n11931, n17888, n17889, n12818, n12892, n12090,
    n12945, n13394, n13400, n12870, n12553, n12007, n11987, n12009, n22812,
    n15966, n12417, n12122, n12559, n12544, n12542, n11916, n11966, n12536,
    n13476, n12338, n12879, n12014, n15777, n12310, n13401, n12334, n12471,
    n13482, n19083, n12849, n15739, n16128, n16039, n15940, n15943, n21950,
    n20068, n19357, n19193, n18739, n12006, n11980, n12407, n12539, n12538,
    n12535, n11971, n11970, n11985, n12985, n12525, n12522, n16712, n13337,
    n13477, n11964, n22813, n22401, n21198, n22913, n12169, n12170, n12171,
    n11994, n11923, n13069, n12327, n13007, n11990, n12847, n12340, n12341,
    n13334, n13270, n13191, n11915, n11983, n11998, n11999, n12000, n12001,
    n13091, n12011, n12309, n13407, n13357, n12845, n16129, n15704, n19346,
    n11973, n11974, n11975, n12331, n12332, n13405, n15968, n15748, n16158,
    n22389, n21034, n19201, n12696, n12734, n12328, n13071, n12552, n12548,
    n12547, n12961, n12405, n12796, n12322, n12530, n12529, n12336, n12335,
    n12337, n20545, n12901, n12897, n21794, n11992, n19333, n19167, n12839,
    n15689, n15691, n16716, n16160, n16041, n15955, n22243, n21964, n21815,
    n21031, n20886, n20409, n12830, n12825, n19696, n12669, n12639, n12642,
    n11936, n13123, n12330, n13009, n12988, n12958, n12943, n12914, n12915,
    n11917, n11932, n12846, n13319, n11969, n11968, n12307, n12308, n11993,
    n12804, n12526, n12802, n12828, n14417, n19213, n22901, n20243, n20081,
    n13152, n13006, n23453, n22863, n11977, n11979, n22784, n13362, n22765,
    n22739, n22645, n13299, n22559, n12694, n11982, n12002, n18818, n11691,
    n11693, n11697, n11698, n11935, n12899, n12883, n11701, n16189, n11929,
    n13159, n21696, n11706, n12608, n15785, n11716, n16185, n11733, n13434,
    n11736, n12706, n19909, n11755, n11756, n15971, n11758, n11759, n11763,
    n11768, n11769, n11842, n11774, n11779, n11780, n12811, n11788, n11984,
    n12916, n12123, n11933, n11793, n11795, n12600, n11799, n11801, n11802,
    n11803, n11981, n11807, n11809, n11810, n11814, n11815, n11817, n11819,
    n12339, n11827, n11830, n16909, n11934, n15125, n12584, n11918, n11976,
    n11922, n11924, n12569, n11928, n12316, n12891, n16826, n11937, n12416,
    n12628, n11965, n19277, n11967, n11972, n12621, n11978, n11986, n12987,
    n12944, n11988, n11989, n11991, n12003, n13487, n12801, n12904, n11995,
    n11996, n11997, P2_U3328_Lock, n12976, n12004, n12005, n12008, n12010,
    n13209, n12012, n12013, n12015, n12016, n13317, n12017, n12018, n13119,
    n12019, n12020, n13118, n12021, n12022, n12922, n12965, n12995, n12641,
    n12637, n12304, n12659, n12305, n12306, n13389, n12312, n12314, n12311,
    n12313, n12755, n12315, n12317, n12318, n12319, n12320, n12321, n13256,
    n12323, n12324, n12325, n13035, n12326, n12561, n12333, n12960, n13554,
    n13380, n12842, n16954, n12419, n12458, n12886, n12470, n12984, n13141,
    n13484, n12554, n12528, n19889, n12517, n12556, n12602, n12520, n12898,
    n12826, n12473, n12472, n13378, n13377, n12475, n12474, n12476, n12599,
    n13363, n12478, n12477, n12596, n13333, n12480, n12479, n12481, n12595,
    n13318, n12483, n12482, n12484, n13298, n12486, n12485, n12487, n12593,
    n13269, n12489, n12488, n12490, n12592, n13255, n12492, n12491, n12493,
    n12587, n13215, n12495, n12494, n12496, n12585, n15172, n13190, n12498,
    n12497, n12499, n12579, n12674, n12501, n12500, n12576, n12578, n12503,
    n12502, n12504, n13124, n12506, n12505, n12571, n12508, n12507, n12568,
    n12570, n12510, n12509, n12567, n12512, n12511, n12566, n12514, n12513,
    n12563, n12565, n12516, n12515, n12562, n13036, n12519, n12518, n12521,
    n13553, n12524, n12523, n12527, n13599, n12531, n12533, n12532, n12534,
    n12537, n13649, n12540, n12541, n12543, n12545, n12546, n13706, n12549,
    n12551, n12550, n12555, n12558, n12557, n12560, n13068, n12564, n13093,
    n13092, n12754, n12731, n12712, n12573, n12572, n12574, n12693, n12575,
    n13151, n12581, n12580, n12582, n12658, n12583, n13216, n12586, n13236,
    n12589, n12588, n12590, n13235, n12591, n12594, n12598, n12597, n12601,
    n12990, n12603, n13095, n12715, n12604, n12605, n13126, n12624, n12606,
    n12626, n12607, n13483, n12610, n12611, n12612, n12613, n12615, n12614,
    n12617, n12616, n12618, n12619, n12620, n12622, n12623, n13127, n12625,
    n12634, n12627, n12629, n12631, n12630, n12632, n12633, n15126, n12635,
    n21658, n15113, n12638, n22929, n12640, n22774, n12645, n12643, n12644,
    n12647, n12860, n12646, n16899, n22820, n12649, n21976, n15118, n12648,
    n12655, n12652, n12650, n12651, n12654, n12653, n16895, n16194, n12656,
    n12657, n21872, n12662, n12660, n12661, n12665, n12663, n12664, n12668,
    n12666, n12667, n12671, n12908, n12938, n17015, n12950, n12977, n17049,
    n13019, n13048, n17266, n13076, n13103, n17095, n12763, n12742, n17228,
    n12725, n12704, n17103, n13138, n13165, n17143, n12685, n13200, n21811,
    n12670, n21939, n13416, n13187, n13395, n12673, n15787, n12672, n21661,
    n12679, n12675, n12677, n12676, n12678, n12690, n12681, n12680, n12684,
    n12682, n12683, n12688, n21706, n12686, n12687, n21788, n21496, n12869,
    n12689, n13183, n12692, n12691, n13182, n13181, n21168, n12701, n12695,
    n12699, n12697, n17155, n17120, n12698, n12700, n12703, n12702, n12711,
    n21211, n12705, n12709, n12707, n12708, n12710, n21364, n13421, n21003,
    n14656, n12722, n12714, n12720, n12716, n12717, n12718, n17210, n17131,
    n12719, n12721, n12724, n12723, n12730, n21044, n12728, n12726, n12727,
    n12729, n21192, n13419, n13121, n15778, n20842, n14637, n12741, n12733,
    n12739, n12757, n12735, n12736, n12737, n17229, n12738, n12740, n20861,
    n12744, n12743, n12749, n12747, n12745, n12746, n12748, n21025, n12751,
    n12750, n12778, n12753, n13418, n12752, n12774, n20677, n14617, n12762,
    n12756, n12760, n17238, n12758, n12759, n12761, n20724, n12772, n20721,
    n12765, n12764, n12770, n12768, n12766, n12767, n12769, n20874, n12771,
    n12775, n20524, n15716, n12773, n12786, n12776, n12781, n12777, n12785,
    n12780, n12779, n12783, n20708, n12782, n12784, n13120, n12788, n12787,
    n12794, n12792, n12790, n12791, n12793, n12808, n12795, n12798, n12797,
    n12799, n12800, n12806, n12803, n18972, n12805, n12807, n12853, n12809,
    n12832, n19078, n12810, n12813, n12812, n12817, n12815, n12814, n12816,
    n12824, n12819, n12822, n12866, n12820, n12821, n12823, n16935, n12827,
    n18819, n12829, n12831, n12834, n12833, n12840, n12835, n12838, n12836,
    n12837, n12851, n16978, n12843, n12844, n13271, n19056, n12848, n12850,
    n12881, n12852, n12854, n12856, n12871, n12855, n19187, n12857, n12859,
    n12858, n12865, n12863, n12861, n12862, n12864, n12868, n18684, n12867,
    n18735, n18671, n12873, n15750, n12872, n12878, n18730, n18667, n12877,
    n12874, n12875, n12876, n12880, n12902, n12885, n12882, n12884, n12890,
    n19210, n12888, n12887, n12889, n12894, n12893, n12895, n19225, n12896,
    n14458, n12900, n12930, n19351, n12903, n12927, n12906, n12905, n12913,
    n12907, n19370, n12911, n12909, n12910, n12912, n19567, n19438, n14478,
    n12924, n12917, n12919, n12918, n12920, n17022, n16996, n12921, n12923,
    n15755, n12925, n12926, n12929, n12928, n15757, n12933, n12931, n12932,
    n12935, n12934, n12937, n12936, n12942, n19593, n12940, n19590, n12939,
    n12941, n15701, n19547, n12949, n12946, n17021, n12947, n12948, n19575,
    n15760, n19589, n19670, n15759, n19572, n19691, n12952, n12951, n12957,
    n12955, n12953, n12954, n12956, n19886, n19556, n12959, n19756, n12967,
    n12962, n12963, n17063, n17037, n12964, n12966, n12968, n15762, n13433,
    n12969, n12970, n12971, n12972, n12973, n12974, n12975, n13005, n19913,
    n12979, n12978, n12983, n12981, n19910, n12980, n12982, n20059, n12999,
    n12998, n12986, n19864, n12997, n12989, n12992, n12991, n12993, n19865,
    n12994, n12996, n19897, n13003, n13004, n13000, n13001, n13002, n13032,
    n13030, n20035, n14539, n13018, n13008, n13016, n13010, n13013, n13011,
    n13012, n13014, n17288, n17086, n13015, n13017, n13028, n20078, n13021,
    n13020, n13026, n13024, n13022, n13023, n13025, n20221, n13027, n13034,
    n19870, n15707, n13029, n13031, n13065, n13033, n13062, n13056, n20196,
    n14558, n13045, n13043, n13038, n13040, n13039, n13041, n17267, n17089,
    n13042, n13044, n13055, n13047, n13046, n13053, n20240, n13051, n13049,
    n13050, n13052, n20382, n13054, n13061, n13060, n20227, n13058, n13057,
    n13059, n13067, n13063, n13064, n13066, n13087, n20360, n14578, n13075,
    n13070, n13073, n13096, n17256, n17082, n13072, n13074, n13085, n20405,
    n13078, n13077, n13083, n13081, n13079, n13080, n13082, n20537, n13084,
    n13088, n15711, n13086, n13089, n13436, n13090, n20519, n14601, n13102,
    n13094, n13100, n13097, n13098, n17105, n13099, n13101, n20561, n13111,
    n20558, n13105, n13104, n13110, n13108, n13106, n13107, n13109, n20702,
    n15773, n13112, n13115, n13113, n13116, n13117, n13144, n13122, n15779,
    n21332, n14695, n13132, n13125, n13130, n13153, n13128, n17196, n17154,
    n13129, n13131, n21358, n13135, n13133, n13134, n13137, n13136, n13140,
    n21352, n13139, n21514, n13169, n13142, n13150, n13143, n13146, n13145,
    n13147, n15781, n13148, n13149, n13174, n21491, n14345, n13158, n13154,
    n17160, n13156, n13155, n13157, n13161, n13160, n13164, n13162, n13163,
    n13167, n21533, n13166, n21686, n15783, n13168, n13172, n13175, n13170,
    n13171, n13173, n13179, n13177, n13176, n13178, n13180, n13185, n13184,
    n13186, n13189, n13188, n22033, n13194, n13192, n13193, n13204, n13197,
    n13195, n13196, n13199, n13198, n13202, n13220, n21961, n13201, n22108,
    n13203, n13210, n13208, n13206, n13205, n13207, n13214, n13212, n13211,
    n13213, n13229, n22204, n13219, n13217, n13218, n13240, n22132, n13227,
    n13223, n13221, n13222, n13225, n13224, n13226, n22255, n13228, n15792,
    n15732, n22122, n13234, n13231, n13230, n13232, n13233, n13249, n13239,
    n13237, n13238, n13261, n22239, n13247, n13243, n13241, n13242, n13245,
    n13244, n13246, n22381, n13248, n15795, n15736, n15794, n13254, n13251,
    n13250, n13252, n13253, n13285, n13260, n13258, n13259, n13276, n22374,
    n13268, n13264, n13262, n13263, n13266, n13265, n13267, n22256, n13274,
    n13272, n13273, n13275, n13303, n15843, n13282, n13278, n15805, n13277,
    n13280, n13279, n13281, n22382, n13283, n15942, n13284, n13291, n15354,
    n13287, n15844, n13286, n13289, n13288, n13290, n13292, n13295, n13294,
    n13296, n13297, n13302, n13300, n13301, n13324, n16042, n13310, n13306,
    n13304, n13305, n13308, n13307, n13309, n16883, n13312, n16161, n13462,
    n13311, n13313, n13315, n13314, n13316, n13332, n13322, n13320, n13321,
    n13323, n13338, n16162, n13331, n13327, n13325, n13326, n13329, n13328,
    n13330, n16886, n13354, n13335, n13336, n13367, n16718, n13339, n13345,
    n13341, n13340, n13343, n16125, n13342, n13344, n16889, n13347, n16192,
    n13355, n13346, n13352, n13349, n16118, n13348, n13350, n13351, n13353,
    n13361, n13356, n13359, n16187, n13358, n13360, n13376, n13366, n13364,
    n13365, n16178, n13368, n13375, n13370, n13369, n13373, n13371, n13372,
    n13374, n16892, n13390, n13379, n13385, n13382, n13381, n13383, n13384,
    n13388, n13386, n13387, n13393, n13391, n13392, n13404, n13398, n13396,
    n13397, n13402, n16268, n16717, n13399, n13403, n13406, n13410, n13408,
    n13409, n13411, n13471, n13413, n13412, n13469, n13414, n13415, n15790,
    n22118, n13417, n15730, n21797, n15776, n13420, n13422, n15752, n13423,
    n19087, n13425, n15753, n13424, n19196, n19091, n13426, n13427, n19360,
    n13429, n13428, n13431, n15766, n13430, n20230, n13443, n20045, n15705,
    n13432, n19678, n13435, n13439, n20391, n18728, n13437, n15120, n13438,
    n13441, n13440, n15765, n13442, n13446, n13444, n15775, n20712, n20549,
    n13445, n13447, n13448, n13449, n13451, n13450, n13455, n21376, n13452,
    n21171, n15725, n21361, n21664, n13453, n15727, n21523, n13454, n13456,
    n13457, n13458, n13460, n13459, n13461, n13464, n13463, n13466, n15974,
    n13465, n13467, n13468, n13470, n13472, n15143, n13473, n13474, n13475,
    n13481, n22148, n13479, n13478, n13480, n13485, n13486, n13496, n14988,
    n22925, n22281, n13491, n13490, n13488, n13489, n22514, n22415, n13494,
    n13492, n22642, n15077, n13495, n14989, n15150, n15818, n16825, n15142,
    n13497, n15159, n15158, n13500, n13498, n13499, n20195, n21490, n15131,
    keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
    keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
    keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
    keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
    keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
    keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
    keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
    keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
    keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
    keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
    keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
    keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
    keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
    keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
    keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
    keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
    keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
    keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
    keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
    keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
    keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
    keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
    keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
    keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
    keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
    keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
    keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
    keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
    keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
    keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
    keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
    keyinput_156, keyinput_157, keyinput_158, keyinput_159, input_0,
    input_1, AND_1, input_2, AND_2, input_3, AND_3, input_4, OR_4, input_5,
    OR_5, input_6, AND_6, input_7, AND_7, input_8, AND_8, input_9, OR_9,
    input_10, OR_10, input_11, AND_11, input_12, OR_12, input_13, OR_13,
    input_14, AND_14, input_15, OR_15, input_16, OR_16, input_17, OR_17,
    input_18, OR_18, input_19, AND_19, input_20, AND_20, input_21, AND_21,
    input_22, OR_22, input_23, OR_23, input_24, AND_24, input_25, OR_25,
    input_26, OR_26, input_27, AND_27, input_28, OR_28, input_29, OR_29,
    input_30, OR_30, input_31, AND_31, input_32, OR_32, input_33, OR_33,
    input_34, AND_34, input_35, AND_35, input_36, AND_36, input_37, OR_37,
    input_38, AND_38, input_39, OR_39, input_40, OR_40, input_41, AND_41,
    input_42, OR_42, input_43, OR_43, input_44, AND_44, input_45, OR_45,
    input_46, OR_46, input_47, AND_47, input_48, OR_48, input_49, AND_49,
    input_50, OR_50, input_51, OR_51, input_52, AND_52, input_53, OR_53,
    input_54, OR_54, input_55, OR_55, input_56, AND_56, input_57, AND_57,
    input_58, OR_58, input_59, AND_59, input_60, AND_60, input_61, OR_61,
    input_62, AND_62, input_63, OR_63, input_64, AND_64, input_65, OR_65,
    input_66, OR_66, input_67, AND_67, input_68, OR_68, input_69, AND_69,
    input_70, AND_70, input_71, AND_71, input_72, OR_72, input_73, AND_73,
    input_74, OR_74, input_75, OR_75, input_76, AND_76, input_77, AND_77,
    input_78, AND_78, input_79, OR_79, input_80, input_81, AND_81,
    input_82, AND_82, input_83, AND_83, input_84, OR_84, input_85, OR_85,
    input_86, AND_86, input_87, AND_87, input_88, AND_88, input_89, OR_89,
    input_90, OR_90, input_91, AND_91, input_92, OR_92, input_93, OR_93,
    input_94, AND_94, input_95, OR_95, input_96, OR_96, input_97, OR_97,
    input_98, OR_98, input_99, AND_99, input_100, AND_100, input_101,
    AND_101, input_102, OR_102, input_103, OR_103, input_104, AND_104,
    input_105, OR_105, input_106, OR_106, input_107, AND_107, input_108,
    OR_108, input_109, OR_109, input_110, OR_110, input_111, AND_111,
    input_112, OR_112, input_113, OR_113, input_114, AND_114, input_115,
    AND_115, input_116, AND_116, input_117, OR_117, input_118, AND_118,
    input_119, OR_119, input_120, OR_120, input_121, AND_121, input_122,
    OR_122, input_123, OR_123, input_124, AND_124, input_125, OR_125,
    input_126, OR_126, input_127, AND_127, input_128, OR_128, input_129,
    AND_129, input_130, OR_130, input_131, OR_131, input_132, AND_132,
    input_133, OR_133, input_134, OR_134, input_135, OR_135, input_136,
    AND_136, input_137, AND_137, input_138, OR_138, input_139, AND_139,
    input_140, AND_140, input_141, OR_141, input_142, AND_142, input_143,
    OR_143, input_144, AND_144, input_145, OR_145, input_146, OR_146,
    input_147, AND_147, input_148, OR_148, input_149, AND_149, input_150,
    AND_150, input_151, AND_151, input_152, OR_152, input_153, AND_153,
    input_154, OR_154, input_155, OR_155, input_156, AND_156, input_157,
    AND_157, input_158, AND_158, input_159, OR_159, OR_159_INV, CASOP;
  assign n13293 = ~n13114;
  assign n13257 = ~n13271;
  assign n11682 = ~n16904;
  assign n16904 = ~n12618 ^ P2_IR_REG_28__SCAN_IN;
  assign n21822 = ~n12627 ^ n12626;
  assign n11667 = n16826 & n13554;
  assign n11671 = ~n11667;
  assign n22473 = n13256 ^ n13255;
  assign n22268 = n13239 & n13238;
  assign n22115 = ~n22135;
  assign n22334 = ~n13236 ^ n12325;
  assign n22135 = n13219 & n13218;
  assign n21536 = n13158 & n13157;
  assign n21716 = n12679 & n12678;
  assign n12577 = n11994 & n11993;
  assign n12713 = ~n12570 & ~n12569;
  assign n12732 = n11928 & n11799;
  assign n19373 = n12924 & n12923;
  assign n12329 = ~n12555 & ~n11733;
  assign n19100 = ~n19083;
  assign n18880 = ~n12817 | ~n12816;
  assign n18900 = ~n15740;
  assign n18756 = n12830 & n12829;
  assign n12841 = ~n13114;
  assign n15740 = n12806 & n12805;
  assign n13114 = ~n15739 | ~n15113;
  assign n11677 = ~n12666;
  assign n11680 = ~n12886;
  assign n22834 = ~n12669;
  assign n12636 = n12634 | P2_IR_REG_19__SCAN_IN;
  assign n12789 = ~n12642 ^ P2_IR_REG_29__SCAN_IN;
  assign n13493 = ~n12416 | ~P2_IR_REG_31__SCAN_IN;
  assign n12609 = ~n13037 & ~n11937;
  assign n13037 = ~n12122 | ~n12123;
  assign n18814 = ~n13554;
  assign n13579 = n13554 | n12520;
  assign n12406 = ~n12407 & ~P2_IR_REG_8__SCAN_IN;
  assign n12418 = n12458 & n12602;
  assign n11931 = n12090 & n12892;
  assign n17888 = P1_ADDR_REG_19__SCAN_IN & P2_ADDR_REG_19__SCAN_IN;
  assign n17889 = ~P2_ADDR_REG_19__SCAN_IN & ~P1_ADDR_REG_19__SCAN_IN;
  assign n12818 = ~P2_IR_REG_1__SCAN_IN & ~P2_IR_REG_0__SCAN_IN;
  assign n12892 = ~P2_IR_REG_4__SCAN_IN;
  assign n12090 = ~P2_IR_REG_2__SCAN_IN & ~P2_IR_REG_3__SCAN_IN;
  assign n12945 = ~P2_IR_REG_6__SCAN_IN;
  assign n13394 = n11967 & n11814;
  assign n13400 = ~n12657 | ~n13394;
  assign n12870 = ~n18880 & ~n18756;
  assign n12553 = SI_7_ | n12552;
  assign n12007 = ~n12418 | ~n11716;
  assign n11987 = n11736 & n12914;
  assign n12009 = ~n13400 | ~n12010;
  assign n22812 = n13366 & n13365;
  assign n15966 = ~n15955 | ~n15942;
  assign n12417 = ~P2_IR_REG_21__SCAN_IN & ~n12611;
  assign n12122 = n12406 & n13011;
  assign n12559 = ~n12558 | ~n12557;
  assign n12544 = ~n12542 | ~n12541;
  assign n12542 = ~P2_DATAO_REG_5__SCAN_IN | ~n13554;
  assign n11916 = ~n12577 | ~n12579;
  assign n11966 = ~n11918 | ~n12536;
  assign n12536 = ~SI_3_ | ~n12535;
  assign n13476 = n13471 & n13470;
  assign n12338 = n13377 & n12339;
  assign n12879 = n12810 | n12853;
  assign n12014 = ~n11701;
  assign n15777 = n20886 | n12751;
  assign n12310 = ~n13388 | ~n12309;
  assign n13401 = ~n13400 | ~n13399;
  assign n12334 = n12471 & P3_ADDR_REG_19__SCAN_IN;
  assign n12471 = ~P1_RD_REG_SCAN_IN;
  assign n13482 = ~n12609 | ~n12608;
  assign n19083 = n12849 & n12848;
  assign n12849 = n12845 & n12844;
  assign n15739 = n21822 & n15125;
  assign n16128 = ~n16158 ^ n16886;
  assign n16039 = ~n13302 | ~n13301;
  assign n15940 = ~n13283 | ~n15966;
  assign n15943 = ~n15955;
  assign n21950 = ~n21964;
  assign n20068 = n13440 & n15765;
  assign n19357 = ~n19373;
  assign n19193 = ~n12901 | ~n12900;
  assign n18739 = ~n15750 | ~n12872;
  assign n12006 = ~n11706 & ~n12007;
  assign n11980 = ~n11981 | ~n12712;
  assign n12407 = ~n11755 | ~n12600;
  assign n12539 = ~n12538 | ~n12537;
  assign n12538 = ~P2_DATAO_REG_4__SCAN_IN | ~n13554;
  assign n12535 = ~n12533 | ~n12532;
  assign n11971 = ~n11973;
  assign n11970 = ~n11973 & ~n12593;
  assign n11985 = n12331 & n11988;
  assign n12985 = ~n12554 ^ SI_8_;
  assign n12525 = ~n11922 | ~n12522;
  assign n12522 = ~n14417 | ~P2_DATAO_REG_0__SCAN_IN;
  assign n16712 = ~n13337 | ~n13336;
  assign n13337 = ~n22765 | ~n13257;
  assign n13477 = ~n11964 | ~n12008;
  assign n11964 = n11965 & n13411;
  assign n22813 = ~n12621 | ~n12620;
  assign n22401 = ~n13260 | ~n13259;
  assign n21198 = n12701 & n12700;
  assign n22913 = ~n13388 | ~n13387;
  assign n12169 = ~n12609 | ~n12170;
  assign n12170 = n11769 & n12417;
  assign n12171 = ~P2_IR_REG_28__SCAN_IN;
  assign n11994 = ~n11923 | ~n11810;
  assign n11923 = n13123 | n13124;
  assign n13069 = ~n12562 & ~n12561;
  assign n12327 = ~n12328 | ~n12560;
  assign n13007 = SI_9_ ^ n12559;
  assign n11990 = ~n12915 | ~n12914;
  assign n12847 = ~n12304 | ~n12531;
  assign n12340 = ~n12598 | ~n11819;
  assign n12341 = ~n13363;
  assign n13334 = ~n12595 | ~n12594;
  assign n13270 = ~n12320 | ~n11809;
  assign n13191 = ~n11915 | ~n12583;
  assign n11915 = ~n11916 | ~n11793;
  assign n11983 = ~n12713;
  assign n11998 = ~n12831 | ~n11999;
  assign n11999 = n12832 & n12852;
  assign n12000 = ~n12855 | ~n12001;
  assign n12001 = n12856 & n12857;
  assign n13091 = n13087 | n13086;
  assign n12011 = ~n11693 | ~n11701;
  assign n12309 = n16899 & n13387;
  assign n13407 = ~n22913;
  assign n13357 = ~n16716 & ~n16889;
  assign n12845 = ~n11667 | ~P1_DATAO_REG_3__SCAN_IN;
  assign n16129 = ~n16160 & ~n16118;
  assign n15704 = n15705 & n13432;
  assign n19346 = ~n19351 | ~n19213;
  assign n11973 = ~n11974 | ~n13298;
  assign n11974 = ~n11975 | ~n12593;
  assign n11975 = ~n13269;
  assign n12331 = ~n11756 | ~n12553;
  assign n12332 = ~n12549;
  assign n13405 = ~n13403 | ~n13404;
  assign n15968 = n15971 & n13462;
  assign n15748 = n13422 | n13421;
  assign n16158 = ~n13322 | ~n13321;
  assign n22389 = ~n22401 ^ n22256;
  assign n21034 = ~n13420 & ~n13419;
  assign n19201 = ~n19346 | ~n12930;
  assign n12696 = ~n13037 & ~n12007;
  assign n12734 = ~n11935 | ~n12418;
  assign n12328 = ~n13036;
  assign n13071 = ~n11935 | ~n12602;
  assign n12552 = ~n12551 | ~n12550;
  assign n12548 = ~n12547 | ~n12546;
  assign n12547 = ~P2_DATAO_REG_6__SCAN_IN | ~n13554;
  assign n12961 = ~n12123 | ~n12600;
  assign n12405 = ~n12818 | ~n12796;
  assign n12796 = ~P2_IR_REG_2__SCAN_IN;
  assign n12322 = ~n12591;
  assign n12530 = ~n12529 | ~n12528;
  assign n12529 = n12527 | n18818;
  assign n12336 = ~n12337 | ~n17888;
  assign n12335 = ~n12334 | ~n17889;
  assign n12337 = ~P3_ADDR_REG_19__SCAN_IN & ~P2_RD_REG_SCAN_IN;
  assign n20545 = ~n13102 | ~n13101;
  assign n12901 = n12897 & n12896;
  assign n12897 = ~n11667 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n21794 = n12662 & n12661;
  assign n11992 = ~n13481 | ~n13480;
  assign n19333 = ~n12890 & ~n12889;
  assign n19167 = ~n12840 & ~n12839;
  assign n12839 = ~n12838 | ~n12837;
  assign n15689 = ~n12794 & ~n12793;
  assign n15691 = ~n12865 & ~n12864;
  assign n16716 = ~n16712;
  assign n16160 = ~n16158;
  assign n16041 = ~n16039;
  assign n15955 = n13274 & n13273;
  assign n22243 = ~n22268;
  assign n21964 = n13194 & n13193;
  assign n21815 = ~n21794;
  assign n21031 = n12722 & n12721;
  assign n20886 = ~n12741 | ~n12740;
  assign n20409 = ~n13075 | ~n13074;
  assign n12830 = n12825 & n12419;
  assign n12825 = ~n11934 | ~n11691;
  assign n19696 = ~n12967 | ~n12966;
  assign n12669 = ~n12639 ^ P2_IR_REG_30__SCAN_IN;
  assign n12639 = ~n22929 | ~P2_IR_REG_31__SCAN_IN;
  assign n12642 = ~n12169 | ~P2_IR_REG_31__SCAN_IN;
  assign n11936 = n12006 & n11763;
  assign n13123 = ~n11924 | ~n11795;
  assign n12330 = ~n13007;
  assign n13009 = ~n12123 | ~n12406;
  assign n12988 = ~n12916 & ~n12407;
  assign n12958 = ~n12552 ^ SI_7_;
  assign n12943 = ~n12548 ^ n13706;
  assign n12914 = ~n12544 ^ n12543;
  assign n12915 = ~n11917 | ~n12540;
  assign n11917 = ~n11966 | ~n12898;
  assign n11932 = ~n12818 | ~n12090;
  assign n12846 = ~n12535 ^ n12534;
  assign n13319 = ~n11968 | ~n11969;
  assign n11969 = ~n11970 & ~n11817;
  assign n11968 = ~n13270 | ~n11971;
  assign n12307 = ~n12308 | ~n12674;
  assign n12308 = ~n12578;
  assign n11993 = ~n13151;
  assign n12804 = ~n11976 | ~n12526;
  assign n12526 = ~SI_1_ | ~n12525;
  assign n12802 = ~n12530 ^ n13599;
  assign n12828 = ~n12525 ^ n13553;
  assign n14417 = n13554 & SI_0_;
  assign n19213 = n12901 & n12900;
  assign n22901 = ~n22813;
  assign n20243 = n13045 & n13044;
  assign n20081 = n13018 & n13017;
  assign n13152 = ~n11994;
  assign n13006 = ~n12555 & ~n12556;
  assign n23453 = ~n13385 ^ n13384;
  assign n22863 = ~n11978 ^ n11977;
  assign n11977 = ~n13377;
  assign n11979 = ~n12340;
  assign n22784 = ~n13363 ^ n13362;
  assign n13362 = ~n12598 | ~n12597;
  assign n22765 = n13334 ^ n13333;
  assign n22739 = n13319 ^ n13318;
  assign n22645 = n13299 ^ n13298;
  assign n13299 = ~n11972 | ~n12593;
  assign n22559 = n13270 ^ n13269;
  assign n12694 = n11982 & n11788;
  assign n11982 = ~n11983 | ~n11984;
  assign n12002 = n12003 & n11830;
  assign n18818 = ~n13554;
  assign n11691 = n11682 & n11933;
  assign n11693 = ~n12015 | ~n11759;
  assign n11697 = n11667 & P1_DATAO_REG_6__SCAN_IN;
  assign n11698 = n11992 & n11827;
  assign n11935 = ~n13037;
  assign n12899 = n16826 & n18814;
  assign n12883 = n22834 | n12789;
  assign n11701 = n13189 | n13188;
  assign n16189 = ~n22812 ^ n16892;
  assign n11929 = ~n18735;
  assign n13159 = n22834 & n22774;
  assign n21696 = ~n15785 & ~n13450;
  assign n11706 = n12624 | n12607;
  assign n12608 = ~P2_IR_REG_21__SCAN_IN;
  assign n15785 = n21716 & n21788;
  assign n11716 = n12715 & n12604;
  assign n16185 = ~n16712 ^ n16889;
  assign n11733 = n12556 | n12330;
  assign n13434 = n19556 | n19696;
  assign n11736 = n12943 & n12553;
  assign n12706 = ~n22834 & ~n12789;
  assign n19909 = n12997 & n12996;
  assign n11755 = n12945 & n12601;
  assign n11756 = n12958 | n12332;
  assign n15971 = ~n16041 | ~n16883;
  assign n11758 = ~n12577 & ~n12578;
  assign n11759 = n12673 | n12672;
  assign n11763 = n12417 & n12612;
  assign n11768 = n12417 & n12470;
  assign n11769 = n12470 & n12171;
  assign n11842 = ~P1_DATAO_REG_1__SCAN_IN;
  assign n11774 = n13292 & n13297;
  assign n11779 = n12971 & n12973;
  assign n11780 = n12879 & n11996;
  assign n12811 = n12669 & n12789;
  assign n11788 = SI_15_ | n12571;
  assign n11984 = ~n12712;
  assign n12916 = ~n11931 | ~n12818;
  assign n12123 = ~n12916;
  assign n11933 = ~n16935;
  assign n11793 = n12306 & n12658;
  assign n11795 = n11980 & n12575;
  assign n12600 = ~P2_IR_REG_5__SCAN_IN;
  assign n11799 = SI_13_ | n12567;
  assign n11801 = SI_12_ | n12566;
  assign n11802 = n13554 & P1_DATAO_REG_2__SCAN_IN;
  assign n11803 = n13554 & P1_DATAO_REG_1__SCAN_IN;
  assign n11981 = n12693 & n11788;
  assign n11807 = n12324 & n13255;
  assign n11809 = n12321 & n12592;
  assign n11810 = SI_17_ | n12504;
  assign n11814 = n12655 | n16194;
  assign n11815 = n12609 & n12417;
  assign n11817 = SI_26_ & n12484;
  assign n11819 = n12341 & n12597;
  assign n12339 = ~n12599;
  assign n11827 = n22281 & n21658;
  assign n11830 = n13500 | n13499;
  assign n16909 = ~n12615 ^ n12614;
  assign n11934 = ~n16909;
  assign n15125 = n12632 & n13482;
  assign n12584 = ~n13191 | ~n13190;
  assign n11918 = ~n12847 | ~n12846;
  assign n11976 = ~n12828 | ~n12826;
  assign n11922 = ~n12521 | ~P1_DATAO_REG_0__SCAN_IN;
  assign n11924 = ~n12713 | ~n11981;
  assign n12569 = ~n12732 & ~n12731;
  assign n11928 = ~n12316 | ~n12315;
  assign n12316 = ~n12317 | ~n11801;
  assign n12891 = ~n11932 | ~P2_IR_REG_31__SCAN_IN;
  assign n16826 = ~n11934 | ~n11682;
  assign n11937 = ~n12006;
  assign n12416 = ~n11936 | ~n11935;
  assign n12628 = ~n12609;
  assign n11965 = ~n13405 | ~n12009;
  assign n19277 = ~n11966 ^ n12898;
  assign n11967 = ~n22813 | ~n13293;
  assign n11972 = ~n13270 | ~n13269;
  assign n12621 = ~n22863 | ~n13257;
  assign n11978 = ~n12599 & ~n11979;
  assign n11986 = ~n12915 | ~n11987;
  assign n12987 = ~n11986 | ~n11985;
  assign n12944 = ~n11990 | ~n12545;
  assign n11988 = ~n11736 | ~n11989;
  assign n11989 = ~n12545;
  assign n11991 = ~n13476 | ~n21976;
  assign n12003 = ~n11991 | ~n11698;
  assign n13487 = ~n11992 | ~n22281;
  assign n12801 = ~n16826 | ~n11802;
  assign n12904 = ~n11997 | ~n11995;
  assign n11995 = ~n11780 | ~n12878;
  assign n11996 = ~n12877 | ~n12876;
  assign n11997 = ~n12000 | ~n11998;
  assign P2_U3328_Lock = ~n12002 | ~n12314;
  assign n12976 = ~n12004 | ~n11779;
  assign n12004 = ~n12005 | ~n12968;
  assign n12005 = ~n12935 | ~n12934;
  assign n12008 = ~n13376 | ~n13405;
  assign n12010 = ~n16189;
  assign n13209 = ~n12012 | ~n12011;
  assign n12012 = ~n13180 | ~n12013;
  assign n12013 = ~n12014 & ~n13186;
  assign n12015 = ~n12016 | ~n13181;
  assign n12016 = ~n13186;
  assign n13317 = ~n12017 | ~n13313;
  assign n12017 = ~n12018 | ~n11774;
  assign n12018 = ~n13285 | ~n13284;
  assign n13119 = ~n12021 | ~n12019;
  assign n12019 = ~n12020 & ~n12786;
  assign n12020 = ~n13117 & ~n13118;
  assign n13118 = ~n13091 | ~n13090;
  assign n12021 = ~n12022 | ~n13113;
  assign n12022 = ~n13112 | ~n13115;
  assign n12922 = ~n11667 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n12965 = ~n11667 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n12995 = ~n11667 | ~P1_DATAO_REG_8__SCAN_IN;
  assign n12641 = ~n12169;
  assign n12637 = ~n12609 | ~n11768;
  assign n12304 = ~n12804 | ~n12802;
  assign n12659 = ~n12305 | ~n12579;
  assign n12305 = n12577 | n12307;
  assign n12306 = ~n12307 | ~n12579;
  assign n13389 = ~n12310 | ~n13293;
  assign n12312 = ~n13476;
  assign n12314 = ~n12313 | ~n12311;
  assign n12311 = ~n12312 | ~n21976;
  assign n12313 = ~n13475 & ~n13487;
  assign n12755 = ~n12316;
  assign n12315 = ~n12754;
  assign n12317 = ~n12319 | ~n12318;
  assign n12318 = ~n13092;
  assign n12319 = ~n13093;
  assign n12320 = ~n13236 | ~n11807;
  assign n12321 = ~n11807 | ~n12322;
  assign n13256 = ~n12323 | ~n12591;
  assign n12323 = ~n13236 | ~n13235;
  assign n12324 = ~n12325 | ~n12591;
  assign n12325 = ~n13235;
  assign n13035 = ~n12326 | ~n12560;
  assign n12326 = ~n12329;
  assign n12561 = ~n12329 & ~n12327;
  assign n12333 = ~n12944 | ~n12943;
  assign n12960 = ~n12333 | ~n12549;
  assign n13554 = ~n12336 | ~n12335;
  assign n13380 = ~n12340 | ~n12338;
  assign n12842 = ~n12405 | ~P2_IR_REG_31__SCAN_IN;
  assign n16954 = ~n12799 | ~n12405;
  assign n12419 = ~n16826 | ~n11803;
  assign n12458 = n12603 & n13095;
  assign n12886 = ~n12811;
  assign n12470 = n12617 & n12616;
  assign n12984 = n13005 | n12999;
  assign n13141 = n13122 & n15779;
  assign n13484 = ~n13482;
  assign n12554 = ~n12519 | ~n12518;
  assign n12528 = ~n18818 | ~P1_DATAO_REG_2__SCAN_IN;
  assign n19889 = ~n15704;
  assign n12517 = ~n12516 | ~n12515;
  assign n12556 = ~SI_8_ & ~n12554;
  assign n12602 = ~P2_IR_REG_10__SCAN_IN;
  assign n12520 = ~SI_0_;
  assign n12898 = ~n12539 ^ n13649;
  assign n12826 = ~n12524 | ~n12523;
  assign n12473 = ~P2_DATAO_REG_30__SCAN_IN | ~n13554;
  assign n12472 = ~n18818 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n13378 = ~n12473 | ~n12472;
  assign n13377 = SI_30_ ^ n13378;
  assign n12475 = ~P2_DATAO_REG_29__SCAN_IN | ~n13554;
  assign n12474 = ~n18814 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n12476 = ~n12475 | ~n12474;
  assign n12599 = ~SI_29_ & ~n12476;
  assign n13363 = ~SI_29_ ^ n12476;
  assign n12478 = ~P2_DATAO_REG_28__SCAN_IN | ~n13554;
  assign n12477 = ~P1_DATAO_REG_28__SCAN_IN | ~n18814;
  assign n12596 = ~n12478 | ~n12477;
  assign n13333 = SI_28_ ^ n12596;
  assign n12480 = ~P2_DATAO_REG_27__SCAN_IN | ~n13554;
  assign n12479 = ~n18814 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n12481 = ~n12480 | ~n12479;
  assign n12595 = ~SI_27_ | ~n12481;
  assign n13318 = SI_27_ ^ n12481;
  assign n12483 = ~P2_DATAO_REG_26__SCAN_IN | ~n13554;
  assign n12482 = ~n18814 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n12484 = ~n12483 | ~n12482;
  assign n13298 = SI_26_ ^ n12484;
  assign n12486 = ~P2_DATAO_REG_25__SCAN_IN | ~n13554;
  assign n12485 = ~n18814 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n12487 = ~n12486 | ~n12485;
  assign n12593 = ~SI_25_ | ~n12487;
  assign n13269 = SI_25_ ^ n12487;
  assign n12489 = ~P2_DATAO_REG_24__SCAN_IN | ~n13554;
  assign n12488 = ~n18814 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n12490 = ~n12489 | ~n12488;
  assign n12592 = ~SI_24_ | ~n12490;
  assign n13255 = SI_24_ ^ n12490;
  assign n12492 = ~P2_DATAO_REG_22__SCAN_IN | ~n13554;
  assign n12491 = ~n18814 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n12493 = ~n12492 | ~n12491;
  assign n12587 = ~SI_22_ | ~n12493;
  assign n13215 = SI_22_ ^ n12493;
  assign n12495 = ~P2_DATAO_REG_21__SCAN_IN | ~n13554;
  assign n12494 = ~n18814 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n12496 = ~n12495 | ~n12494;
  assign n12585 = ~SI_21_ | ~n12496;
  assign n15172 = ~SI_21_;
  assign n13190 = ~n15172 ^ n12496;
  assign n12498 = ~P2_DATAO_REG_19__SCAN_IN | ~n13554;
  assign n12497 = ~n18814 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n12499 = ~n12498 | ~n12497;
  assign n12579 = ~SI_19_ | ~n12499;
  assign n12674 = SI_19_ ^ n12499;
  assign n12501 = ~P2_DATAO_REG_18__SCAN_IN | ~n13554;
  assign n12500 = ~n18814 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n12576 = ~n12501 | ~n12500;
  assign n12578 = ~SI_18_ & ~n12576;
  assign n12503 = ~P2_DATAO_REG_17__SCAN_IN | ~n13554;
  assign n12502 = ~n18814 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n12504 = ~n12503 | ~n12502;
  assign n13124 = ~SI_17_ ^ n12504;
  assign n12506 = ~P2_DATAO_REG_15__SCAN_IN | ~n13554;
  assign n12505 = ~n18814 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n12571 = ~n12506 | ~n12505;
  assign n12508 = ~P2_DATAO_REG_14__SCAN_IN | ~n13554;
  assign n12507 = ~n18814 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n12568 = ~n12508 | ~n12507;
  assign n12570 = ~SI_14_ & ~n12568;
  assign n12510 = ~P2_DATAO_REG_13__SCAN_IN | ~n13554;
  assign n12509 = ~n18814 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n12567 = ~n12510 | ~n12509;
  assign n12512 = ~P2_DATAO_REG_12__SCAN_IN | ~n13554;
  assign n12511 = ~n18814 | ~P1_DATAO_REG_12__SCAN_IN;
  assign n12566 = ~n12512 | ~n12511;
  assign n12514 = ~P2_DATAO_REG_11__SCAN_IN | ~n13554;
  assign n12513 = ~n18814 | ~P1_DATAO_REG_11__SCAN_IN;
  assign n12563 = ~n12514 | ~n12513;
  assign n12565 = ~SI_11_ & ~n12563;
  assign n12516 = ~P2_DATAO_REG_10__SCAN_IN | ~n13554;
  assign n12515 = ~n18814 | ~P1_DATAO_REG_10__SCAN_IN;
  assign n12562 = ~SI_10_ & ~n12517;
  assign n13036 = ~SI_10_ ^ n12517;
  assign n12519 = ~P2_DATAO_REG_8__SCAN_IN | ~n13554;
  assign n12518 = ~n18814 | ~P1_DATAO_REG_8__SCAN_IN;
  assign n12521 = ~n13579;
  assign n13553 = ~SI_1_;
  assign n12524 = n13554 | n11842;
  assign n12523 = ~n13554 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n12527 = ~P2_DATAO_REG_2__SCAN_IN;
  assign n13599 = ~SI_2_;
  assign n12531 = ~SI_2_ | ~n12530;
  assign n12533 = ~P2_DATAO_REG_3__SCAN_IN | ~n13554;
  assign n12532 = ~n18814 | ~P1_DATAO_REG_3__SCAN_IN;
  assign n12534 = ~SI_3_;
  assign n12537 = ~n18814 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n13649 = ~SI_4_;
  assign n12540 = ~SI_4_ | ~n12539;
  assign n12541 = ~n18814 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n12543 = ~SI_5_;
  assign n12545 = ~SI_5_ | ~n12544;
  assign n12546 = ~n18814 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n13706 = ~SI_6_;
  assign n12549 = ~SI_6_ | ~n12548;
  assign n12551 = ~P2_DATAO_REG_7__SCAN_IN | ~n13554;
  assign n12550 = ~n18814 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n12555 = ~n12987 & ~n12985;
  assign n12558 = ~P2_DATAO_REG_9__SCAN_IN | ~n13554;
  assign n12557 = ~n18814 | ~P1_DATAO_REG_9__SCAN_IN;
  assign n12560 = ~SI_9_ | ~n12559;
  assign n13068 = ~SI_11_ ^ n12563;
  assign n12564 = ~n13069 & ~n13068;
  assign n13093 = ~n12565 & ~n12564;
  assign n13092 = ~SI_12_ ^ n12566;
  assign n12754 = ~SI_13_ ^ n12567;
  assign n12731 = ~SI_14_ ^ n12568;
  assign n12712 = ~SI_15_ ^ n12571;
  assign n12573 = ~P2_DATAO_REG_16__SCAN_IN | ~n13554;
  assign n12572 = ~n18814 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n12574 = ~n12573 | ~n12572;
  assign n12693 = SI_16_ ^ n12574;
  assign n12575 = ~SI_16_ | ~n12574;
  assign n13151 = ~SI_18_ ^ n12576;
  assign n12581 = ~P2_DATAO_REG_20__SCAN_IN | ~n13554;
  assign n12580 = ~n18814 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n12582 = ~n12581 | ~n12580;
  assign n12658 = SI_20_ ^ n12582;
  assign n12583 = ~SI_20_ | ~n12582;
  assign n13216 = ~n12585 | ~n12584;
  assign n12586 = ~n13215 | ~n13216;
  assign n13236 = ~n12587 | ~n12586;
  assign n12589 = ~P2_DATAO_REG_23__SCAN_IN | ~n13554;
  assign n12588 = ~n18814 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n12590 = ~n12589 | ~n12588;
  assign n13235 = SI_23_ ^ n12590;
  assign n12591 = ~SI_23_ | ~n12590;
  assign n12594 = ~n13318 | ~n13319;
  assign n12598 = ~n13333 | ~n13334;
  assign n12597 = ~SI_28_ | ~n12596;
  assign n12601 = ~P2_IR_REG_7__SCAN_IN;
  assign n12990 = ~P2_IR_REG_8__SCAN_IN;
  assign n12603 = ~P2_IR_REG_12__SCAN_IN;
  assign n13095 = ~P2_IR_REG_11__SCAN_IN;
  assign n12715 = ~P2_IR_REG_13__SCAN_IN & ~P2_IR_REG_14__SCAN_IN;
  assign n12604 = ~P2_IR_REG_15__SCAN_IN;
  assign n12605 = ~P2_IR_REG_18__SCAN_IN;
  assign n13126 = ~P2_IR_REG_17__SCAN_IN;
  assign n12624 = ~n12605 | ~n13126;
  assign n12606 = ~P2_IR_REG_16__SCAN_IN & ~P2_IR_REG_19__SCAN_IN;
  assign n12626 = ~P2_IR_REG_20__SCAN_IN;
  assign n12607 = ~n12606 | ~n12626;
  assign n13483 = ~P2_IR_REG_22__SCAN_IN;
  assign n12610 = ~P2_IR_REG_23__SCAN_IN;
  assign n12611 = ~n13483 | ~n12610;
  assign n12612 = ~P2_IR_REG_24__SCAN_IN & ~P2_IR_REG_25__SCAN_IN;
  assign n12613 = ~P2_IR_REG_31__SCAN_IN | ~P2_IR_REG_26__SCAN_IN;
  assign n12615 = ~n13493 | ~n12613;
  assign n12614 = ~P2_IR_REG_27__SCAN_IN;
  assign n12617 = ~P2_IR_REG_24__SCAN_IN & ~P2_IR_REG_26__SCAN_IN;
  assign n12616 = ~P2_IR_REG_27__SCAN_IN & ~P2_IR_REG_25__SCAN_IN;
  assign n12618 = ~n12637 | ~P2_IR_REG_31__SCAN_IN;
  assign n12619 = ~P1_DATAO_REG_30__SCAN_IN;
  assign n12620 = n11671 | n12619;
  assign n12622 = ~P2_IR_REG_16__SCAN_IN;
  assign n12623 = ~n12696 | ~n12622;
  assign n13127 = ~n12623 | ~P2_IR_REG_31__SCAN_IN;
  assign n12625 = ~n12624 | ~P2_IR_REG_31__SCAN_IN;
  assign n12634 = ~n13127 | ~n12625;
  assign n12627 = ~n12636 | ~P2_IR_REG_31__SCAN_IN;
  assign n12629 = ~n12628 | ~P2_IR_REG_31__SCAN_IN;
  assign n12631 = ~n12629 | ~P2_IR_REG_21__SCAN_IN;
  assign n12630 = ~n12608 | ~P2_IR_REG_31__SCAN_IN;
  assign n12632 = ~n12631 | ~n12630;
  assign n12633 = ~n13482 | ~P2_IR_REG_31__SCAN_IN;
  assign n15126 = ~n12633 ^ P2_IR_REG_22__SCAN_IN;
  assign n12635 = ~n12634 | ~P2_IR_REG_19__SCAN_IN;
  assign n21658 = ~n12636 | ~n12635;
  assign n15113 = ~n15126 & ~n21658;
  assign n12638 = ~P2_IR_REG_29__SCAN_IN;
  assign n22929 = ~n12641 | ~n12638;
  assign n12640 = ~P2_IR_REG_31__SCAN_IN;
  assign n22774 = ~n12789;
  assign n12645 = ~n11677 | ~P2_REG0_REG_31__SCAN_IN;
  assign n12643 = ~P2_REG2_REG_31__SCAN_IN;
  assign n12644 = n12883 | n12643;
  assign n12647 = n12645 & n12644;
  assign n12860 = n22834 & n12789;
  assign n12646 = ~n12860 | ~P2_REG1_REG_31__SCAN_IN;
  assign n16899 = ~n12647 | ~n12646;
  assign n22820 = ~n16899;
  assign n12649 = ~n22820 & ~n21822;
  assign n21976 = ~n15125;
  assign n15118 = ~n21822 & ~n21976;
  assign n12648 = ~n12869 & ~n15118;
  assign n12655 = ~n12649 & ~n12648;
  assign n12652 = ~n12860 | ~P2_REG1_REG_30__SCAN_IN;
  assign n12650 = ~P2_REG2_REG_30__SCAN_IN;
  assign n12651 = n12883 | n12650;
  assign n12654 = n12652 & n12651;
  assign n12653 = ~n13159 | ~P2_REG0_REG_30__SCAN_IN;
  assign n16895 = ~n12654 | ~n12653;
  assign n16194 = ~n16895;
  assign n12656 = ~n16895 | ~n13293;
  assign n12657 = ~n22901 | ~n12656;
  assign n21872 = n12659 ^ n12658;
  assign n12662 = ~n21872 | ~n13257;
  assign n12660 = ~P1_DATAO_REG_20__SCAN_IN;
  assign n12661 = n11671 | n12660;
  assign n12665 = ~n12860 | ~P2_REG1_REG_20__SCAN_IN;
  assign n12663 = ~P2_REG2_REG_20__SCAN_IN;
  assign n12664 = n12883 | n12663;
  assign n12668 = ~n12665 | ~n12664;
  assign n12666 = ~n13159;
  assign n12667 = n13159 & P2_REG0_REG_20__SCAN_IN;
  assign n12671 = ~n12668 & ~n12667;
  assign n12908 = P2_REG3_REG_4__SCAN_IN & P2_REG3_REG_3__SCAN_IN;
  assign n12938 = ~n12908 | ~P2_REG3_REG_5__SCAN_IN;
  assign n17015 = ~P2_REG3_REG_6__SCAN_IN;
  assign n12950 = ~n12938 & ~n17015;
  assign n12977 = ~n12950 | ~P2_REG3_REG_7__SCAN_IN;
  assign n17049 = ~P2_REG3_REG_8__SCAN_IN;
  assign n13019 = ~n12977 & ~n17049;
  assign n13048 = ~n13019 | ~P2_REG3_REG_9__SCAN_IN;
  assign n17266 = ~P2_REG3_REG_10__SCAN_IN;
  assign n13076 = ~n13048 & ~n17266;
  assign n13103 = ~n13076 | ~P2_REG3_REG_11__SCAN_IN;
  assign n17095 = ~P2_REG3_REG_12__SCAN_IN;
  assign n12763 = ~n13103 & ~n17095;
  assign n12742 = ~n12763 | ~P2_REG3_REG_13__SCAN_IN;
  assign n17228 = ~P2_REG3_REG_14__SCAN_IN;
  assign n12725 = ~n12742 & ~n17228;
  assign n12704 = ~n12725 | ~P2_REG3_REG_15__SCAN_IN;
  assign n17103 = ~P2_REG3_REG_16__SCAN_IN;
  assign n13138 = ~n12704 & ~n17103;
  assign n13165 = ~n13138 | ~P2_REG3_REG_17__SCAN_IN;
  assign n17143 = ~P2_REG3_REG_18__SCAN_IN;
  assign n12685 = ~n13165 & ~n17143;
  assign n13200 = n12685 & P2_REG3_REG_19__SCAN_IN;
  assign n21811 = P2_REG3_REG_20__SCAN_IN ^ n13200;
  assign n12670 = ~n21811 | ~n11680;
  assign n21939 = ~n12671 | ~n12670;
  assign n13416 = ~n21939;
  assign n13187 = ~n21815 & ~n13416;
  assign n13395 = ~n12841;
  assign n12673 = ~n13187 & ~n13395;
  assign n15787 = ~n21794 & ~n21939;
  assign n12672 = ~n15787 & ~n13293;
  assign n21661 = n11758 ^ n12674;
  assign n12679 = ~n21661 | ~n13257;
  assign n12675 = ~P1_DATAO_REG_19__SCAN_IN;
  assign n12677 = n11671 | n12675;
  assign n12676 = n16826 | n21658;
  assign n12678 = n12677 & n12676;
  assign n12690 = ~n21716 | ~n12841;
  assign n12681 = ~n12860 | ~P2_REG1_REG_19__SCAN_IN;
  assign n12680 = ~n13159 | ~P2_REG0_REG_19__SCAN_IN;
  assign n12684 = ~n12681 | ~n12680;
  assign n12682 = ~P2_REG2_REG_19__SCAN_IN;
  assign n12683 = ~n12883 & ~n12682;
  assign n12688 = n12684 | n12683;
  assign n21706 = ~P2_REG3_REG_19__SCAN_IN ^ n12685;
  assign n12686 = ~n21706;
  assign n12687 = n11680 & n12686;
  assign n21788 = n12688 | n12687;
  assign n21496 = ~n21788;
  assign n12869 = ~n13114;
  assign n12689 = ~n21496 | ~n13114;
  assign n13183 = n12690 & n12689;
  assign n12692 = ~n21716 | ~n13114;
  assign n12691 = ~n21496 | ~n13293;
  assign n13182 = ~n12692 | ~n12691;
  assign n13181 = ~n13183 & ~n13182;
  assign n21168 = n12694 ^ n12693;
  assign n12701 = ~n21168 | ~n13257;
  assign n12695 = ~P1_DATAO_REG_16__SCAN_IN;
  assign n12699 = n11671 | n12695;
  assign n12697 = n12696 | n12640;
  assign n17155 = ~n12697 ^ P2_IR_REG_16__SCAN_IN;
  assign n17120 = ~n17155;
  assign n12698 = n16826 | n17120;
  assign n12700 = n12699 & n12698;
  assign n12703 = ~n12860 | ~P2_REG1_REG_16__SCAN_IN;
  assign n12702 = ~n11677 | ~P2_REG0_REG_16__SCAN_IN;
  assign n12711 = n12703 & n12702;
  assign n21211 = P2_REG3_REG_16__SCAN_IN ^ n12704;
  assign n12705 = ~n21211;
  assign n12709 = ~n11680 | ~n12705;
  assign n12707 = ~P2_REG2_REG_16__SCAN_IN;
  assign n12708 = n12883 | n12707;
  assign n12710 = n12709 & n12708;
  assign n21364 = ~n12711 | ~n12710;
  assign n13421 = ~n21198 & ~n21364;
  assign n21003 = n12713 ^ n12712;
  assign n14656 = ~n21003;
  assign n12722 = ~n14656 | ~n13257;
  assign n12714 = ~P1_DATAO_REG_15__SCAN_IN;
  assign n12720 = n11671 | n12714;
  assign n12716 = ~n12734;
  assign n12717 = ~n12716 | ~n12715;
  assign n12718 = ~n12717 | ~P2_IR_REG_31__SCAN_IN;
  assign n17210 = ~n12718 ^ P2_IR_REG_15__SCAN_IN;
  assign n17131 = ~n17210;
  assign n12719 = n16826 | n17131;
  assign n12721 = n12720 & n12719;
  assign n12724 = ~n12860 | ~P2_REG1_REG_15__SCAN_IN;
  assign n12723 = ~n11677 | ~P2_REG0_REG_15__SCAN_IN;
  assign n12730 = n12724 & n12723;
  assign n21044 = P2_REG3_REG_15__SCAN_IN ^ n12725;
  assign n12728 = ~n11680 | ~n21044;
  assign n12726 = ~P2_REG2_REG_15__SCAN_IN;
  assign n12727 = n12883 | n12726;
  assign n12729 = n12728 & n12727;
  assign n21192 = ~n12730 | ~n12729;
  assign n13419 = ~n21031 & ~n21192;
  assign n13121 = ~n13421 & ~n13419;
  assign n15778 = ~n21031 | ~n21192;
  assign n20842 = n12732 ^ n12731;
  assign n14637 = ~n20842;
  assign n12741 = ~n14637 | ~n13257;
  assign n12733 = ~P1_DATAO_REG_14__SCAN_IN;
  assign n12739 = n11671 | n12733;
  assign n12757 = ~n12734 | ~P2_IR_REG_31__SCAN_IN;
  assign n12735 = ~n12757;
  assign n12736 = ~n12735 & ~P2_IR_REG_13__SCAN_IN;
  assign n12737 = ~n12736 & ~n12640;
  assign n17229 = ~P2_IR_REG_14__SCAN_IN ^ n12737;
  assign n12738 = n17229 | n16826;
  assign n12740 = n12739 & n12738;
  assign n20861 = ~P2_REG3_REG_14__SCAN_IN ^ n12742;
  assign n12744 = ~n11680 | ~n20861;
  assign n12743 = ~n12860 | ~P2_REG1_REG_14__SCAN_IN;
  assign n12749 = n12744 & n12743;
  assign n12747 = ~n11677 | ~P2_REG0_REG_14__SCAN_IN;
  assign n12745 = ~P2_REG2_REG_14__SCAN_IN;
  assign n12746 = n12883 | n12745;
  assign n12748 = n12747 & n12746;
  assign n21025 = ~n12749 | ~n12748;
  assign n12751 = ~n21025;
  assign n12750 = n15777 & n13293;
  assign n12778 = n15778 & n12750;
  assign n12753 = ~n15777 | ~n13114;
  assign n13418 = ~n20886 | ~n12751;
  assign n12752 = ~n13418 | ~n12869;
  assign n12774 = ~n12753 | ~n12752;
  assign n20677 = n12755 ^ n12754;
  assign n14617 = ~n20677;
  assign n12762 = ~n14617 | ~n13257;
  assign n12756 = ~P1_DATAO_REG_13__SCAN_IN;
  assign n12760 = n11671 | n12756;
  assign n17238 = ~n12757 ^ P2_IR_REG_13__SCAN_IN;
  assign n12758 = ~n17238;
  assign n12759 = n16826 | n12758;
  assign n12761 = n12760 & n12759;
  assign n20724 = n12762 & n12761;
  assign n12772 = ~n20724 | ~n12841;
  assign n20721 = P2_REG3_REG_13__SCAN_IN ^ n12763;
  assign n12765 = ~n11680 | ~n20721;
  assign n12764 = ~n11677 | ~P2_REG0_REG_13__SCAN_IN;
  assign n12770 = n12765 & n12764;
  assign n12768 = ~n12860 | ~P2_REG1_REG_13__SCAN_IN;
  assign n12766 = ~P2_REG2_REG_13__SCAN_IN;
  assign n12767 = n12883 | n12766;
  assign n12769 = n12768 & n12767;
  assign n20874 = ~n12770 | ~n12769;
  assign n12771 = n20874 | n13293;
  assign n12775 = ~n12772 | ~n12771;
  assign n20524 = ~n20874;
  assign n15716 = ~n20724 & ~n20524;
  assign n12773 = n12775 | n15716;
  assign n12786 = ~n12774 | ~n12773;
  assign n12776 = ~n12775;
  assign n12781 = ~n12786 & ~n12776;
  assign n12777 = ~n12781 | ~n20874;
  assign n12785 = ~n12778 | ~n12777;
  assign n12780 = ~n13419;
  assign n12779 = n13418 & n13114;
  assign n12783 = n12780 & n12779;
  assign n20708 = ~n20724;
  assign n12782 = ~n12781 | ~n20708;
  assign n12784 = ~n12783 | ~n12782;
  assign n13120 = ~n12785 | ~n12784;
  assign n12788 = ~n12860 | ~P2_REG1_REG_2__SCAN_IN;
  assign n12787 = ~n13159 | ~P2_REG0_REG_2__SCAN_IN;
  assign n12794 = ~n12788 | ~n12787;
  assign n12792 = ~n12811 | ~P2_REG3_REG_2__SCAN_IN;
  assign n12790 = ~P2_REG2_REG_2__SCAN_IN;
  assign n12791 = n12883 | n12790;
  assign n12793 = ~n12792 | ~n12791;
  assign n12808 = ~n15689 | ~n12841;
  assign n12795 = n12640 | n12818;
  assign n12798 = ~n12795 | ~P2_IR_REG_2__SCAN_IN;
  assign n12797 = ~n12796 | ~P2_IR_REG_31__SCAN_IN;
  assign n12799 = ~n12798 | ~n12797;
  assign n12800 = n16826 | n16954;
  assign n12806 = n12801 & n12800;
  assign n12803 = ~n12802;
  assign n18972 = ~n12804 ^ n12803;
  assign n12805 = ~n12899 | ~n18972;
  assign n12807 = ~n15740 | ~n13114;
  assign n12853 = ~n12808 | ~n12807;
  assign n12809 = ~n12853 | ~n18900;
  assign n12832 = n12809 & n13293;
  assign n19078 = ~n15689;
  assign n12810 = n19078 & n18900;
  assign n12813 = ~n12706 | ~P2_REG2_REG_1__SCAN_IN;
  assign n12812 = ~n12811 | ~P2_REG3_REG_1__SCAN_IN;
  assign n12817 = n12813 & n12812;
  assign n12815 = ~n12860 | ~P2_REG1_REG_1__SCAN_IN;
  assign n12814 = ~n13159 | ~P2_REG0_REG_1__SCAN_IN;
  assign n12816 = n12815 & n12814;
  assign n12824 = ~n12818;
  assign n12819 = ~P2_IR_REG_1__SCAN_IN;
  assign n12822 = ~n12819 | ~P2_IR_REG_31__SCAN_IN;
  assign n12866 = ~P2_IR_REG_0__SCAN_IN;
  assign n12820 = ~P2_IR_REG_31__SCAN_IN | ~P2_IR_REG_0__SCAN_IN;
  assign n12821 = ~n12820 | ~P2_IR_REG_1__SCAN_IN;
  assign n12823 = ~n12822 | ~n12821;
  assign n16935 = ~n12824 | ~n12823;
  assign n12827 = ~n12826;
  assign n18819 = ~n12828 ^ n12827;
  assign n12829 = ~n12899 | ~n18819;
  assign n12831 = ~n12879 | ~n12870;
  assign n12834 = ~n12860 | ~P2_REG1_REG_3__SCAN_IN;
  assign n12833 = ~n11677 | ~P2_REG0_REG_3__SCAN_IN;
  assign n12840 = ~n12834 | ~n12833;
  assign n12835 = ~P2_REG3_REG_3__SCAN_IN;
  assign n12838 = ~n11680 | ~n12835;
  assign n12836 = ~P2_REG2_REG_3__SCAN_IN;
  assign n12837 = n12883 | n12836;
  assign n12851 = ~n19167 | ~n12841;
  assign n16978 = ~n12842 ^ P2_IR_REG_3__SCAN_IN;
  assign n12843 = ~n16978;
  assign n12844 = n16826 | n12843;
  assign n13271 = ~n12899;
  assign n19056 = ~n12847 ^ n12846;
  assign n12848 = n13271 | n19056;
  assign n12850 = ~n19083 | ~n13114;
  assign n12881 = ~n12851 | ~n12850;
  assign n12852 = ~n12881 | ~n19100;
  assign n12854 = ~n12853 | ~n19078;
  assign n12856 = n12854 & n13114;
  assign n12871 = n18880 & n18756;
  assign n12855 = ~n12879 | ~n12871;
  assign n19187 = ~n19167;
  assign n12857 = ~n12881 | ~n19187;
  assign n12859 = ~n12811 | ~P2_REG3_REG_0__SCAN_IN;
  assign n12858 = ~n11677 | ~P2_REG0_REG_0__SCAN_IN;
  assign n12865 = ~n12859 | ~n12858;
  assign n12863 = ~n12860 | ~P2_REG1_REG_0__SCAN_IN;
  assign n12861 = ~P2_REG2_REG_0__SCAN_IN;
  assign n12862 = n12883 | n12861;
  assign n12864 = ~n12863 | ~n12862;
  assign n12868 = n16826 | n12866;
  assign n18684 = ~n13579 ^ P1_DATAO_REG_0__SCAN_IN;
  assign n12867 = ~n16826 | ~n18684;
  assign n18735 = ~n12868 | ~n12867;
  assign n18671 = ~n15691 | ~n18735;
  assign n12873 = ~n18671 & ~n12869;
  assign n15750 = ~n12870;
  assign n12872 = ~n12871;
  assign n12878 = ~n12873 & ~n18739;
  assign n18730 = ~n15691;
  assign n18667 = ~n18730 | ~n11929;
  assign n12877 = n18667 | n12841;
  assign n12874 = ~n15739;
  assign n12875 = n12874 | n15113;
  assign n12876 = ~n18667 | ~n12875;
  assign n12880 = n19187 & n19100;
  assign n12902 = ~n12881 & ~n12880;
  assign n12885 = ~n13159 | ~P2_REG0_REG_4__SCAN_IN;
  assign n12882 = ~P2_REG2_REG_4__SCAN_IN;
  assign n12884 = n12883 | n12882;
  assign n12890 = ~n12885 | ~n12884;
  assign n19210 = P2_REG3_REG_4__SCAN_IN ^ P2_REG3_REG_3__SCAN_IN;
  assign n12888 = ~n11680 | ~n19210;
  assign n12887 = ~n12860 | ~P2_REG1_REG_4__SCAN_IN;
  assign n12889 = ~n12888 | ~n12887;
  assign n12894 = ~n12891 | ~P2_IR_REG_4__SCAN_IN;
  assign n12893 = ~n12892 | ~P2_IR_REG_31__SCAN_IN;
  assign n12895 = ~n12894 | ~n12893;
  assign n19225 = ~n12895 | ~n12916;
  assign n12896 = n16826 | n19225;
  assign n14458 = ~n19277;
  assign n12900 = ~n12899 | ~n14458;
  assign n12930 = ~n19333 | ~n19193;
  assign n19351 = ~n19333;
  assign n12903 = ~n12902 & ~n19201;
  assign n12927 = ~n12904 | ~n12903;
  assign n12906 = ~n12860 | ~P2_REG1_REG_5__SCAN_IN;
  assign n12905 = ~n11677 | ~P2_REG0_REG_5__SCAN_IN;
  assign n12913 = n12906 & n12905;
  assign n12907 = ~P2_REG3_REG_5__SCAN_IN;
  assign n19370 = ~n12908 ^ n12907;
  assign n12911 = ~n11680 | ~n19370;
  assign n12909 = ~P2_REG2_REG_5__SCAN_IN;
  assign n12910 = n12883 | n12909;
  assign n12912 = n12911 & n12910;
  assign n19567 = ~n12913 | ~n12912;
  assign n19438 = ~n12915 ^ n12914;
  assign n14478 = ~n19438;
  assign n12924 = ~n14478 | ~n13257;
  assign n12917 = ~n12916 | ~P2_IR_REG_31__SCAN_IN;
  assign n12919 = ~n12917 | ~P2_IR_REG_5__SCAN_IN;
  assign n12918 = ~n12600 | ~P2_IR_REG_31__SCAN_IN;
  assign n12920 = ~n12919 | ~n12918;
  assign n17022 = n12920 & n12961;
  assign n16996 = ~n17022;
  assign n12921 = n16826 | n16996;
  assign n12923 = n12922 & n12921;
  assign n15755 = ~n19567 | ~n19373;
  assign n12925 = ~n15755 | ~n19346;
  assign n12926 = ~n12925 | ~n13114;
  assign n12929 = ~n12927 | ~n12926;
  assign n12928 = ~n19567;
  assign n15757 = ~n12928 | ~n19357;
  assign n12933 = ~n12929 | ~n15757;
  assign n12931 = ~n15757 | ~n12930;
  assign n12932 = ~n12931 | ~n12841;
  assign n12935 = ~n12933 | ~n12932;
  assign n12934 = n15755 | n13114;
  assign n12937 = ~n12860 | ~P2_REG1_REG_6__SCAN_IN;
  assign n12936 = ~n11677 | ~P2_REG0_REG_6__SCAN_IN;
  assign n12942 = ~n12937 | ~n12936;
  assign n19593 = ~n12938 ^ P2_REG3_REG_6__SCAN_IN;
  assign n12940 = ~n11680 | ~n19593;
  assign n19590 = ~P2_REG2_REG_6__SCAN_IN;
  assign n12939 = n12883 | n19590;
  assign n12941 = ~n12940 | ~n12939;
  assign n15701 = ~n12942 & ~n12941;
  assign n19547 = ~n12944 ^ n12943;
  assign n12949 = n19547 | n13271;
  assign n12946 = ~n12961 | ~P2_IR_REG_31__SCAN_IN;
  assign n17021 = ~n12946 ^ n12945;
  assign n12947 = ~n16826 & ~n17021;
  assign n12948 = ~n11697 & ~n12947;
  assign n19575 = ~n12949 | ~n12948;
  assign n15760 = ~n15701 | ~n19575;
  assign n19589 = ~n19575;
  assign n19670 = ~n15701;
  assign n15759 = ~n19589 | ~n19670;
  assign n19572 = n15760 & n15759;
  assign n19691 = P2_REG3_REG_7__SCAN_IN ^ n12950;
  assign n12952 = ~n11680 | ~n19691;
  assign n12951 = ~n11677 | ~P2_REG0_REG_7__SCAN_IN;
  assign n12957 = n12952 & n12951;
  assign n12955 = ~n12860 | ~P2_REG1_REG_7__SCAN_IN;
  assign n12953 = ~P2_REG2_REG_7__SCAN_IN;
  assign n12954 = n12883 | n12953;
  assign n12956 = n12955 & n12954;
  assign n19886 = ~n12957 | ~n12956;
  assign n19556 = ~n19886;
  assign n12959 = ~n12958;
  assign n19756 = ~n12960 ^ n12959;
  assign n12967 = n19756 | n13271;
  assign n12962 = n12961 | P2_IR_REG_6__SCAN_IN;
  assign n12963 = ~n12962 | ~P2_IR_REG_31__SCAN_IN;
  assign n17063 = ~n12963 ^ P2_IR_REG_7__SCAN_IN;
  assign n17037 = ~n17063;
  assign n12964 = n16826 | n17037;
  assign n12966 = n12965 & n12964;
  assign n12968 = n19572 & n13434;
  assign n15762 = ~n13434;
  assign n13433 = ~n19556 | ~n19696;
  assign n12969 = ~n13433 | ~n15760;
  assign n12970 = ~n12969 | ~n13114;
  assign n12971 = n15762 | n12970;
  assign n12972 = ~n13434 | ~n15759;
  assign n12973 = ~n12972 | ~n12841;
  assign n12974 = ~n19886 & ~n13395;
  assign n12975 = ~n12974 | ~n19696;
  assign n13005 = ~n12976 | ~n12975;
  assign n19913 = ~P2_REG3_REG_8__SCAN_IN ^ n12977;
  assign n12979 = ~n11680 | ~n19913;
  assign n12978 = ~n12860 | ~P2_REG1_REG_8__SCAN_IN;
  assign n12983 = n12979 & n12978;
  assign n12981 = ~n11677 | ~P2_REG0_REG_8__SCAN_IN;
  assign n19910 = ~P2_REG2_REG_8__SCAN_IN;
  assign n12980 = n12883 | n19910;
  assign n12982 = n12981 & n12980;
  assign n20059 = ~n12983 | ~n12982;
  assign n12999 = ~n20059 | ~n13293;
  assign n12998 = ~n12984 | ~n13293;
  assign n12986 = ~n12985;
  assign n19864 = ~n12987 ^ n12986;
  assign n12997 = n19864 | n13271;
  assign n12989 = n12988 | n12640;
  assign n12992 = ~n12989 | ~P2_IR_REG_8__SCAN_IN;
  assign n12991 = ~n12990 | ~P2_IR_REG_31__SCAN_IN;
  assign n12993 = ~n12992 | ~n12991;
  assign n19865 = ~n12993 | ~n13009;
  assign n12994 = n16826 | n19865;
  assign n12996 = n12995 & n12994;
  assign n19897 = ~n19909;
  assign n13003 = ~n12998 | ~n19897;
  assign n13004 = n20059 & n13114;
  assign n13000 = n13005 | n13004;
  assign n13001 = ~n13000 | ~n12999;
  assign n13002 = ~n13001 | ~n19909;
  assign n13032 = ~n13003 | ~n13002;
  assign n13030 = ~n13005 | ~n13004;
  assign n20035 = ~n13007 ^ n13006;
  assign n14539 = ~n20035;
  assign n13018 = ~n14539 | ~n13257;
  assign n13008 = ~P1_DATAO_REG_9__SCAN_IN;
  assign n13016 = n11671 | n13008;
  assign n13010 = ~n13009 | ~P2_IR_REG_31__SCAN_IN;
  assign n13013 = ~n13010 | ~P2_IR_REG_9__SCAN_IN;
  assign n13011 = ~P2_IR_REG_9__SCAN_IN;
  assign n13012 = ~n13011 | ~P2_IR_REG_31__SCAN_IN;
  assign n13014 = ~n13013 | ~n13012;
  assign n17288 = n13037 & n13014;
  assign n17086 = ~n17288;
  assign n13015 = n16826 | n17086;
  assign n13017 = n13016 & n13015;
  assign n13028 = ~n20081 | ~n13395;
  assign n20078 = P2_REG3_REG_9__SCAN_IN ^ n13019;
  assign n13021 = ~n11680 | ~n20078;
  assign n13020 = ~n12860 | ~P2_REG1_REG_9__SCAN_IN;
  assign n13026 = n13021 & n13020;
  assign n13024 = ~n11677 | ~P2_REG0_REG_9__SCAN_IN;
  assign n13022 = ~P2_REG2_REG_9__SCAN_IN;
  assign n13023 = n12883 | n13022;
  assign n13025 = n13024 & n13023;
  assign n20221 = ~n13026 | ~n13025;
  assign n13027 = n20221 | n13114;
  assign n13034 = ~n13028 | ~n13027;
  assign n19870 = ~n20221;
  assign n15707 = ~n20081 | ~n19870;
  assign n13029 = ~n13034 | ~n15707;
  assign n13031 = n13030 & n13029;
  assign n13065 = ~n13032 | ~n13031;
  assign n13033 = ~n20081 & ~n19870;
  assign n13062 = n13034 | n13033;
  assign n13056 = ~n13065 | ~n13062;
  assign n20196 = n13036 ^ n13035;
  assign n14558 = ~n20196;
  assign n13045 = ~n14558 | ~n13257;
  assign n13043 = n11671 | n20195;
  assign n13038 = ~n13037 | ~P2_IR_REG_31__SCAN_IN;
  assign n13040 = ~n13038 | ~P2_IR_REG_10__SCAN_IN;
  assign n13039 = ~n12602 | ~P2_IR_REG_31__SCAN_IN;
  assign n13041 = ~n13040 | ~n13039;
  assign n17267 = n13041 & n13071;
  assign n17089 = ~n17267;
  assign n13042 = n16826 | n17089;
  assign n13044 = n13043 & n13042;
  assign n13055 = ~n20243 | ~n13395;
  assign n13047 = ~n12860 | ~P2_REG1_REG_10__SCAN_IN;
  assign n13046 = ~n11677 | ~P2_REG0_REG_10__SCAN_IN;
  assign n13053 = n13047 & n13046;
  assign n20240 = ~P2_REG3_REG_10__SCAN_IN ^ n13048;
  assign n13051 = ~n11680 | ~n20240;
  assign n13049 = ~P2_REG2_REG_10__SCAN_IN;
  assign n13050 = n12883 | n13049;
  assign n13052 = n13051 & n13050;
  assign n20382 = ~n13053 | ~n13052;
  assign n13054 = n20382 | n13114;
  assign n13061 = n13055 & n13054;
  assign n13060 = ~n13056 | ~n13061;
  assign n20227 = ~n20243;
  assign n13058 = ~n20227 | ~n13293;
  assign n13057 = ~n20382 | ~n13395;
  assign n13059 = ~n13058 | ~n13057;
  assign n13067 = ~n13060 | ~n13059;
  assign n13063 = ~n13061;
  assign n13064 = n13063 & n13062;
  assign n13066 = ~n13065 | ~n13064;
  assign n13087 = ~n13067 | ~n13066;
  assign n20360 = n13069 ^ n13068;
  assign n14578 = ~n20360;
  assign n13075 = ~n14578 | ~n13257;
  assign n13070 = ~P1_DATAO_REG_11__SCAN_IN;
  assign n13073 = n11671 | n13070;
  assign n13096 = ~n13071 | ~P2_IR_REG_31__SCAN_IN;
  assign n17256 = ~n13096 ^ P2_IR_REG_11__SCAN_IN;
  assign n17082 = ~n17256;
  assign n13072 = n16826 | n17082;
  assign n13074 = n13073 & n13072;
  assign n13085 = n20409 | n12841;
  assign n20405 = P2_REG3_REG_11__SCAN_IN ^ n13076;
  assign n13078 = ~n11680 | ~n20405;
  assign n13077 = ~n11677 | ~P2_REG0_REG_11__SCAN_IN;
  assign n13083 = n13078 & n13077;
  assign n13081 = ~n12860 | ~P2_REG1_REG_11__SCAN_IN;
  assign n13079 = ~P2_REG2_REG_11__SCAN_IN;
  assign n13080 = n12883 | n13079;
  assign n13082 = n13081 & n13080;
  assign n20537 = ~n13083 | ~n13082;
  assign n13084 = n20537 | n13114;
  assign n13088 = ~n13085 | ~n13084;
  assign n15711 = n20409 | n20537;
  assign n13086 = n13088 & n15711;
  assign n13089 = ~n13088;
  assign n13436 = ~n20409 | ~n20537;
  assign n13090 = ~n13089 | ~n13436;
  assign n20519 = n13093 ^ n13092;
  assign n14601 = ~n20519;
  assign n13102 = ~n14601 | ~n13257;
  assign n13094 = ~P1_DATAO_REG_12__SCAN_IN;
  assign n13100 = n11671 | n13094;
  assign n13097 = n13096 & n13095;
  assign n13098 = ~n13097 & ~n12640;
  assign n17105 = ~P2_IR_REG_12__SCAN_IN ^ n13098;
  assign n13099 = n16826 | n17105;
  assign n13101 = n13100 & n13099;
  assign n20561 = ~n20545;
  assign n13111 = ~n13118 | ~n20561;
  assign n20558 = ~P2_REG3_REG_12__SCAN_IN ^ n13103;
  assign n13105 = ~n11680 | ~n20558;
  assign n13104 = ~n11677 | ~P2_REG0_REG_12__SCAN_IN;
  assign n13110 = n13105 & n13104;
  assign n13108 = ~n12860 | ~P2_REG1_REG_12__SCAN_IN;
  assign n13106 = ~P2_REG2_REG_12__SCAN_IN;
  assign n13107 = n12883 | n13106;
  assign n13109 = n13108 & n13107;
  assign n20702 = ~n13110 | ~n13109;
  assign n15773 = ~n20702;
  assign n13112 = ~n13111 | ~n15773;
  assign n13115 = ~n20702 | ~n13395;
  assign n13113 = ~n20545 | ~n13395;
  assign n13116 = ~n20545 | ~n13293;
  assign n13117 = n13116 & n13115;
  assign n13144 = ~n13120 | ~n13119;
  assign n13122 = ~n13121 | ~n13144;
  assign n15779 = ~n21198 | ~n21364;
  assign n21332 = n13124 ^ n13123;
  assign n14695 = ~n21332;
  assign n13132 = ~n14695 | ~n13257;
  assign n13125 = ~P1_DATAO_REG_17__SCAN_IN;
  assign n13130 = n11671 | n13125;
  assign n13153 = n13127 & n13126;
  assign n13128 = ~n13127 & ~n13126;
  assign n17196 = ~n13153 & ~n13128;
  assign n17154 = ~n17196;
  assign n13129 = n16826 | n17154;
  assign n13131 = n13130 & n13129;
  assign n21358 = n13132 & n13131;
  assign n13135 = ~n11677 | ~P2_REG0_REG_17__SCAN_IN;
  assign n13133 = ~P2_REG2_REG_17__SCAN_IN;
  assign n13134 = n12883 | n13133;
  assign n13137 = ~n13135 | ~n13134;
  assign n13136 = n12860 & P2_REG1_REG_17__SCAN_IN;
  assign n13140 = ~n13137 & ~n13136;
  assign n21352 = P2_REG3_REG_17__SCAN_IN ^ n13138;
  assign n13139 = ~n11680 | ~n21352;
  assign n21514 = ~n13140 | ~n13139;
  assign n13169 = ~n21358 | ~n21514;
  assign n13142 = ~n13141 | ~n13169;
  assign n13150 = ~n13142 | ~n13293;
  assign n13143 = n15779 & n15778;
  assign n13146 = ~n13144 | ~n13143;
  assign n13145 = ~n13421;
  assign n13147 = ~n13146 | ~n13145;
  assign n15781 = ~n21358 & ~n21514;
  assign n13148 = n13147 | n15781;
  assign n13149 = ~n13148 | ~n13395;
  assign n13174 = ~n13150 | ~n13149;
  assign n21491 = n13152 ^ n13151;
  assign n14345 = ~n21491;
  assign n13158 = ~n14345 | ~n13257;
  assign n13154 = ~n13153 & ~n12640;
  assign n17160 = ~P2_IR_REG_18__SCAN_IN ^ n13154;
  assign n13156 = ~n17160 & ~n16826;
  assign n13155 = ~n11671 & ~n21490;
  assign n13157 = ~n13156 & ~n13155;
  assign n13161 = ~n12860 | ~P2_REG1_REG_18__SCAN_IN;
  assign n13160 = ~n13159 | ~P2_REG0_REG_18__SCAN_IN;
  assign n13164 = ~n13161 | ~n13160;
  assign n13162 = ~P2_REG2_REG_18__SCAN_IN;
  assign n13163 = ~n12883 & ~n13162;
  assign n13167 = n13164 | n13163;
  assign n21533 = ~P2_REG3_REG_18__SCAN_IN ^ n13165;
  assign n13166 = n11680 & n21533;
  assign n21686 = n13167 | n13166;
  assign n15783 = n21536 | n21686;
  assign n13168 = ~n15781 & ~n13395;
  assign n13172 = ~n15783 | ~n13168;
  assign n13175 = ~n21536 | ~n21686;
  assign n13170 = n13169 & n13114;
  assign n13171 = ~n13175 | ~n13170;
  assign n13173 = ~n13172 | ~n13171;
  assign n13179 = ~n13174 | ~n13173;
  assign n13177 = ~n15783 | ~n13395;
  assign n13176 = ~n13175 | ~n13293;
  assign n13178 = ~n13177 | ~n13176;
  assign n13180 = ~n13179 | ~n13178;
  assign n13185 = ~n13182;
  assign n13184 = ~n13183;
  assign n13186 = ~n13185 & ~n13184;
  assign n13189 = ~n13187 & ~n12841;
  assign n13188 = ~n15787 & ~n13395;
  assign n22033 = n13191 ^ n13190;
  assign n13194 = ~n22033 | ~n13257;
  assign n13192 = ~P1_DATAO_REG_21__SCAN_IN;
  assign n13193 = n11671 | n13192;
  assign n13204 = ~n21950 & ~n13293;
  assign n13197 = ~n12860 | ~P2_REG1_REG_21__SCAN_IN;
  assign n13195 = ~P2_REG2_REG_21__SCAN_IN;
  assign n13196 = n12883 | n13195;
  assign n13199 = ~n13197 | ~n13196;
  assign n13198 = n11677 & P2_REG0_REG_21__SCAN_IN;
  assign n13202 = ~n13199 & ~n13198;
  assign n13220 = n13200 & P2_REG3_REG_20__SCAN_IN;
  assign n21961 = P2_REG3_REG_21__SCAN_IN ^ n13220;
  assign n13201 = ~n21961 | ~n11680;
  assign n22108 = ~n13202 | ~n13201;
  assign n13203 = ~n22108 & ~n13395;
  assign n13210 = ~n13204 & ~n13203;
  assign n13208 = ~n13209 & ~n13210;
  assign n13206 = ~n21950 & ~n13395;
  assign n13205 = ~n22108 & ~n13293;
  assign n13207 = ~n13206 & ~n13205;
  assign n13214 = ~n13208 & ~n13207;
  assign n13212 = ~n13209;
  assign n13211 = ~n13210;
  assign n13213 = ~n13212 & ~n13211;
  assign n13229 = ~n13214 & ~n13213;
  assign n22204 = n13216 ^ n13215;
  assign n13219 = ~n22204 | ~n13257;
  assign n13217 = ~P1_DATAO_REG_22__SCAN_IN;
  assign n13218 = n11671 | n13217;
  assign n13240 = n13220 & P2_REG3_REG_21__SCAN_IN;
  assign n22132 = P2_REG3_REG_22__SCAN_IN ^ n13240;
  assign n13227 = ~n22132 | ~n11680;
  assign n13223 = ~n11677 | ~P2_REG0_REG_22__SCAN_IN;
  assign n13221 = ~P2_REG2_REG_22__SCAN_IN;
  assign n13222 = n12883 | n13221;
  assign n13225 = ~n13223 | ~n13222;
  assign n13224 = n12860 & P2_REG1_REG_22__SCAN_IN;
  assign n13226 = ~n13225 & ~n13224;
  assign n22255 = ~n13227 | ~n13226;
  assign n13228 = ~n22115 | ~n22255;
  assign n15792 = ~n22255;
  assign n15732 = ~n22135 | ~n15792;
  assign n22122 = ~n13228 | ~n15732;
  assign n13234 = ~n13229 | ~n22122;
  assign n13231 = ~n22135 | ~n13395;
  assign n13230 = ~n15792 | ~n12841;
  assign n13232 = ~n13231 | ~n13230;
  assign n13233 = ~n13232 | ~n15732;
  assign n13249 = ~n13234 | ~n13233;
  assign n13239 = ~n22334 | ~n13257;
  assign n13237 = ~P1_DATAO_REG_23__SCAN_IN;
  assign n13238 = n11671 | n13237;
  assign n13261 = n13240 & P2_REG3_REG_22__SCAN_IN;
  assign n22239 = P2_REG3_REG_23__SCAN_IN ^ n13261;
  assign n13247 = ~n22239 | ~n11680;
  assign n13243 = ~n12860 | ~P2_REG1_REG_23__SCAN_IN;
  assign n13241 = ~P2_REG2_REG_23__SCAN_IN;
  assign n13242 = n12883 | n13241;
  assign n13245 = ~n13243 | ~n13242;
  assign n13244 = n11677 & P2_REG0_REG_23__SCAN_IN;
  assign n13246 = ~n13245 & ~n13244;
  assign n22381 = ~n13247 | ~n13246;
  assign n13248 = ~n22243 | ~n22381;
  assign n15795 = ~n22381;
  assign n15736 = ~n22268 | ~n15795;
  assign n15794 = ~n13248 | ~n15736;
  assign n13254 = ~n13249 | ~n15794;
  assign n13251 = ~n22268 | ~n13395;
  assign n13250 = ~n15795 | ~n12841;
  assign n13252 = ~n13251 | ~n13250;
  assign n13253 = ~n13252 | ~n15736;
  assign n13285 = ~n13254 | ~n13253;
  assign n13260 = ~n22473 | ~n13257;
  assign n13258 = ~P1_DATAO_REG_24__SCAN_IN;
  assign n13259 = n11671 | n13258;
  assign n13276 = ~n13261 | ~P2_REG3_REG_23__SCAN_IN;
  assign n22374 = ~P2_REG3_REG_24__SCAN_IN ^ n13276;
  assign n13268 = ~n22374 | ~n11680;
  assign n13264 = ~n12860 | ~P2_REG1_REG_24__SCAN_IN;
  assign n13262 = ~P2_REG2_REG_24__SCAN_IN;
  assign n13263 = n12883 | n13262;
  assign n13266 = ~n13264 | ~n13263;
  assign n13265 = n11677 & P2_REG0_REG_24__SCAN_IN;
  assign n13267 = ~n13266 & ~n13265;
  assign n22256 = ~n13268 | ~n13267;
  assign n13274 = ~n22559 | ~n13257;
  assign n13272 = ~P1_DATAO_REG_25__SCAN_IN;
  assign n13273 = n11671 | n13272;
  assign n13275 = ~P2_REG3_REG_24__SCAN_IN;
  assign n13303 = ~n13276 & ~n13275;
  assign n15843 = P2_REG3_REG_25__SCAN_IN ^ n13303;
  assign n13282 = ~n15843 | ~n11680;
  assign n13278 = ~n11677 | ~P2_REG0_REG_25__SCAN_IN;
  assign n15805 = ~P2_REG2_REG_25__SCAN_IN;
  assign n13277 = n12883 | n15805;
  assign n13280 = ~n13278 | ~n13277;
  assign n13279 = n12860 & P2_REG1_REG_25__SCAN_IN;
  assign n13281 = ~n13280 & ~n13279;
  assign n22382 = ~n13282 | ~n13281;
  assign n13283 = ~n15943 | ~n22382;
  assign n15942 = ~n22382;
  assign n13284 = n22389 & n15940;
  assign n13291 = ~n15940;
  assign n15354 = ~n22401;
  assign n13287 = ~n15354 | ~n13395;
  assign n15844 = ~n22256;
  assign n13286 = ~n15844 | ~n13293;
  assign n13289 = ~n13287 | ~n13286;
  assign n13288 = ~n15354 | ~n15844;
  assign n13290 = ~n13289 | ~n13288;
  assign n13292 = n13291 | n13290;
  assign n13295 = ~n15955 | ~n13395;
  assign n13294 = ~n15942 | ~n13293;
  assign n13296 = ~n13295 | ~n13294;
  assign n13297 = ~n13296 | ~n15966;
  assign n13302 = ~n22645 | ~n13257;
  assign n13300 = ~P1_DATAO_REG_26__SCAN_IN;
  assign n13301 = n11671 | n13300;
  assign n13324 = ~n13303 | ~P2_REG3_REG_25__SCAN_IN;
  assign n16042 = ~P2_REG3_REG_26__SCAN_IN ^ n13324;
  assign n13310 = ~n16042 | ~n11680;
  assign n13306 = ~n11677 | ~P2_REG0_REG_26__SCAN_IN;
  assign n13304 = ~P2_REG2_REG_26__SCAN_IN;
  assign n13305 = n12883 | n13304;
  assign n13308 = ~n13306 | ~n13305;
  assign n13307 = n12860 & P2_REG1_REG_26__SCAN_IN;
  assign n13309 = ~n13308 & ~n13307;
  assign n16883 = ~n13310 | ~n13309;
  assign n13312 = ~n15971 | ~n12869;
  assign n16161 = ~n16883;
  assign n13462 = ~n16039 | ~n16161;
  assign n13311 = ~n13462 | ~n13395;
  assign n13313 = ~n13312 | ~n13311;
  assign n13315 = ~n15971 | ~n13395;
  assign n13314 = ~n13462 | ~n12841;
  assign n13316 = ~n13315 | ~n13314;
  assign n13332 = ~n13317 | ~n13316;
  assign n13322 = ~n22739 | ~n13257;
  assign n13320 = ~P1_DATAO_REG_27__SCAN_IN;
  assign n13321 = n11671 | n13320;
  assign n13323 = ~P2_REG3_REG_26__SCAN_IN;
  assign n13338 = ~n13324 & ~n13323;
  assign n16162 = P2_REG3_REG_27__SCAN_IN ^ n13338;
  assign n13331 = ~n16162 | ~n11680;
  assign n13327 = ~n12860 | ~P2_REG1_REG_27__SCAN_IN;
  assign n13325 = ~P2_REG2_REG_27__SCAN_IN;
  assign n13326 = n12883 | n13325;
  assign n13329 = ~n13327 | ~n13326;
  assign n13328 = n13159 & P2_REG0_REG_27__SCAN_IN;
  assign n13330 = ~n13329 & ~n13328;
  assign n16886 = ~n13331 | ~n13330;
  assign n13354 = ~n13332 | ~n16128;
  assign n13335 = ~P1_DATAO_REG_28__SCAN_IN;
  assign n13336 = n11671 | n13335;
  assign n13367 = n13338 & P2_REG3_REG_27__SCAN_IN;
  assign n16718 = ~P2_REG3_REG_28__SCAN_IN ^ n13367;
  assign n13339 = ~n16718;
  assign n13345 = ~n13339 | ~n11680;
  assign n13341 = ~n12860 | ~P2_REG1_REG_28__SCAN_IN;
  assign n13340 = ~n11677 | ~P2_REG0_REG_28__SCAN_IN;
  assign n13343 = ~n13341 | ~n13340;
  assign n16125 = ~P2_REG2_REG_28__SCAN_IN;
  assign n13342 = ~n12883 & ~n16125;
  assign n13344 = ~n13343 & ~n13342;
  assign n16889 = ~n13345 | ~n13344;
  assign n13347 = ~n13357 & ~n13395;
  assign n16192 = ~n16889;
  assign n13355 = ~n16712 & ~n16192;
  assign n13346 = ~n13355 & ~n12841;
  assign n13352 = ~n13347 & ~n13346;
  assign n13349 = ~n16160 & ~n13395;
  assign n16118 = ~n16886;
  assign n13348 = ~n16118 & ~n12841;
  assign n13350 = ~n13349 & ~n13348;
  assign n13351 = ~n13350 & ~n16129;
  assign n13353 = ~n13352 & ~n13351;
  assign n13361 = ~n13354 | ~n13353;
  assign n13356 = ~n13355;
  assign n13359 = ~n13356 | ~n12841;
  assign n16187 = ~n13357;
  assign n13358 = ~n16187 | ~n13395;
  assign n13360 = ~n13359 | ~n13358;
  assign n13376 = ~n13361 | ~n13360;
  assign n13366 = ~n22784 | ~n12899;
  assign n13364 = ~P1_DATAO_REG_29__SCAN_IN;
  assign n13365 = n11671 | n13364;
  assign n16178 = ~n13367 | ~P2_REG3_REG_28__SCAN_IN;
  assign n13368 = ~n16178;
  assign n13375 = ~n13368 | ~n11680;
  assign n13370 = ~n12860 | ~P2_REG1_REG_29__SCAN_IN;
  assign n13369 = ~n13159 | ~P2_REG0_REG_29__SCAN_IN;
  assign n13373 = ~n13370 | ~n13369;
  assign n13371 = ~P2_REG2_REG_29__SCAN_IN;
  assign n13372 = ~n12883 & ~n13371;
  assign n13374 = ~n13373 & ~n13372;
  assign n16892 = ~n13375 | ~n13374;
  assign n13390 = ~n13394 & ~n16895;
  assign n13379 = ~SI_30_ | ~n13378;
  assign n13385 = ~n13380 | ~n13379;
  assign n13382 = ~n13554 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n13381 = ~n18818 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n13383 = ~n13382 | ~n13381;
  assign n13384 = ~n13383 ^ SI_31_;
  assign n13388 = ~n23453 | ~n13257;
  assign n13386 = ~P1_DATAO_REG_31__SCAN_IN;
  assign n13387 = n11671 | n13386;
  assign n13393 = ~n13390 & ~n13389;
  assign n13391 = ~n22812 & ~n16892;
  assign n13392 = ~n13400 | ~n13391;
  assign n13404 = ~n13393 | ~n13392;
  assign n13398 = ~n13394 & ~n22813;
  assign n13396 = ~n22913 | ~n22820;
  assign n13397 = ~n13396 | ~n13395;
  assign n13402 = ~n13398 & ~n13397;
  assign n16268 = ~n22812;
  assign n16717 = ~n16892;
  assign n13399 = ~n16268 & ~n16717;
  assign n13403 = ~n13402 | ~n13401;
  assign n13406 = ~n16899 | ~n13395;
  assign n13410 = ~n13407 | ~n13406;
  assign n13408 = ~n22820 | ~n13293;
  assign n13409 = ~n22913 | ~n13408;
  assign n13411 = ~n13410 | ~n13409;
  assign n13471 = ~n13477 | ~n21822;
  assign n13413 = ~n22820 ^ n22913;
  assign n13412 = ~n16194 ^ n22813;
  assign n13469 = ~n13413 & ~n13412;
  assign n13414 = ~n22108;
  assign n13415 = ~n21950 | ~n13414;
  assign n15790 = ~n21964 | ~n22108;
  assign n22118 = ~n13415 | ~n15790;
  assign n13417 = ~n21815 | ~n21939;
  assign n15730 = ~n21794 | ~n13416;
  assign n21797 = ~n13417 | ~n15730;
  assign n15776 = ~n15777 | ~n13418;
  assign n13420 = ~n15778;
  assign n13422 = ~n15779;
  assign n15752 = ~n15689 | ~n18900;
  assign n13423 = n18900 | n15689;
  assign n19087 = ~n15752 | ~n13423;
  assign n13425 = ~n19087 & ~n18739;
  assign n15753 = ~n19167 | ~n19100;
  assign n13424 = n19100 | n19167;
  assign n19196 = ~n15753 | ~n13424;
  assign n19091 = ~n19196;
  assign n13426 = ~n13425 | ~n19091;
  assign n13427 = ~n13426 & ~n19201;
  assign n19360 = n15757 & n15755;
  assign n13429 = ~n13427 | ~n19360;
  assign n13428 = ~n19572;
  assign n13431 = ~n13429 & ~n13428;
  assign n15766 = n20243 & n20382;
  assign n13430 = ~n20243 & ~n20382;
  assign n20230 = ~n15766 & ~n13430;
  assign n13443 = ~n13431 | ~n20230;
  assign n20045 = ~n20059;
  assign n15705 = ~n19909 | ~n20045;
  assign n13432 = n19909 | n20045;
  assign n19678 = ~n13434 | ~n13433;
  assign n13435 = ~n19678;
  assign n13439 = ~n19889 | ~n13435;
  assign n20391 = ~n15711 | ~n13436;
  assign n18728 = ~n18671;
  assign n13437 = ~n18667;
  assign n15120 = ~n18728 & ~n13437;
  assign n13438 = ~n20391 | ~n15120;
  assign n13441 = ~n13439 & ~n13438;
  assign n13440 = n20081 | n20221;
  assign n15765 = ~n20081 | ~n20221;
  assign n13442 = ~n13441 | ~n20068;
  assign n13446 = ~n13443 & ~n13442;
  assign n13444 = n20724 | n20874;
  assign n15775 = ~n20724 | ~n20874;
  assign n20712 = ~n13444 | ~n15775;
  assign n20549 = ~n20545 ^ n15773;
  assign n13445 = ~n20712 & ~n20549;
  assign n13447 = ~n13446 | ~n13445;
  assign n13448 = ~n15748 & ~n13447;
  assign n13449 = ~n21034 | ~n13448;
  assign n13451 = ~n15776 & ~n13449;
  assign n13450 = ~n21716 & ~n21788;
  assign n13455 = ~n13451 | ~n21696;
  assign n21376 = ~n21358;
  assign n13452 = ~n21376 | ~n21514;
  assign n21171 = ~n21514;
  assign n15725 = ~n21358 | ~n21171;
  assign n21361 = ~n13452 | ~n15725;
  assign n21664 = ~n21686;
  assign n13453 = n21536 | n21664;
  assign n15727 = ~n21536 | ~n21664;
  assign n21523 = ~n13453 | ~n15727;
  assign n13454 = ~n21361 | ~n21523;
  assign n13456 = ~n13455 & ~n13454;
  assign n13457 = ~n21797 | ~n13456;
  assign n13458 = ~n22118 & ~n13457;
  assign n13460 = ~n22122 | ~n13458;
  assign n13459 = ~n22389 | ~n15794;
  assign n13461 = ~n13460 & ~n13459;
  assign n13464 = ~n13461 | ~n15940;
  assign n13463 = ~n16185 | ~n15968;
  assign n13466 = ~n13464 & ~n13463;
  assign n15974 = ~n16128;
  assign n13465 = ~n15974 & ~n21822;
  assign n13467 = ~n13466 | ~n13465;
  assign n13468 = ~n13467 & ~n16189;
  assign n13470 = ~n13469 | ~n13468;
  assign n13472 = ~n15118;
  assign n15143 = ~n15126 | ~n15125;
  assign n13473 = ~n13472 | ~n15143;
  assign n13474 = ~n13477 | ~n13473;
  assign n13475 = ~n13474 | ~n15131;
  assign n13481 = ~n13477;
  assign n22148 = ~n15126;
  assign n13479 = ~n15739 | ~n22148;
  assign n13478 = ~n15125 | ~n21658;
  assign n13480 = ~n13479 | ~n13478;
  assign n13485 = ~n13484 | ~n13483;
  assign n13486 = ~n13485 | ~P2_IR_REG_31__SCAN_IN;
  assign n13496 = ~n13486 ^ P2_IR_REG_23__SCAN_IN;
  assign n14988 = ~n13496;
  assign n22925 = ~P2_STATE_REG_SCAN_IN;
  assign n22281 = ~n14988 & ~n22925;
  assign n13491 = n11815 | n12640;
  assign n13490 = ~P2_IR_REG_24__SCAN_IN;
  assign n13488 = n13491 & n13490;
  assign n13489 = ~n12640 & ~n13488;
  assign n22514 = ~n13489 ^ P2_IR_REG_25__SCAN_IN;
  assign n22415 = ~n13491 ^ n13490;
  assign n13494 = ~n22415;
  assign n13492 = ~P2_IR_REG_26__SCAN_IN;
  assign n22642 = ~n13493 ^ n13492;
  assign n15077 = ~n22642;
  assign n13495 = ~n13494 | ~n15077;
  assign n14989 = ~n22514 & ~n13495;
  assign n15150 = ~n13496 & ~n14989;
  assign n15818 = ~P2_STATE_REG_SCAN_IN | ~n15150;
  assign n16825 = ~n13496 & ~n15143;
  assign n15142 = n21822 & n21658;
  assign n13497 = ~n16825 | ~n15142;
  assign n15159 = ~n15818 & ~n13497;
  assign n15158 = ~n15159 | ~n16904;
  assign n13500 = ~n15158 & ~n11934;
  assign n13498 = ~n22281 | ~n22148;
  assign n13499 = ~n13498 | ~P2_B_REG_SCAN_IN;
  assign n20195 = ~P1_DATAO_REG_10__SCAN_IN;
  assign n21490 = ~P1_DATAO_REG_18__SCAN_IN;
  assign n15131 = ~n21658;
  assign keyinput_0 = 1'b1;
  assign keyinput_1 = 1'b1;
  assign keyinput_2 = 1'b0;
  assign keyinput_3 = 1'b1;
  assign keyinput_4 = 1'b1;
  assign keyinput_5 = 1'b0;
  assign keyinput_6 = 1'b1;
  assign keyinput_7 = 1'b1;
  assign keyinput_8 = 1'b0;
  assign keyinput_9 = 1'b0;
  assign keyinput_10 = 1'b0;
  assign keyinput_11 = 1'b1;
  assign keyinput_12 = 1'b0;
  assign keyinput_13 = 1'b0;
  assign keyinput_14 = 1'b0;
  assign keyinput_15 = 1'b0;
  assign keyinput_16 = 1'b0;
  assign keyinput_17 = 1'b1;
  assign keyinput_18 = 1'b1;
  assign keyinput_19 = 1'b0;
  assign keyinput_20 = 1'b1;
  assign keyinput_21 = 1'b1;
  assign keyinput_22 = 1'b0;
  assign keyinput_23 = 1'b0;
  assign keyinput_24 = 1'b0;
  assign keyinput_25 = 1'b1;
  assign keyinput_26 = 1'b1;
  assign keyinput_27 = 1'b1;
  assign keyinput_28 = 1'b0;
  assign keyinput_29 = 1'b0;
  assign keyinput_30 = 1'b0;
  assign keyinput_31 = 1'b1;
  assign keyinput_32 = 1'b0;
  assign keyinput_33 = 1'b1;
  assign keyinput_34 = 1'b1;
  assign keyinput_35 = 1'b0;
  assign keyinput_36 = 1'b1;
  assign keyinput_37 = 1'b1;
  assign keyinput_38 = 1'b0;
  assign keyinput_39 = 1'b1;
  assign keyinput_40 = 1'b0;
  assign keyinput_41 = 1'b1;
  assign keyinput_42 = 1'b0;
  assign keyinput_43 = 1'b1;
  assign keyinput_44 = 1'b0;
  assign keyinput_45 = 1'b1;
  assign keyinput_46 = 1'b0;
  assign keyinput_47 = 1'b0;
  assign keyinput_48 = 1'b1;
  assign keyinput_49 = 1'b0;
  assign keyinput_50 = 1'b1;
  assign keyinput_51 = 1'b0;
  assign keyinput_52 = 1'b1;
  assign keyinput_53 = 1'b1;
  assign keyinput_54 = 1'b1;
  assign keyinput_55 = 1'b1;
  assign keyinput_56 = 1'b0;
  assign keyinput_57 = 1'b1;
  assign keyinput_58 = 1'b0;
  assign keyinput_59 = 1'b1;
  assign keyinput_60 = 1'b0;
  assign keyinput_61 = 1'b1;
  assign keyinput_62 = 1'b0;
  assign keyinput_63 = 1'b0;
  assign keyinput_64 = 1'b0;
  assign keyinput_65 = 1'b0;
  assign keyinput_66 = 1'b0;
  assign keyinput_67 = 1'b1;
  assign keyinput_68 = 1'b1;
  assign keyinput_69 = 1'b1;
  assign keyinput_70 = 1'b0;
  assign keyinput_71 = 1'b0;
  assign keyinput_72 = 1'b0;
  assign keyinput_73 = 1'b1;
  assign keyinput_74 = 1'b0;
  assign keyinput_75 = 1'b0;
  assign keyinput_76 = 1'b1;
  assign keyinput_77 = 1'b0;
  assign keyinput_78 = 1'b0;
  assign keyinput_79 = 1'b0;
  assign keyinput_80 = 1'b1;
  assign keyinput_81 = 1'b1;
  assign keyinput_82 = 1'b1;
  assign keyinput_83 = 1'b0;
  assign keyinput_84 = 1'b0;
  assign keyinput_85 = 1'b0;
  assign keyinput_86 = 1'b0;
  assign keyinput_87 = 1'b0;
  assign keyinput_88 = 1'b0;
  assign keyinput_89 = 1'b0;
  assign keyinput_90 = 1'b0;
  assign keyinput_91 = 1'b0;
  assign keyinput_92 = 1'b0;
  assign keyinput_93 = 1'b0;
  assign keyinput_94 = 1'b1;
  assign keyinput_95 = 1'b0;
  assign keyinput_96 = 1'b0;
  assign keyinput_97 = 1'b1;
  assign keyinput_98 = 1'b1;
  assign keyinput_99 = 1'b0;
  assign keyinput_100 = 1'b0;
  assign keyinput_101 = 1'b1;
  assign keyinput_102 = 1'b0;
  assign keyinput_103 = 1'b0;
  assign keyinput_104 = 1'b0;
  assign keyinput_105 = 1'b1;
  assign keyinput_106 = 1'b0;
  assign keyinput_107 = 1'b1;
  assign keyinput_108 = 1'b0;
  assign keyinput_109 = 1'b0;
  assign keyinput_110 = 1'b1;
  assign keyinput_111 = 1'b1;
  assign keyinput_112 = 1'b1;
  assign keyinput_113 = 1'b0;
  assign keyinput_114 = 1'b0;
  assign keyinput_115 = 1'b0;
  assign keyinput_116 = 1'b1;
  assign keyinput_117 = 1'b1;
  assign keyinput_118 = 1'b0;
  assign keyinput_119 = 1'b1;
  assign keyinput_120 = 1'b1;
  assign keyinput_121 = 1'b0;
  assign keyinput_122 = 1'b1;
  assign keyinput_123 = 1'b1;
  assign keyinput_124 = 1'b1;
  assign keyinput_125 = 1'b1;
  assign keyinput_126 = 1'b1;
  assign keyinput_127 = 1'b0;
  assign keyinput_128 = 1'b0;
  assign keyinput_129 = 1'b1;
  assign keyinput_130 = 1'b0;
  assign keyinput_131 = 1'b0;
  assign keyinput_132 = 1'b1;
  assign keyinput_133 = 1'b1;
  assign keyinput_134 = 1'b1;
  assign keyinput_135 = 1'b1;
  assign keyinput_136 = 1'b1;
  assign keyinput_137 = 1'b0;
  assign keyinput_138 = 1'b1;
  assign keyinput_139 = 1'b1;
  assign keyinput_140 = 1'b1;
  assign keyinput_141 = 1'b0;
  assign keyinput_142 = 1'b0;
  assign keyinput_143 = 1'b0;
  assign keyinput_144 = 1'b0;
  assign keyinput_145 = 1'b1;
  assign keyinput_146 = 1'b1;
  assign keyinput_147 = 1'b0;
  assign keyinput_148 = 1'b1;
  assign keyinput_149 = 1'b0;
  assign keyinput_150 = 1'b0;
  assign keyinput_151 = 1'b0;
  assign keyinput_152 = 1'b0;
  assign keyinput_153 = 1'b0;
  assign keyinput_154 = 1'b0;
  assign keyinput_155 = 1'b0;
  assign keyinput_156 = 1'b0;
  assign keyinput_157 = 1'b0;
  assign keyinput_158 = 1'b0;
  assign keyinput_159 = 1'b0;
  assign input_0 = keyinput_0 ^ SI_31_;
  assign input_1 = keyinput_1 ^ SI_30_;
  assign AND_1 = input_0 & input_1;
  assign input_2 = keyinput_2 ^ SI_29_;
  assign AND_2 = input_2 & AND_1;
  assign input_3 = keyinput_3 ^ SI_28_;
  assign AND_3 = input_3 & AND_2;
  assign input_4 = keyinput_4 ^ SI_27_;
  assign OR_4 = input_4 | AND_3;
  assign input_5 = keyinput_5 ^ SI_26_;
  assign OR_5 = input_5 | OR_4;
  assign input_6 = keyinput_6 ^ SI_25_;
  assign AND_6 = input_6 & OR_5;
  assign input_7 = keyinput_7 ^ SI_24_;
  assign AND_7 = input_7 & AND_6;
  assign input_8 = keyinput_8 ^ SI_23_;
  assign AND_8 = input_8 & AND_7;
  assign input_9 = keyinput_9 ^ SI_22_;
  assign OR_9 = input_9 | AND_8;
  assign input_10 = keyinput_10 ^ SI_21_;
  assign OR_10 = input_10 | OR_9;
  assign input_11 = keyinput_11 ^ SI_20_;
  assign AND_11 = input_11 & OR_10;
  assign input_12 = keyinput_12 ^ SI_19_;
  assign OR_12 = input_12 | AND_11;
  assign input_13 = keyinput_13 ^ SI_18_;
  assign OR_13 = input_13 | OR_12;
  assign input_14 = keyinput_14 ^ SI_17_;
  assign AND_14 = input_14 & OR_13;
  assign input_15 = keyinput_15 ^ SI_16_;
  assign OR_15 = input_15 | AND_14;
  assign input_16 = keyinput_16 ^ SI_15_;
  assign OR_16 = input_16 | OR_15;
  assign input_17 = keyinput_17 ^ SI_14_;
  assign OR_17 = input_17 | OR_16;
  assign input_18 = keyinput_18 ^ SI_13_;
  assign OR_18 = input_18 | OR_17;
  assign input_19 = keyinput_19 ^ SI_12_;
  assign AND_19 = input_19 & OR_18;
  assign input_20 = keyinput_20 ^ SI_11_;
  assign AND_20 = input_20 & AND_19;
  assign input_21 = keyinput_21 ^ SI_10_;
  assign AND_21 = input_21 & AND_20;
  assign input_22 = keyinput_22 ^ SI_9_;
  assign OR_22 = input_22 | AND_21;
  assign input_23 = keyinput_23 ^ SI_8_;
  assign OR_23 = input_23 | OR_22;
  assign input_24 = keyinput_24 ^ SI_7_;
  assign AND_24 = input_24 & OR_23;
  assign input_25 = keyinput_25 ^ SI_6_;
  assign OR_25 = input_25 | AND_24;
  assign input_26 = keyinput_26 ^ SI_5_;
  assign OR_26 = input_26 | OR_25;
  assign input_27 = keyinput_27 ^ SI_4_;
  assign AND_27 = input_27 & OR_26;
  assign input_28 = keyinput_28 ^ SI_3_;
  assign OR_28 = input_28 | AND_27;
  assign input_29 = keyinput_29 ^ SI_2_;
  assign OR_29 = input_29 | OR_28;
  assign input_30 = keyinput_30 ^ SI_1_;
  assign OR_30 = input_30 | OR_29;
  assign input_31 = keyinput_31 ^ SI_0_;
  assign AND_31 = input_31 & OR_30;
  assign input_32 = keyinput_32 ^ P1_ADDR_REG_19__SCAN_IN;
  assign OR_32 = input_32 | AND_31;
  assign input_33 = keyinput_33 ^ P1_DATAO_REG_0__SCAN_IN;
  assign OR_33 = input_33 | OR_32;
  assign input_34 = keyinput_34 ^ P1_DATAO_REG_1__SCAN_IN;
  assign AND_34 = input_34 & OR_33;
  assign input_35 = keyinput_35 ^ P1_DATAO_REG_2__SCAN_IN;
  assign AND_35 = input_35 & AND_34;
  assign input_36 = keyinput_36 ^ P1_DATAO_REG_3__SCAN_IN;
  assign AND_36 = input_36 & AND_35;
  assign input_37 = keyinput_37 ^ P1_DATAO_REG_4__SCAN_IN;
  assign OR_37 = input_37 | AND_36;
  assign input_38 = keyinput_38 ^ P1_DATAO_REG_5__SCAN_IN;
  assign AND_38 = input_38 & OR_37;
  assign input_39 = keyinput_39 ^ P1_DATAO_REG_6__SCAN_IN;
  assign OR_39 = input_39 | AND_38;
  assign input_40 = keyinput_40 ^ P1_DATAO_REG_7__SCAN_IN;
  assign OR_40 = input_40 | OR_39;
  assign input_41 = keyinput_41 ^ P1_DATAO_REG_8__SCAN_IN;
  assign AND_41 = input_41 & OR_40;
  assign input_42 = keyinput_42 ^ P1_DATAO_REG_9__SCAN_IN;
  assign OR_42 = input_42 | AND_41;
  assign input_43 = keyinput_43 ^ P1_DATAO_REG_10__SCAN_IN;
  assign OR_43 = input_43 | OR_42;
  assign input_44 = keyinput_44 ^ P1_DATAO_REG_11__SCAN_IN;
  assign AND_44 = input_44 & OR_43;
  assign input_45 = keyinput_45 ^ P1_DATAO_REG_12__SCAN_IN;
  assign OR_45 = input_45 | AND_44;
  assign input_46 = keyinput_46 ^ P1_DATAO_REG_13__SCAN_IN;
  assign OR_46 = input_46 | OR_45;
  assign input_47 = keyinput_47 ^ P1_DATAO_REG_14__SCAN_IN;
  assign AND_47 = input_47 & OR_46;
  assign input_48 = keyinput_48 ^ P1_DATAO_REG_15__SCAN_IN;
  assign OR_48 = input_48 | AND_47;
  assign input_49 = keyinput_49 ^ P1_DATAO_REG_16__SCAN_IN;
  assign AND_49 = input_49 & OR_48;
  assign input_50 = keyinput_50 ^ P1_DATAO_REG_17__SCAN_IN;
  assign OR_50 = input_50 | AND_49;
  assign input_51 = keyinput_51 ^ P1_DATAO_REG_18__SCAN_IN;
  assign OR_51 = input_51 | OR_50;
  assign input_52 = keyinput_52 ^ P1_DATAO_REG_19__SCAN_IN;
  assign AND_52 = input_52 & OR_51;
  assign input_53 = keyinput_53 ^ P1_DATAO_REG_20__SCAN_IN;
  assign OR_53 = input_53 | AND_52;
  assign input_54 = keyinput_54 ^ P1_DATAO_REG_21__SCAN_IN;
  assign OR_54 = input_54 | OR_53;
  assign input_55 = keyinput_55 ^ P1_DATAO_REG_22__SCAN_IN;
  assign OR_55 = input_55 | OR_54;
  assign input_56 = keyinput_56 ^ P1_DATAO_REG_23__SCAN_IN;
  assign AND_56 = input_56 & OR_55;
  assign input_57 = keyinput_57 ^ P1_DATAO_REG_24__SCAN_IN;
  assign AND_57 = input_57 & AND_56;
  assign input_58 = keyinput_58 ^ P1_DATAO_REG_25__SCAN_IN;
  assign OR_58 = input_58 | AND_57;
  assign input_59 = keyinput_59 ^ P1_DATAO_REG_26__SCAN_IN;
  assign AND_59 = input_59 & OR_58;
  assign input_60 = keyinput_60 ^ P1_DATAO_REG_27__SCAN_IN;
  assign AND_60 = input_60 & AND_59;
  assign input_61 = keyinput_61 ^ P1_DATAO_REG_28__SCAN_IN;
  assign OR_61 = input_61 | AND_60;
  assign input_62 = keyinput_62 ^ P1_DATAO_REG_29__SCAN_IN;
  assign AND_62 = input_62 & OR_61;
  assign input_63 = keyinput_63 ^ P1_DATAO_REG_30__SCAN_IN;
  assign OR_63 = input_63 | AND_62;
  assign input_64 = keyinput_64 ^ P1_DATAO_REG_31__SCAN_IN;
  assign AND_64 = input_64 & OR_63;
  assign input_65 = keyinput_65 ^ P1_RD_REG_SCAN_IN;
  assign OR_65 = input_65 | AND_64;
  assign input_66 = keyinput_66 ^ P2_IR_REG_0__SCAN_IN;
  assign OR_66 = input_66 | OR_65;
  assign input_67 = keyinput_67 ^ P2_IR_REG_1__SCAN_IN;
  assign AND_67 = input_67 & OR_66;
  assign input_68 = keyinput_68 ^ P2_IR_REG_2__SCAN_IN;
  assign OR_68 = input_68 | AND_67;
  assign input_69 = keyinput_69 ^ P2_IR_REG_3__SCAN_IN;
  assign AND_69 = input_69 & OR_68;
  assign input_70 = keyinput_70 ^ P2_IR_REG_4__SCAN_IN;
  assign AND_70 = input_70 & AND_69;
  assign input_71 = keyinput_71 ^ P2_IR_REG_5__SCAN_IN;
  assign AND_71 = input_71 & AND_70;
  assign input_72 = keyinput_72 ^ P2_IR_REG_6__SCAN_IN;
  assign OR_72 = input_72 | AND_71;
  assign input_73 = keyinput_73 ^ P2_IR_REG_7__SCAN_IN;
  assign AND_73 = input_73 & OR_72;
  assign input_74 = keyinput_74 ^ P2_IR_REG_8__SCAN_IN;
  assign OR_74 = input_74 | AND_73;
  assign input_75 = keyinput_75 ^ P2_IR_REG_9__SCAN_IN;
  assign OR_75 = input_75 | OR_74;
  assign input_76 = keyinput_76 ^ P2_IR_REG_10__SCAN_IN;
  assign AND_76 = input_76 & OR_75;
  assign input_77 = keyinput_77 ^ P2_IR_REG_11__SCAN_IN;
  assign AND_77 = input_77 & AND_76;
  assign input_78 = keyinput_78 ^ P2_IR_REG_12__SCAN_IN;
  assign AND_78 = input_78 & AND_77;
  assign input_79 = keyinput_79 ^ P2_IR_REG_13__SCAN_IN;
  assign OR_79 = input_79 | AND_78;
  assign input_80 = keyinput_80 ^ SI_31_;
  assign input_81 = keyinput_81 ^ SI_30_;
  assign AND_81 = input_80 & input_81;
  assign input_82 = keyinput_82 ^ SI_29_;
  assign AND_82 = input_82 & AND_81;
  assign input_83 = keyinput_83 ^ SI_28_;
  assign AND_83 = input_83 & AND_82;
  assign input_84 = keyinput_84 ^ SI_27_;
  assign OR_84 = input_84 | AND_83;
  assign input_85 = keyinput_85 ^ SI_26_;
  assign OR_85 = input_85 | OR_84;
  assign input_86 = keyinput_86 ^ SI_25_;
  assign AND_86 = input_86 & OR_85;
  assign input_87 = keyinput_87 ^ SI_24_;
  assign AND_87 = input_87 & AND_86;
  assign input_88 = keyinput_88 ^ SI_23_;
  assign AND_88 = input_88 & AND_87;
  assign input_89 = keyinput_89 ^ SI_22_;
  assign OR_89 = input_89 | AND_88;
  assign input_90 = keyinput_90 ^ SI_21_;
  assign OR_90 = input_90 | OR_89;
  assign input_91 = keyinput_91 ^ SI_20_;
  assign AND_91 = input_91 & OR_90;
  assign input_92 = keyinput_92 ^ SI_19_;
  assign OR_92 = input_92 | AND_91;
  assign input_93 = keyinput_93 ^ SI_18_;
  assign OR_93 = input_93 | OR_92;
  assign input_94 = keyinput_94 ^ SI_17_;
  assign AND_94 = input_94 & OR_93;
  assign input_95 = keyinput_95 ^ SI_16_;
  assign OR_95 = input_95 | AND_94;
  assign input_96 = keyinput_96 ^ SI_15_;
  assign OR_96 = input_96 | OR_95;
  assign input_97 = keyinput_97 ^ SI_14_;
  assign OR_97 = input_97 | OR_96;
  assign input_98 = keyinput_98 ^ SI_13_;
  assign OR_98 = input_98 | OR_97;
  assign input_99 = keyinput_99 ^ SI_12_;
  assign AND_99 = input_99 & OR_98;
  assign input_100 = keyinput_100 ^ SI_11_;
  assign AND_100 = input_100 & AND_99;
  assign input_101 = keyinput_101 ^ SI_10_;
  assign AND_101 = input_101 & AND_100;
  assign input_102 = keyinput_102 ^ SI_9_;
  assign OR_102 = input_102 | AND_101;
  assign input_103 = keyinput_103 ^ SI_8_;
  assign OR_103 = input_103 | OR_102;
  assign input_104 = keyinput_104 ^ SI_7_;
  assign AND_104 = input_104 & OR_103;
  assign input_105 = keyinput_105 ^ SI_6_;
  assign OR_105 = input_105 | AND_104;
  assign input_106 = keyinput_106 ^ SI_5_;
  assign OR_106 = input_106 | OR_105;
  assign input_107 = keyinput_107 ^ SI_4_;
  assign AND_107 = input_107 & OR_106;
  assign input_108 = keyinput_108 ^ SI_3_;
  assign OR_108 = input_108 | AND_107;
  assign input_109 = keyinput_109 ^ SI_2_;
  assign OR_109 = input_109 | OR_108;
  assign input_110 = keyinput_110 ^ SI_1_;
  assign OR_110 = input_110 | OR_109;
  assign input_111 = keyinput_111 ^ SI_0_;
  assign AND_111 = input_111 & OR_110;
  assign input_112 = keyinput_112 ^ P1_ADDR_REG_19__SCAN_IN;
  assign OR_112 = input_112 | AND_111;
  assign input_113 = keyinput_113 ^ P1_DATAO_REG_0__SCAN_IN;
  assign OR_113 = input_113 | OR_112;
  assign input_114 = keyinput_114 ^ P1_DATAO_REG_1__SCAN_IN;
  assign AND_114 = input_114 & OR_113;
  assign input_115 = keyinput_115 ^ P1_DATAO_REG_2__SCAN_IN;
  assign AND_115 = input_115 & AND_114;
  assign input_116 = keyinput_116 ^ P1_DATAO_REG_3__SCAN_IN;
  assign AND_116 = input_116 & AND_115;
  assign input_117 = keyinput_117 ^ P1_DATAO_REG_4__SCAN_IN;
  assign OR_117 = input_117 | AND_116;
  assign input_118 = keyinput_118 ^ P1_DATAO_REG_5__SCAN_IN;
  assign AND_118 = input_118 & OR_117;
  assign input_119 = keyinput_119 ^ P1_DATAO_REG_6__SCAN_IN;
  assign OR_119 = input_119 | AND_118;
  assign input_120 = keyinput_120 ^ P1_DATAO_REG_7__SCAN_IN;
  assign OR_120 = input_120 | OR_119;
  assign input_121 = keyinput_121 ^ P1_DATAO_REG_8__SCAN_IN;
  assign AND_121 = input_121 & OR_120;
  assign input_122 = keyinput_122 ^ P1_DATAO_REG_9__SCAN_IN;
  assign OR_122 = input_122 | AND_121;
  assign input_123 = keyinput_123 ^ P1_DATAO_REG_10__SCAN_IN;
  assign OR_123 = input_123 | OR_122;
  assign input_124 = keyinput_124 ^ P1_DATAO_REG_11__SCAN_IN;
  assign AND_124 = input_124 & OR_123;
  assign input_125 = keyinput_125 ^ P1_DATAO_REG_12__SCAN_IN;
  assign OR_125 = input_125 | AND_124;
  assign input_126 = keyinput_126 ^ P1_DATAO_REG_13__SCAN_IN;
  assign OR_126 = input_126 | OR_125;
  assign input_127 = keyinput_127 ^ P1_DATAO_REG_14__SCAN_IN;
  assign AND_127 = input_127 & OR_126;
  assign input_128 = keyinput_128 ^ P1_DATAO_REG_15__SCAN_IN;
  assign OR_128 = input_128 | AND_127;
  assign input_129 = keyinput_129 ^ P1_DATAO_REG_16__SCAN_IN;
  assign AND_129 = input_129 & OR_128;
  assign input_130 = keyinput_130 ^ P1_DATAO_REG_17__SCAN_IN;
  assign OR_130 = input_130 | AND_129;
  assign input_131 = keyinput_131 ^ P1_DATAO_REG_18__SCAN_IN;
  assign OR_131 = input_131 | OR_130;
  assign input_132 = keyinput_132 ^ P1_DATAO_REG_19__SCAN_IN;
  assign AND_132 = input_132 & OR_131;
  assign input_133 = keyinput_133 ^ P1_DATAO_REG_20__SCAN_IN;
  assign OR_133 = input_133 | AND_132;
  assign input_134 = keyinput_134 ^ P1_DATAO_REG_21__SCAN_IN;
  assign OR_134 = input_134 | OR_133;
  assign input_135 = keyinput_135 ^ P1_DATAO_REG_22__SCAN_IN;
  assign OR_135 = input_135 | OR_134;
  assign input_136 = keyinput_136 ^ P1_DATAO_REG_23__SCAN_IN;
  assign AND_136 = input_136 & OR_135;
  assign input_137 = keyinput_137 ^ P1_DATAO_REG_24__SCAN_IN;
  assign AND_137 = input_137 & AND_136;
  assign input_138 = keyinput_138 ^ P1_DATAO_REG_25__SCAN_IN;
  assign OR_138 = input_138 | AND_137;
  assign input_139 = keyinput_139 ^ P1_DATAO_REG_26__SCAN_IN;
  assign AND_139 = input_139 & OR_138;
  assign input_140 = keyinput_140 ^ P1_DATAO_REG_27__SCAN_IN;
  assign AND_140 = input_140 & AND_139;
  assign input_141 = keyinput_141 ^ P1_DATAO_REG_28__SCAN_IN;
  assign OR_141 = input_141 | AND_140;
  assign input_142 = keyinput_142 ^ P1_DATAO_REG_29__SCAN_IN;
  assign AND_142 = input_142 & OR_141;
  assign input_143 = keyinput_143 ^ P1_DATAO_REG_30__SCAN_IN;
  assign OR_143 = input_143 | AND_142;
  assign input_144 = keyinput_144 ^ P1_DATAO_REG_31__SCAN_IN;
  assign AND_144 = input_144 & OR_143;
  assign input_145 = keyinput_145 ^ P1_RD_REG_SCAN_IN;
  assign OR_145 = input_145 | AND_144;
  assign input_146 = keyinput_146 ^ P2_IR_REG_0__SCAN_IN;
  assign OR_146 = input_146 | OR_145;
  assign input_147 = keyinput_147 ^ P2_IR_REG_1__SCAN_IN;
  assign AND_147 = input_147 & OR_146;
  assign input_148 = keyinput_148 ^ P2_IR_REG_2__SCAN_IN;
  assign OR_148 = input_148 | AND_147;
  assign input_149 = keyinput_149 ^ P2_IR_REG_3__SCAN_IN;
  assign AND_149 = input_149 & OR_148;
  assign input_150 = keyinput_150 ^ P2_IR_REG_4__SCAN_IN;
  assign AND_150 = input_150 & AND_149;
  assign input_151 = keyinput_151 ^ P2_IR_REG_5__SCAN_IN;
  assign AND_151 = input_151 & AND_150;
  assign input_152 = keyinput_152 ^ P2_IR_REG_6__SCAN_IN;
  assign OR_152 = input_152 | AND_151;
  assign input_153 = keyinput_153 ^ P2_IR_REG_7__SCAN_IN;
  assign AND_153 = input_153 & OR_152;
  assign input_154 = keyinput_154 ^ P2_IR_REG_8__SCAN_IN;
  assign OR_154 = input_154 | AND_153;
  assign input_155 = keyinput_155 ^ P2_IR_REG_9__SCAN_IN;
  assign OR_155 = input_155 | OR_154;
  assign input_156 = keyinput_156 ^ P2_IR_REG_10__SCAN_IN;
  assign AND_156 = input_156 & OR_155;
  assign input_157 = keyinput_157 ^ P2_IR_REG_11__SCAN_IN;
  assign AND_157 = input_157 & AND_156;
  assign input_158 = keyinput_158 ^ P2_IR_REG_12__SCAN_IN;
  assign AND_158 = input_158 & AND_157;
  assign input_159 = keyinput_159 ^ P2_IR_REG_13__SCAN_IN;
  assign OR_159 = input_159 | AND_158;
  assign OR_159_INV = ~OR_159;
  assign CASOP = OR_79 & OR_159_INV;
  assign P2_U3328 = P2_U3328_Lock ^ CASOP;
endmodule


