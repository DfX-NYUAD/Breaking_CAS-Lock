// Benchmark "b20_C" written by ABC on Thu Mar  5 01:04:56 2020

module b20_C ( 
    P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
    SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_,
    SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_,
    SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN,
    P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
    P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
    P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
    P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
    P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
    P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
    P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
    P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
    P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
    P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
    P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
    P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
    P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
    P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
    P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
    P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
    P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
    P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
    P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
    P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
    P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
    P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
    P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
    P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
    P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
    P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
    P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
    P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
    P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
    P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
    P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
    P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
    P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
    P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
    P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
    P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
    P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
    P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
    P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
    P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
    P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
    P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
    P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
    P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
    P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
    P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
    P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
    P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
    P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
    P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
    P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
    P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
    P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
    P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
    P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
    P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
    P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
    P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
    P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
    P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
    P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
    P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
    P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
    P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
    P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
    P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
    P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
    P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
    P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
    P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
    P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
    P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
    P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
    P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
    P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
    P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
    P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
    P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
    P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465,
    P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486,
    P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507,
    P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
    P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
    P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
    P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
    P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
    P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
    P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554,
    P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
    P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
    P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
    P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
    P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290,
    P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283,
    P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276,
    P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269,
    P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377,
    P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257,
    P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250,
    P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243,
    P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236,
    P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402,
    P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423,
    P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444,
    P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452,
    P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459,
    P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466,
    P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473,
    P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480,
    P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487,
    P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230,
    P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223,
    P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216,
    P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209,
    P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202,
    P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195,
    P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188,
    P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491,
    P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498,
    P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505,
    P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
    P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
    P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179,
    P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
    P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
    P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
    P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150,
    P2_U3893  );
  input  P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_,
    SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
    SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
    SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN,
    P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
    P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
    P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
    P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
    P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
    P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
    P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
    P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
    P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
    P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
    P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
    P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
    P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
    P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
    P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
    P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
    P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
    P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
    P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
    P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
    P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
    P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
    P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
    P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
    P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
    P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
    P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
    P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
    P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
    P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
    P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
    P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
    P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
    P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
    P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
    P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
    P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
    P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
    P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
    P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
    P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
    P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
    P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
    P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
    P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
    P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
    P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
    P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
    P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
    P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
    P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
    P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
    P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
    P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
    P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
    P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
    P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
    P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
    P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
    P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
    P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
    P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
    P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
    P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
    P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
    P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
    P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
    P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
    P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
    P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
    P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
    P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
    P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
    P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
    P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
    P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
    P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
    P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
    P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465,
    P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486,
    P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507,
    P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
    P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
    P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
    P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
    P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
    P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
    P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554,
    P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
    P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
    P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
    P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
    P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290,
    P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283,
    P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276,
    P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269,
    P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377,
    P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257,
    P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250,
    P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243,
    P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236,
    P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402,
    P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423,
    P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444,
    P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452,
    P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459,
    P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466,
    P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473,
    P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480,
    P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487,
    P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230,
    P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223,
    P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216,
    P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209,
    P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202,
    P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195,
    P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188,
    P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491,
    P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498,
    P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505,
    P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
    P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
    P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179,
    P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
    P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
    P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
    P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150,
    P2_U3893;
  wire n10912, n16383, n16378, n15414, n15532, n16419, n16358, n15323,
    n15670, n10299, n13348, n16702, n9283, n15388, n9325, n9001, n11910,
    n9343, n10218, n16149, n8932, n8931, n14970, n9347, n9087, n9053,
    n8919, n9493, n9043, n13718, n10624, n13314, n10280, n15674, n9770,
    n8950, n8933, n16453, n9012, n10297, n10904, n10906, n11382, n15429,
    n10806, n14900, n15602, n15338, n16936, n15240, n16442, n16438, n10958,
    n15516, n15999, n13672, n9024, n10963, n8924, n8928, n10714, n9810,
    n10969, n9430, n16045, n14804, n8918, n14149, n9957, n16446, n16441,
    n16430, n16222, n16421, n16352, n16221, n16220, n15571, n16219, n15628,
    n16326, n16144, n16921, n16944, n16920, n16943, n16429, n16343, n15466,
    n16143, n15294, n16142, n16150, n16041, n16342, n15297, n15558, n16428,
    n15507, n15326, n15459, n15622, n15491, n14689, n16432, n16040, n16949,
    n14692, n15506, n16140, n16321, n15616, n15325, n16916, n16211, n15556,
    n15621, n16141, n15327, n15023, n16843, n16837, n16319, n16911, n16036,
    n15082, n16209, n16363, n15246, n15026, n16029, n16931, n16320, n15016,
    n14539, n16316, n15053, n16930, n16909, n16832, n15177, n14574, n14979,
    n16027, n14542, n15289, n15312, n16362, n15483, n16210, n15365, n16814,
    n16946, n15069, n16136, n10941, n15415, n15450, n14963, n14953, n16915,
    n16907, n15081, n15102, n16908, n16312, n16835, n16311, n16836, n16039,
    n15319, n16026, n10940, n15615, n15029, n14966, n15663, n15480, n14978,
    n14540, n15351, n14433, n14943, n16309, n16904, n16372, n16315, n16131,
    n15662, n16137, n14905, n15614, n10922, n15109, n15317, n15154, n10939,
    n14360, n16820, n16826, n16829, n15066, n16804, n15067, n16028, n14537,
    n16015, n16139, n10937, n15315, n14923, n15619, n16434, n15416, n15304,
    n14570, n14904, n15226, n15158, n10357, n14840, n14869, n14800, n16427,
    n14803, n14982, n16934, n16902, n14887, n14952, n16314, n14872, n15482,
    n14843, n15065, n15465, n14793, n15594, n14862, n15412, n15541, n16818,
    n16310, n16006, n14959, n15332, n15618, n16800, n16017, n15469, n15063,
    n14998, n14161, n14153, n16215, n15504, n15658, n14968, n14801, n10935,
    n15302, n14941, n10350, n15301, n14973, n15079, n15500, n15060, n14886,
    n16361, n10920, n15108, n10910, n10933, n10905, n14877, n16792, n14425,
    n15411, n15539, n16398, n16007, n10883, n16408, n16306, n16806, n15078,
    n16403, n10707, n14684, n15593, n14890, n16008, n14837, n16896, n16791,
    n14829, n14997, n14816, n15613, n15599, n15499, n15364, n15107, n15530,
    n15538, n15477, n10902, n10908, n15409, n15061, n14747, n14681, n15015,
    n14668, n14658, n15568, n10688, n16206, n10913, n16304, n15528, n15578,
    n15623, n16407, n16124, n16339, n16790, n14665, n10706, n14148, n15646,
    n14939, n16400, n14934, n15019, n10721, n15552, n15975, n15526, n15468,
    n14733, n14894, n15361, n15310, n15007, n10724, n15077, n14778, n14533,
    n15463, n14536, n14679, n16898, n14566, n15437, n13886, n13854, n16773,
    n15153, n10861, n14621, n16783, n14728, n15588, n15573, n14635, n14523,
    n14513, n14958, n14950, n15306, n14861, n14828, n14866, n15997, n14932,
    n16301, n16227, n14534, n10622, n14565, n14520, n14860, n14827, n14317,
    n14531, n15054, n15244, n14421, n13678, n14320, n14957, n15151, n14865,
    n9742, n14645, n15163, n13685, n14949, n15519, n15576, n10840, n14955,
    n14420, n14884, n15162, n10898, n15052, n10682, n14387, n10866, n14797,
    n15242, n14948, n14836, n14792, n14397, n10831, n14347, n14350, n14255,
    n10839, n10838, n10487, n14394, n15149, n13682, n14448, n16766, n14530,
    n15987, n14552, n14315, n14223, n15148, n14254, n14294, n14835, n14272,
    n14544, n14791, n14226, n15443, n10858, n15982, n13680, n14503, n14306,
    n15161, n10837, n10835, n14291, n14929, n15350, n14796, n15051, n10664,
    n10692, n10662, n16121, n16054, n15176, n10657, n14345, n14662, n14881,
    n14995, n15972, n10836, n14676, n15348, n15962, n13458, n14564, n14314,
    n10663, n14248, n14657, n14204, n14675, n10811, n15175, n14271, n13456,
    n9735, n15013, n15956, n14927, n15225, n15346, n14409, n14834, n14517,
    n14661, n15228, n14512, n14221, n14203, n14313, n14369, n14656, n15155,
    n13993, n15166, n14502, n13307, n10660, n14211, n15223, n14095, n16745,
    n16200, n14419, n14671, n14107, n14516, n14821, n14859, n14286, n14220,
    n15959, n9734, n10679, n14528, n14344, n14241, n13996, n16895, n14146,
    n14815, n15227, n16746, n14124, n15958, n14732, n16747, n14527, n15214,
    n15965, n14844, n14281, n13949, n15005, n14922, n16050, n14823, n15101,
    n13946, n14562, n14343, n14674, n15221, n13305, n13936, n14238, n14391,
    n14386, n15948, n14090, n14096, n13826, n14192, n14106, n13991, n14289,
    n13968, n13983, n14305, n14811, n10640, n10824, n14921, n14132, n10776,
    n15943, n14525, n14128, n14775, n14730, n14210, n13935, n13762, n13943,
    n13122, n14285, n14288, n14725, n14918, n10320, n14746, n14110, n13825,
    n14089, n14909, n14312, n14543, n16890, n14083, n16728, n15287, n14105,
    n14634, n13128, n14390, n13713, n13765, n14385, n13629, n13972, n10815,
    n13632, n16112, n10645, n14311, n14632, n13922, n14545, n15932, n15278,
    n16735, n14555, n13990, n10638, n10778, n14607, n14100, n16740, n14744,
    n10791, n14209, n13879, n13942, n15407, n13963, n13894, n14474, n14485,
    n10773, n15913, n14771, n14786, n14284, n14620, n13759, n14436, n14310,
    n13989, n13712, n10259, n14087, n14606, n10771, n15277, n14342, n10607,
    n10606, n15405, n14770, n13589, n13891, n13628, n13615, n13814, n13900,
    n13700, n13966, n10642, n13612, n13737, n13579, n13565, n14341, n15272,
    n13661, n13758, n14401, n13875, n13921, n13958, n14736, n14233, n13982,
    n10774, n15404, n14472, n16720, n14435, n15919, n13888, n13965, n13962,
    n14650, n14333, n13534, n10759, n14473, n13669, n10757, n14231, n15271,
    n15910, n14340, n12976, n13920, n13626, n14219, n13625, n14336, n14447,
    n14175, n13740, n13601, n13751, n15408, n14218, n13915, n15269, n13726,
    n13657, n16289, n15393, n13610, n10741, n15213, n14649, n13666, n13734,
    n16107, n16099, n16706, n13600, n13868, n13562, n13575, n10756, n13988,
    n10611, n10573, n13210, n14496, n10484, n15204, n13663, n13449, n10556,
    n15384, n10739, n15383, n13750, n13479, n10737, n13699, n15895, n9705,
    n10164, n13733, n16155, n14487, n14379, n16291, n14261, n13519, n13561,
    n10555, n13985, n14363, n14489, n13300, n15382, n10726, n14723, n15202,
    n15260, n14495, n10736, n10593, n13652, n13698, n13477, n13446, n14262,
    n10461, n14373, n14378, n14179, n15286, n13609, n15406, n13207, n15370,
    n16689, n14227, n13441, n13574, n13941, n14181, n15368, n13214, n13354,
    n13397, n13515, n9700, n15201, n13250, n13353, n10437, n10577, n13573,
    n13664, n13247, n13445, n13558, n15366, n13383, n10412, n14708, n15205,
    n15279, n14705, n13692, n13557, n14605, n10402, n15283, n13244, n13179,
    n10435, n10411, n10537, n15375, n10410, n10545, n13375, n13442, n13238,
    n13809, n13206, n16882, n14375, n13176, n13387, n10409, n13803, n15284,
    n15140, n9692, n10434, n15195, n10432, n10406, n10401, n14040, n15212,
    n13333, n15253, n13897, n14769, n13154, n13219, n13754, n15130, n16228,
    n13235, n10407, n14714, n10408, n13175, n16156, n13137, n13817, n14701,
    n15873, n13245, n13800, n13686, n13898, n12915, n10384, n13232, n15128,
    n14722, n16056, n14597, n13611, n14765, n12912, n10403, n14135, n9278,
    n15251, n14471, n16625, n14711, n13865, n10397, n13618, n14767, n14468,
    n16603, n14590, n13688, n10296, n13952, n14763, n10508, n12944, n13131,
    n12758, n13522, n15125, n10263, n15135, n14467, n13603, n10373, n16875,
    n13544, n14712, n14018, n10075, n13548, n10261, n13380, n16062, n16624,
    n10295, n15134, n13078, n15863, n10279, n13521, n15123, n10358, n10237,
    n16458, n15853, n14720, n16059, n10213, n10074, n14758, n13581, n10277,
    n16872, n14750, n13715, n10394, n13546, n14748, n14756, n13190, n13781,
    n10076, n13637, n10071, n13728, n13717, n10273, n16622, n15830, n13186,
    n13184, n13727, n16274, n12929, n13202, n14453, n10286, n16465, n10252,
    n14460, n16276, n16061, n13645, n13648, n14451, n9687, n13261, n15562,
    n14572, n14458, n14029, n10050, n16415, n10270, n15449, n13008, n10210,
    n10047, n10062, n12814, n16349, n14686, n13508, n10202, n16179, n14037,
    n13833, n16809, n15237, n16870, n13841, n9686, n13044, n13039, n10048,
    n10200, n12858, n10044, n16775, n16597, n16905, n16088, n13437, n13425,
    n15643, n16779, n13320, n10501, n16868, n12521, n15001, n9685, n15575,
    n13360, n13089, n15572, n13064, n13488, n10012, n10700, n9992, n16076,
    n16866, n12965, n13290, n13483, n12516, n13271, n13011, n16173, n15669,
    n13268, n12113, n12560, n9684, n13409, n14429, n13390, n15579, n15446,
    n9639, n13293, n10495, n16424, n13279, n16582, n15796, n12572, n9608,
    n14781, n15234, n12108, n12558, n16570, n9989, n9984, n16573, n9683,
    n12889, n15112, n15334, n16454, n16078, n10001, n12155, n16574, n10896,
    n12164, n13275, n15308, n16018, n13029, n12837, n12015, n16734, n12530,
    n12010, n10930, n12161, n15045, n12836, n12152, n15969, n16439, n15520,
    n15495, n15964, n16721, n10620, n14826, n10889, n10872, n10718, n11864,
    n10828, n16444, n12531, n11892, n9682, n16703, n10871, n10888, n16560,
    n11598, n11610, n10807, n9394, n11889, n15953, n12440, n9938, n11987,
    n15497, n11859, n11070, n12538, n15659, n14547, n10849, n15439, n11986,
    n11534, n15937, n16851, n15601, n16553, n10887, n14641, n16696, n11563,
    n11596, n12539, n12100, n11503, n15518, n9681, n12535, n10869, n10821,
    n16259, n11630, n15511, n11643, n11644, n15428, n15933, n15094, n16548,
    n12364, n15167, n11886, n11550, n9399, n11533, n11508, n11501, n15342,
    n9398, n11557, n16631, n11296, n12435, n14611, n9649, n11890, n11304,
    n12006, n16542, n10788, n15455, n15426, n9680, n10847, n11834, n11391,
    n11990, n11302, n15028, n12007, n11553, n11293, n14610, n11786, n9364,
    n16540, n16482, n16665, n9527, n11884, n13730, n10767, n14737, n10804,
    n9389, n13101, n13694, n10818, n13023, n16960, n15916, n16065, n11763,
    n12900, n11301, n15836, n11292, n9383, n9387, n13571, n9678, n14079,
    n15564, n12022, n11835, n11883, n11661, n15557, n15901, n11832, n11428,
    n11172, n12023, n16133, n11209, n11982, n11426, n16313, n13808, n10546,
    n14177, n15850, n10123, n13283, n10785, n12407, n11855, n11277, n15654,
    n10827, n10653, n10634, n10604, n10587, n10561, n10569, n10674, n10552,
    n10525, n10527, n10533, n10515, n10171, n10192, n10224, n9638, n10764,
    n11984, n14874, n11272, n15182, n9676, n11275, n11077, n11891, n10747,
    n16345, n10251, n13769, n10488, n11574, n10544, n15371, n9385, n11875,
    n10131, n11873, n13276, n10579, n10269, n10595, n10421, n11575, n16346,
    n10711, n11322, n16365, n10613, n10733, n9674, n10644, n10028, n15536,
    n10393, n13789, n11025, n11573, n10228, n8925, n10470, n11754, n10285,
    n10671, n13258, n9089, n11587, n16367, n8927, n10061, n11662, n9973,
    n15479, n15584, n10450, n10962, n11588, n10116, n11554, n16146, n11560,
    n12517, n11572, n13040, n12109, n9755, n10452, n12011, n11860, n9633,
    n11569, n10966, n11537, n10425, n11586, n10226, n9002, n9323, n14685,
    n12101, n10239, n9261, n9242, n9137, n10024, n9564, n10375, n9271,
    n9628, n9251, n11584, n12125, n9224, n10053, n16956, n9620, n9733,
    n9610, n9233, n9196, n12121, n9384, n9380, n10151, n10322, n9223,
    n9212, n9136, n11581, n9232, n11211, n9616, n12536, n10955, n11856,
    n9065, n11876, n9724, n9184, n9709, n9920, n9731, n9203, n9179, n9197,
    n9150, n9189, n9719, n9135, n10021, n9070, n9258, n9231, n9230, n9619,
    n9249, n10332, n9268, n9694, n9239, n9248, n10150, n9240, n10414,
    n9221, n10337, n9699, n9133, n9229, n9219, n9149, n9188, n10035, n9194,
    n9183, n9178, n11872, n9997, n9523, n9727, n9728, n9356, n9569, n9996,
    n9696, n14154, n13679, n9544, n9217, n9284, n9273, n9148, n11568,
    n9131, n13683, n11583, n9264, n10388, n11571, n10324, n9598, n9280,
    n13123, n10002, n9707, n9590, n9761, n9067, n9968, n9702, n9712, n9519,
    n9717, n9054, n9285, n9697, n9943, n9551, n9287, n9132, n9975, n11344,
    n9520, n9552, n9950, n9925, n9031, n9501, n9336, n9749, n9008, n8990,
    n8995, n8961, n9502, n9078, n10374, n10478, n10417, n8951, n10445,
    n9084, n10520, n10282, n10489, n14047, n10166, n9662, n8954, n8964,
    n9025, n9631, n9882, n9618, n9027, n8984, n8983, n8985, n9028, n9006,
    n11267, n16967, n16957, n16393, n16922, n16364, n16396, n15633, n16848,
    n15630, n16437, n15667, n15508, n15549, n15546, n16152, n16376, n15563,
    n16404, n15494, n15476, n16952, n16325, n15473, n15514, n16833, n16213,
    n15420, n16323, n15423, n15513, n15085, n15118, n15441, n16828, n16416,
    n15648, n15115, n15542, n15033, n15492, n15036, n15457, n16390, n15292,
    n15438, n15418, n15486, n16842, n14986, n16389, n14687, n16034, n14989,
    n15031, n14980, n15030, n15010, n15320, n15321, n16409, n16841, n16797,
    n16813, n15110, n16929, n15238, n16033, n16373, n16830, n16831, n14983,
    n14984, n15008, n15080, n14888, n15164, n14906, n16914, n15627, n16928,
    n15580, n16935, n15600, n15470, n16368, n15089, n15336, n14960, n10917,
    n16308, n16822, n16923, n14974, n16819, n16899, n10911, n10915, n16214,
    n15464, n15456, n14852, n16927, n10921, n14784, n16426, n15661, n14951,
    n16132, n14879, n16371, n16788, n15577, n16897, n15657, n14838, n15634,
    n16226, n14009, n15424, n16786, n15996, n15978, n14940, n14850, n16769,
    n16812, n15291, n16360, n14782, n16207, n10932, n10914, n15249, n14004,
    n14885, n15299, n15498, n15537, n15598, n16049, n10879, n15590, n16388,
    n10723, n14897, n15105, n14780, n15994, n15020, n16002, n15612, n15014,
    n16354, n14647, n15106, n14666, n15037, n14567, n15496, n16047, n15488,
    n10880, n10876, n15550, n15073, n13998, n15525, n15489, n15436, n15410,
    n15300, n10878, n10875, n14663, n16297, n14521, n14554, n10862, n15452,
    n14422, n14505, n15989, n14678, n16205, n14546, n15988, n14486, n16122,
    n14931, n16296, n14318, n13465, n14677, n10857, n15973, n14518, n10854,
    n15986, n15288, n15058, n16752, n14411, n14371, n14256, n14883, n14348,
    n15241, n15230, n14395, n15985, n16120, n10856, n14205, n10853, n16744,
    n14224, n14259, n14945, n15984, n14292, n14392, n14824, n14298, n14529,
    n14334, n10656, n10832, n10659, n16754, n15159, n15968, n16760, n15018,
    n16749, n16201, n14295, n10729, n10830, n16743, n16051, n14257, n14092,
    n15344, n14833, n14831, n14176, n13453, n10844, n14925, n10813, n16748,
    n13313, n14511, n14270, n14184, n15086, n14194, n10810, n14817, n13994,
    n16738, n14418, n14557, n14232, n15940, n14093, n10655, n14069, n14785,
    n15951, n14501, n15088, n10825, n16115, n13302, n13827, n15219, n14790,
    n14731, n10801, n15100, n13925, n14819, n14054, n14404, n14830, n10677,
    n14246, n13971, n14991, n15004, n13947, n14561, n14864, n14809, n15942,
    n13301, n15925, n14526, n13944, n14182, n15935, n13969, n14304, n14729,
    n16741, n15930, n10792, n14789, n13120, n14854, n16718, n13895, n13816,
    n10608, n13763, n13910, n13934, n13127, n16727, n14414, n16055, n16294,
    n15905, n13703, n13892, n14727, n13631, n14743, n14631, n13876, n9715,
    n14244, n16194, n16712, n13739, n14202, n16726, n13736, n13760, n13804,
    n13711, n13670, n14434, n10770, n13667, n10258, n14309, n14412, n14242,
    n12978, n14773, n15927, n14660, n10614, n10782, n15898, n13981, n13658,
    n15912, n13614, n16715, n13563, n14374, n13588, n13801, n16687, n15915,
    n10761, n14230, n16686, n14195, n16286, n13533, n15896, n10596, n14515,
    n16714, n16708, n16707, n14337, n16101, n13877, n10571, n13863, n13914,
    n13867, n13559, n13889, n10554, n12652, n14493, n14287, n10580, n14389,
    n10139, n14377, n15882, n10746, n14229, n14213, n14187, n15908, n13644,
    n10460, n14178, n13296, n10467, n16675, n13568, n14361, n14376, n13295,
    n13513, n13651, n10734, n15256, n15377, n10562, n13912, n10451, n13547,
    n15199, n13444, n13511, n14273, n16654, n13243, n12176, n15373, n10405,
    n13553, n13805, n10535, n15887, n15190, n10431, n14088, n10441, n13552,
    n13927, n14372, n14282, n16880, n14275, n13189, n13802, n14130, n14059,
    n13174, n10386, n14072, n15180, n10404, n10400, n15254, n13200, n10383,
    n13798, n10422, n13550, n14696, n13087, n13926, n16626, n16627, n14076,
    n15209, n16636, n10505, n10399, n16060, n16634, n13065, n12968, n16642,
    n13704, n10396, n16282, n16633, n13950, n14113, n14585, n13719, n13887,
    n13545, n14719, n16617, n10254, n13595, n10301, n13720, n14577, n16620,
    n16183, n13604, n10294, n14013, n10193, n12891, n10212, n10211, n13541,
    n13061, n10275, n13364, n16615, n16621, n12746, n10272, n14028, n16467,
    n16604, n16271, n14601, n13776, n12744, n15781, n10225, n10049, n13256,
    n13073, n16834, n13835, n13843, n15560, n12582, n14036, n15447, n13768,
    n10056, n12365, n9646, n13066, n12689, n15561, n15235, n10017, n13376,
    n13143, n13839, n10046, n13832, n13402, n10057, n12888, n10043, n13792,
    n13378, n16270, n16607, n13362, n9991, n13270, n16592, n16539, n12418,
    n16085, n16356, n16425, n13407, n9626, n10029, n10011, n13480, n9609,
    n9625, n13278, n12373, n15413, n16586, n12080, n16759, n12372, n12747,
    n16514, n12424, n15540, n12238, n13031, n13010, n9960, n10874, n10855,
    n9624, n10877, n10852, n15485, n15792, n12370, n10722, n16576, n12994,
    n15772, n12547, n16170, n12045, n16513, n11904, n16494, n12367, n13055,
    n12160, n16512, n14779, n9949, n13053, n11988, n9911, n15655, n12151,
    n12050, n11708, n15502, n12528, n11535, n15068, n11722, n14878, n16505,
    n10850, n9934, n9561, n9204, n15617, n11814, n15754, n9914, n9393,
    n15521, n16381, n9801, n16377, n15324, n16487, n12810, n16486, n9913,
    n15146, n12459, n12187, n9653, n12762, n16551, n14914, n16501, n12235,
    n12098, n16235, n11811, n12322, n9889, n11532, n12765, n12400, n11724,
    n10646, n11679, n9924, n12124, n10553, n13634, n12122, n15731, n11529,
    n12420, n11526, n12675, n11659, n9020, n14450, n11530, n13503, n15777,
    n13731, n12004, n16475, n16608, n16466, n13859, n15883, n12997, n10179,
    n13960, n13015, n10534, n12769, n15820, n10476, n12375, n15803, n14060,
    n15789, n14136, n15751, n15840, n15773, n11655, n10199, n11524, n9603,
    n11997, n16516, n10172, n9362, n9425, n16496, n9645, n9656, n13871,
    n9019, n9331, n9832, n15394, n11812, n10157, n10158, n16847, n11528,
    n11853, n12019, n10209, n9791, n10458, n10112, n16507, n11759, n10115,
    n11663, n9623, n9411, n9512, n9015, n11761, n10851, n10119, n10560,
    n10926, n10180, n10524, n15268, n15398, n10639, n10678, n10684, n10693,
    n10191, n10223, n11949, n10514, n10198, n10111, n9324, n10549, n16845,
    n10372, n9841, n11751, n10000, n15639, n10118, n14935, n10110, n11101,
    n11833, n10420, n9463, n13779, n10865, n10268, n9101, n15484, n10843,
    n16333, n9813, n8926, n9342, n8920, n10745, n15369, n10005, n14971,
    n10781, n10864, n14892, n9023, n10719, n10899, n10814, n10206, n9098,
    n13454, n14967, n9756, n15281, n10120, n10204, n15381, n9088, n10216,
    n10240, n10188, n10363, n8921, n9474, n9329, n9344, n14156, n9632,
    n9752, n15386, n13303, n14426, n8968, n8953, n10135, n9322, n9750,
    n9286, n10576, n9011, n9630, n9732, n8973, n8962, n14598, n13119,
    n9328, n14717, n16433, n9459, n9259, n9269, n10327, n9747, n9213,
    n9408, n8960, n10676, n9014, n9511, n10342, n9379, n9069, n9210,
    n10341, n8970, n9202, n16939, n10336, n9969, n9079, n8959, n9617,
    n14351, n9591, n14157, n9052, n9570, n9721, n9245, n9068, n9235, n9208,
    n9254, n9226, n9201, n9244, n14034, n16322, n9182, n10032, n9192,
    n9706, n9279, n10247, n9187, n9711, n9186, n9274, n9181, n9044, n9058,
    n9200, n9916, n9207, n9191, n9722, n9216, n9517, n10265, n9139, n9494,
    n10219, n8981, n9030, n9138, n9516, n8997, n9134, n9096, n8965, n8986,
    n8987, n8949, n9518, n8943, n9026, n8974, n9543, n8996, n9491, n9038,
    n9046, n9334, n9335, n9341, n9107, n8975, n8963, n9743, n8979, n9748,
    n9729, n10364, n16134, n16900, n13431, n8922, n16940, n9405, n11100,
    n8923, n16918, n16774, n16044, n8929, n8930, n10730, n16958, n10826,
    n9428, n9446, n15591, n9037, n9726, n9199, n15087, n13103, n10795,
    n10777, n13346, n9367, n9368, n9355, n16533, n16661, n11773, n10015,
    n9993, n9964, n9959, n11683, n9263, n9206, n14074, n10517, n10589,
    n9509, n9361, n11556, n12020, n10667, n10627, n13322, n10222, n9492,
    n10433, n10833, n9872, n12872, n10276, n10274, n10796, n10907, n14237,
    n13067, n10800, n9220, n9478, n9641, n14041, n9354, n10572, n9371,
    n10208, n9366, n13389, n13233, n9521, n10742, n10743, n15998, n9998,
    n15132, n16485, n16503, n16614, n15944, n16232, n16795, n9536, n9431,
    n10016, n10045, n9246, n10661, n10658, n10686, n10253, n16917, n9485,
    n9094, n9146, n9147, n12014, n12123, n13470, n10647, n10617, n9450,
    n16347, n14846, n16884, n9622, n16863, n16859, n9939, n10882, n10298,
    n10293, n10740, n10738, n10725, n10775, n10758, n10779, n10772, n10077,
    n10069, n12217, n10834, n10809, n9988, n9982, n9986, n13509, n10042,
    n9874, n14108, n10454, n10453, n10147, n10148, n10156, n11486, n15535,
    n15311, n14928, n14405, n13152, n11684, n10440, n10416, n9266, n9256,
    n10387, n9237, n9211, n9193, n9860, n9056, n12990, n16462, n15328,
    n9640, n9601, n10598, n14622, n10518, n16669, n15333, n15329, n10590,
    n16676, n9353, n10681, n15352, n10586, n10550, n10169, n10197, n10174,
    n10229, n9370, n9363, n9440, n13430, n9145, n9155, n9130, n11580,
    n11552, n11567, n11626, n11636, n11562, n12005, n12021, n12099, n13793,
    n14602, n15267, n16357, n15239, n15341, n15218, n14808, n14507, n14381,
    n14300, n13746, n13356, n13367, n14659, n14644, n14514, n14388, n10559,
    n10526, n10523, n10513, n10190, n12939, n12830, n9497, n9480, n16476,
    n9522, n10909, n12873, n14726, n15885, n15160, n10812, n10797, n14125,
    n10786, n10783, n10765, n10762, n10427, n10040, n10041, n9852, n9807,
    n9754, n13834, n13842, n14760, n15517, n10419, n13617, n10267, n13213,
    n13241, n9923, n15649, n14550, n14190, n14260, n13937, n13753, n13756,
    n12636, n12694, n12696, n9691, n9222, n9228, n9995, n10020, n9563,
    n10344, n10705, n10503, n13026, n13349, n13977, n13469, n9659, n9654,
    n15354, n15360, n16605, n13410, n14035, n14032, n14718, n14579, n14596,
    n14594, n14713, n14715, n15252, n15183, n14654, n14509, n13743, n13395,
    n13336, n13335, n13234, n14352, n9737, n14439, n10936, n13525, n13523,
    n13819, n10469, n15136, n15127, n14307, n14252, n14268, n13984, n13217,
    n13215, n13156, n10637, n16504, n16502, n16558, n16556, n16568, n16571,
    n16589, n16587, n15782, n16619, n16616, n16459, n16460, n16457, n16640,
    n16648, n16647, n15833, n15855, n16668, n16662, n15867, n16711, n16709,
    n16700, n15893, n15904, n15900, n16737, n15921, n15923, n15946, n16757,
    n16763, n15991, n15679, n16190, n16189, n16116, n16111, n16110, n16796,
    n16891, n16889, n16887, n16020, n16019, n16013, n16014, n16058, n16252,
    n16817, n16821, n14637, n16303, n16300, n16129, n16126, n16125, n16135,
    n16109, n16164, n16168, n16256, n16073, n9205, n9583, n9605, n16825,
    n16824, n16925, n13257, n14014, n16630, n16924, n16913, n14992, n16731,
    n16666, n16660, n9635, n16584, n9937, n9933, n9932, n9798, n16307,
    n16154, n14924, n16113, n10732, n13690, n16260, n16248, n16249, n10330,
    n10329, n10325, n9253, n9234, n9209, n9568, n9029, n9060, n13013,
    n9488, n9508, n10623, n9647, n12671, n10680, n10194, n10196, n10177,
    n10173, n9360, n9156, n11419, n9167, n11629, n11854, n11863, n12009,
    n12107, n12515, n13038, n13255, n13775, n13032, n14012, n14584, n14695,
    n14578, n15189, n15198, n15265, n15181, n15565, n10498, n10207, n12392,
    n12391, n11760, n9382, n16412, n15574, n15445, n14994, n15003, n14855,
    n14640, n14506, n14491, n16886, n14365, n14277, n14078, n13954, n16878,
    n13722, n9476, n9388, n11527, n9327, n9326, n8994, n8993, n8989, n9515,
    n12839, n9915, n10903, n10436, n9965, n9966, n10464, n10459, n11480,
    n11485, n11481, n11280, n11305, n10149, n13484, n13491, n14899, n15298,
    n14944, n10848, n10845, n14413, n14556, n10371, n10392, n11308, n9896,
    n12596, n12348, n15309, n14825, n14207, n13810, n13693, n13580, n13570,
    n13196, n13082, n13088, n13141, n9999, n16175, n12740, n15057, n9814,
    n11653, n11660, n10107, n14147, n13997, n10897, n10690, n10610, n10592,
    n10575, n10415, n9272, n11615, n9218, n9629, n9214, n9215, n9587,
    n9198, n9586, n9021, n9548, n12550, n12199, n14321, n15595, n15583,
    n15582, n14624, n15142, n15141, n9352, n10165, n15603, n13714, n13466,
    n13468, n10214, n9365, n14162, n14164, n10538, n10536, n9392, n9395,
    n15604, n9657, n16948, n10698, n10490, n10673, n10633, n10652, n10618,
    n10603, n10568, n10532, n9486, n9464, n9144, n9095, n11416, n11858,
    n11874, n11319, n12529, n13030, n13269, n13056, n13767, n14027, n14576,
    n14710, n15179, n14704, n15282, n15374, n15389, n15367, n15385, n15376,
    n15460, n16659, n14101, n14071, n12662, n9438, n9439, n9417, n9413,
    n11525, n16387, n16348, n15467, n15017, n14863, n14849, n14794, n16723,
    n14299, n13976, n13745, n13866, n13650, n13332, n9621, n13129, n13132,
    n11887, n9391, n9346, n8988, n9338, n15184, n15192, n14698, n14015,
    n10205, n9614, n11628, n9157, n15509, n10881, n15510, n10841, n10859,
    n10860, n15738, n12434, n14056, n9898, n12086, n9990, n10146, n14724,
    n10744, n10278, n10025, n15829, n13512, n9803, n11744, n11745, n10727,
    n10144, n12439, n16318, n16224, n16331, n10894, n10805, n10819, n10752,
    n10457, n10155, n11241, n11300, n11597, n11504, n12561, n11197, n15126,
    n10716, n15104, n15430, n15042, n15070, n15091, n15952, n14398, n15936,
    n13938, n14116, n13607, n15826, n12953, n11841, n15684, n15318, n14954,
    n14832, n14880, n14239, n13987, n13986, n13940, n13939, n13192, n13193,
    n13170, n13153, n12955, n12904, n12892, n12038, n11675, n10961, n11674,
    n10984, n15585, n10691, n8958, n10114, n9720, n10636, n9710, n10641,
    n16236, n9010, n12785, n12181, n14755, n11962, n14457, n11804, n13840,
    n10390, n11714, n13487, n12571, n11519, n12158, n10058, n11262, n11163,
    n11114, n11282, n9945, n11054, n9185, n9540, n11251, n10991, n9071,
    n9176, n11044, n9460, n11009, n12825, n15355, n13596, n15215, n15222,
    n13419, n9644, n13418, n12301, n14324, n14322, n14331, n15611, n9604,
    n12429, n9427, n14652, n14625, n14623, n15143, n15150, n13901, n14044,
    n14042, n15337, n15335, n15347, n9507, n9506, n12981, n12972, n14476,
    n14483, n14805, n14810, n14165, n14163, n14173, n16550, n15596, n9651,
    n10256, n10257, n10585, n10551, n10170, n16645, n10233, n10231, n9374,
    n13325, n9581, n9535, n12402, n9441, n13429, n12110, n9125, n9123,
    n12537, n13054, n13277, n13791, n14600, n15208, n15378, n15273, n15285,
    n15255, n15395, n15372, n15380, n16359, n15626, n13744, n15290, n13382,
    n13381, n13370, n13115, n12938, n12782, n12649, n11531, n9738, n8999,
    n10541, n15206, n9634, n12518, n12012, n11585, n11570, n11418, n11002,
    n11356, n10980, n10133, n12847, n15527, n15524, n10303, n15090, n13292,
    n14438, n14445, n14444, n12877, n12875, n14735, n14734, n10124, n14133,
    n14131, n14058, n14057, n15165, n10009, n10008, n9784, n14609, n14608,
    n14618, n14617, n13520, n14919, n14911, n10142, n15427, n10137, n10136,
    n10134, n14111, n10808, n10822, n10789, n10768, n10475, n10428, n10429,
    n10311, n10291, n13076, n9885, n9858, n9806, n15690, n9760, n11507,
    n13497, n14766, n15027, n14981, n15501, n14873, n14670, n14524, n14335,
    n14201, n13071, n13069, n11918, n16382, n13757, n13627, n13624, n12604,
    n12388, n12272, n12359, n10349, n14155, n14005, n9751, n13880, n13459,
    n9736, n13308, n13452, n16328, n13124, n16324, n12315, n14754, n12564,
    n11600, n10055, n11609, n10022, n11299, n9566, n9567, n11492, n9919,
    n11039, n11473, n10996, n11007, n10953, n9672, n10710, n9660, n15363,
    n13163, n13796, n14039, n14604, n14603, n14721, n15211, n14573, n14432,
    n14655, n14510, n14384, n13752, n13393, n13450, n13340, n13239, n13447,
    n13337, n13236, n12654, n10942, n10486, n15139, n15138, n14253, n14269,
    n13824, n13933, n13227, n13162, n13208, n13251, n13180, n13211, n13248,
    n13177, n12913, n13169, n12887, n9332, n16021, n13226, n8934, n16401,
    n15707, n16554, n16564, n16575, n16623, n16657, n16699, n16048, n13646,
    n9471, n11582, n9386, n9940, n9559, n9542, n9093, n15554, n10558,
    n9612, n12587, n10236, n14636, n16594, n15229, n14638, n9987, n10126,
    n15696, n9195, n10687, n10650, n10530, n14787, n16405, n16730, n13870,
    n9821, n10462, n10863, n14926, n11668, n9225, n9944, n9457, n9003,
    n12793, n16410, n14428, n15625, n8972, n14129, n15835, n10141, n16130,
    n14402, n14235, n11249, n12484, n9477, n9004, n9600, n11852, n13741,
    n11989, n14000, n15776, n10353, n13461, n12733, n13490, n11359, n11658,
    n12882, n8936, n8935, n8940, n8938, n8937, n8939, n8944, n8941, n9811,
    n9833, n8942, n9859, n8946, n8945, n8947, n8948, n9005, n8952, n13165,
    n9013, n8955, n8957, n8956, n8966, n8969, n8967, n9017, n13460, n8971,
    n10121, n8976, n8977, n8982, n8978, n8980, n9589, n9080, n9077, n8991,
    n8992, n8998, n9085, n9000, n9007, n9009, n11667, n9744, n9016, n11686,
    n9018, n9022, n10345, n9032, n9418, n9034, n9033, n9036, n9035, n9040,
    n9048, n9039, n9763, n9042, n9041, n9045, n9047, n9050, n9049, n9051,
    n9436, n9434, n9055, n9437, n9456, n9057, n9063, n9059, n9064, n9061,
    n9062, n9066, n9177, n9076, n9893, n9072, n9074, n13309, n9073, n9075,
    n16961, n9081, n9082, n9345, n9083, n9086, n9090, n11327, n9091, n9092,
    n9097, n9105, n9099, n9100, n9103, n9102, n9104, n9111, n11991, n9106,
    n11349, n9108, n11348, n9109, n9110, n9129, n9113, n9112, n9116,
    n11342, n9115, n9114, n11316, n11341, n9119, n9117, n9118, n9121,
    n9120, n9154, n9122, n9127, n9124, n15396, n9126, n9128, n9140, n9143,
    n12465, n9141, n9142, n9153, n9151, n9152, n9175, n9160, n9158, n9159,
    n9163, n9161, n9162, n9164, n9166, n9165, n11425, n9168, n9170, n9169,
    n9171, n9173, n9172, n9174, n9180, n9541, n9190, n9565, n9611, n10052,
    n9227, n10217, n9236, n9238, n9241, n10215, n9243, n10241, n9247,
    n9250, n9252, n10189, n9255, n9257, n9260, n10187, n9262, n9265, n9267,
    n9270, n10362, n9275, n9276, n9277, n10439, n9281, n9282, n9693, n9292,
    n9288, n9290, n9289, n9291, n13037, n9294, n9293, n9295, n9320, n9297,
    n9296, n9301, n9299, n9298, n9300, n9317, n9303, n9302, n9307, n9305,
    n9304, n9306, n9315, n9309, n9308, n9313, n9311, n9310, n9312, n9314,
    n9316, n9318, n9319, n9321, n9330, n11888, n9333, n9337, n10521,
    n10540, n9339, n9340, n16798, n11539, n9348, n14355, n9359, n9349,
    n13999, n9358, n13434, n9351, n9350, n9357, n10631, n9377, n9369,
    n9375, n9373, n9372, n9376, n9378, n9402, n9381, n11767, n9403, n9650,
    n11885, n9390, n9400, n12653, n12316, n9396, n9397, n9401, n9661,
    n16947, n9404, n9407, n9406, n11026, n9409, n9410, n9412, n9415, n9414,
    n9416, n9420, n9419, n11540, n9422, n9421, n9426, n9424, n9423, n16471,
    n16470, n16472, n12430, n9429, n11971, n9433, n9432, n9435, n9455,
    n9453, n11001, n12255, n9445, n9443, n9442, n9444, n12421, n11969,
    n9448, n9447, n16495, n11970, n12201, n9449, n9452, n9451, n9462,
    n9454, n9458, n9461, n9465, n9469, n9467, n9466, n9468, n16506, n9470,
    n9473, n16517, n9472, n12458, n9475, n11049, n9479, n16523, n9482,
    n9481, n9487, n9483, n12659, n9484, n16522, n9490, n9489, n12186,
    n9498, n9496, n9495, n9500, n9499, n9528, n9503, n12790, n9505, n9504,
    n12467, n9510, n12673, n9513, n9514, n9525, n9524, n9526, n9529,
    n12684, n9531, n9530, n9533, n9532, n9534, n9539, n9537, n12761, n9538,
    n12548, n9546, n9545, n9547, n9558, n9550, n9549, n9557, n9577, n9553,
    n9555, n9554, n9556, n9560, n9562, n9574, n9572, n9571, n9573, n13016,
    n9576, n9575, n9582, n9578, n9580, n9579, n9585, n9584, n12966, n9595,
    n9588, n9593, n9613, n9592, n9594, n13315, n9597, n9596, n9599, n9602,
    n9606, n9607, n13406, n9615, n13052, n13041, n13230, n9627, n10201,
    n9637, n9636, n16610, n9643, n9642, n9648, n9652, n9655, n9658, n9690,
    n13182, n13006, n12687, n12416, n12078, n11902, n11706, n11548, n11389,
    n9679, n9677, n9675, n9673, n10967, n9671, n9669, n9667, n10951, n9665,
    n10943, n10946, n10945, n9663, n10949, n10948, n9664, n10950, n9666,
    n10952, n9668, n10954, n9670, n11024, n11076, n11171, n11390, n11549,
    n11707, n11903, n12079, n12417, n12688, n13007, n13183, n9688, n9689,
    n9695, n9698, n9701, n9703, n9704, n9708, n9713, n9714, n9716, n9718,
    n9723, n9725, n9730, n10321, n10323, n9740, n14356, n9739, n9741,
    n9746, n9745, n9781, n9753, n9758, n9757, n9759, n11719, n9762, n11843,
    n15534, n11840, n9769, n9765, n9764, n11922, n9767, n9766, n9768,
    n11377, n9775, n9774, n10901, n9772, n9771, n9773, n11378, n9778,
    n9776, n9777, n9794, n9780, n9779, n9785, n9783, n9782, n15683, n9792,
    n9788, n9786, n11198, n9787, n9790, n11014, n9789, n9793, n9797,
    n11723, n9796, n15701, n9795, n9802, n9800, n9799, n11747, n9805,
    n9804, n9809, n9808, n12496, n9817, n9815, n9834, n11407, n9812,
    n12480, n9816, n9818, n9822, n9820, n9819, n9823, n9825, n9824, n12509,
    n9827, n9826, n9828, n9830, n9829, n9831, n15715, n9843, n10842, n9835,
    n9836, n11226, n9839, n9837, n9838, n9840, n15714, n9842, n9844, n9848,
    n9846, n9845, n9849, n9847, n12506, n9851, n9850, n12507, n12085,
    n9853, n9854, n12084, n9856, n9855, n9857, n15722, n9868, n9866, n9861,
    n11203, n9864, n9862, n9863, n9865, n15723, n9867, n9869, n9873, n9871,
    n9870, n9875, n12324, n9879, n9877, n9876, n9878, n12349, n9888, n9881,
    n9880, n9886, n12707, n9884, n9883, n15739, n9887, n9891, n9890, n9892,
    n9912, n9897, n9895, n9894, n12371, n9906, n12449, n9900, n9899, n9904,
    n9902, n9901, n9903, n9905, n9907, n9909, n9908, n9910, n9918, n9917,
    n9922, n11019, n9921, n15750, n12850, n9927, n9926, n9931, n9929,
    n9928, n9930, n9936, n9935, n9941, n9963, n9942, n11055, n9947, n9946,
    n9948, n12879, n9952, n9951, n9956, n9954, n9953, n9955, n9958, n12870,
    n9962, n9961, n9967, n12871, n12857, n9974, n9972, n9970, n9971,
    n15788, n9983, n12920, n9977, n9976, n9981, n9979, n9978, n9980, n9985,
    n9994, n15802, n13298, n10004, n10003, n10007, n10006, n10010, n13288,
    n10014, n10013, n10019, n10018, n13289, n10023, n11497, n10027, n10026,
    n13517, n10031, n10030, n10034, n10033, n10036, n13501, n10037, n10039,
    n10038, n10051, n10262, n10054, n11435, n10060, n10059, n15819, n10070,
    n13060, n10064, n10063, n10068, n10066, n10065, n10067, n10073, n10072,
    n10078, n10080, n10079, n10081, n10106, n10083, n10082, n10087, n10085,
    n10084, n10086, n10103, n10089, n10088, n10093, n10091, n10090, n10092,
    n10101, n10095, n10094, n10099, n10097, n10096, n10098, n10100, n10102,
    n10104, n10105, n10113, n10108, n10109, n10117, n13221, n10122, n16369,
    n10129, n10125, n10140, n10127, n16332, n11911, n10128, n10130, n10132,
    n10968, n10138, n11654, n10162, n10143, n10145, n11603, n10160, n13881,
    n15515, n10153, n10152, n10154, n10159, n10161, n10163, n14583, n10184,
    n10168, n10167, n13973, n10182, n10176, n10175, n13869, n10178, n10181,
    n10183, n10186, n10185, n10260, n10510, n16637, n10507, n10195, n10203,
    n13635, n10221, n10220, n16461, n10227, n13653, n10230, n10234, n10232,
    n10235, n10238, n13594, n10242, n10250, n10244, n10243, n10246, n10245,
    n10248, n14587, n10249, n16628, n10255, n10506, n10264, n13524, n10368,
    n10266, n15839, n10271, n10365, n10281, n10284, n10283, n15849, n13536,
    n10288, n10287, n10292, n10290, n10289, n10360, n10359, n10302, n10300,
    n10318, n10316, n10304, n10305, n12565, n10314, n10306, n14112, n10308,
    n10307, n10312, n10310, n10309, n10313, n10315, n10317, n10319, n10326,
    n10328, n10331, n10333, n10335, n10334, n10338, n10340, n10339, n10343,
    n10347, n10346, n10348, n10351, n10352, n10355, n10354, n10356, n10361,
    n14109, n10366, n10367, n10369, n10370, n13797, n14134, n10377, n10376,
    n10381, n10379, n10378, n10380, n10382, n10385, n10389, n10391, n13619,
    n10395, n10398, n10413, n14055, n10443, n10418, n15888, n10424, n10423,
    n10426, n10430, n10438, n10465, n10463, n10442, n10444, n10446, n10449,
    n10447, n10448, n15880, n10456, n10455, n10728, n10468, n10466, n10485,
    n10483, n10477, n10472, n10471, n10473, n10474, n10481, n10479, n14762,
    n10480, n10482, n10563, n10581, n10491, n10493, n10492, n10494, n10504,
    n10497, n10496, n10502, n10697, n13400, n10500, n10499, n15589, n10509,
    n10516, n10511, n10512, n14075, n10519, n14043, n10522, n16658, n10529,
    n10528, n10531, n10539, n10543, n10542, n16679, n10548, n10547, n14296,
    n16680, n10557, n14323, n16695, n10570, n10565, n10564, n10566, n10567,
    n14492, n10574, n14475, n12490, n10578, n10588, n10583, n10582, n10584,
    n10591, n10594, n10597, n10605, n10600, n10599, n10601, n10602, n16724,
    n10609, n10612, n10616, n10615, n10621, n10619, n10626, n10625, n15330,
    n10635, n10629, n10628, n10630, n10632, n15343, n10643, n10654, n10649,
    n10648, n10651, n10665, n10666, n10675, n10669, n10668, n10670, n10672,
    n10683, n15353, n10685, n10689, n10694, n16778, n10696, n10695, n10701,
    n10699, n10702, n10708, n10704, n10703, n10709, n10886, n10713, n10712,
    n15322, n10715, n10717, n10720, n13674, n14437, n10731, n15902, n10735,
    n12491, n10754, n10749, n10748, n10750, n10751, n10753, n10755, n10760,
    n14400, n10763, n10766, n10769, n10780, n12883, n10784, n10787, n10790,
    n14908, n10794, n10793, n10799, n10798, n14907, n10803, n10802, n13125,
    n10817, n10816, n10820, n15949, n10823, n10829, n15038, n10846, n15983,
    n15039, n15425, n10868, n10867, n10873, n10870, n10884, n10885, n10891,
    n10890, n10892, n10893, n10895, n15673, n10900, n13882, n10919, n10916,
    n10918, n10924, n10923, n10928, n10925, n10927, n10929, n10938, n10934,
    n10931, n10944, n10947, n10957, n10956, n10960, n10959, n10965, n10964,
    n10979, n10971, n10970, n10972, n13673, n11185, n10975, n10973, n10974,
    n11381, n10976, n10977, n10978, n10983, n10981, n15122, n10982, n10985,
    n10988, n10986, n10987, n10990, n10989, n10993, n10992, n10995, n10994,
    n10998, n10997, n11000, n10999, n11004, n11003, n11006, n11005, n11013,
    n11008, n11011, n11010, n11012, n11018, n11016, n11455, n11015, n11017,
    n11023, n11021, n11020, n11022, n11028, n11027, n11030, n11029, n11032,
    n11031, n11034, n11033, n11036, n11035, n11038, n11037, n11041, n11040,
    n11043, n11042, n11046, n11201, n11045, n11048, n11047, n11051, n11050,
    n11053, n11052, n11059, n11057, n11056, n11058, n12312, n11061, n11060,
    n11063, n11062, n11065, n11064, n11067, n11066, n11069, n11068, n11071,
    n11073, n11072, n11075, n11074, n11083, n11079, n11078, n11081, n11080,
    n11082, n11085, n11084, n11087, n11086, n11089, n11088, n11091, n11090,
    n11093, n11092, n11095, n11094, n11097, n11096, n11099, n11098, n11107,
    n11103, n11102, n11105, n11104, n11106, n11109, n11108, n11111, n11110,
    n11113, n11112, n11116, n11115, n11118, n11117, n11120, n11119, n11122,
    n11121, n11124, n11123, n11126, n11125, n11128, n11127, n11130, n11129,
    n11132, n11131, n11134, n11133, n11136, n11135, n11138, n11137, n11140,
    n11139, n11142, n11141, n11144, n11143, n11146, n11145, n11148, n11147,
    n11150, n11149, n11152, n11151, n11154, n11153, n11156, n11155, n11158,
    n11157, n11160, n11159, n11162, n11161, n11166, n11164, n11165, n11168,
    n11167, n11170, n11169, n11174, n11173, n11176, n11175, n11178, n11177,
    n11180, n11179, n11182, n11181, n11184, n11183, n12853, n11193, n11447,
    n11446, n11448, n11186, n11394, n11393, n11395, n11187, n11222, n11221,
    n11223, n11188, n11371, n11370, n11372, n11189, n11466, n11465, n11467,
    n11190, n11240, n11239, n11191, n11484, n11207, n11192, n11276, n11194,
    n11195, n11216, n11196, n15119, n11214, n16330, n15137, n11210, n11273,
    n11442, n11441, n11443, n11199, n11399, n11398, n11400, n11200, n11228,
    n11227, n11229, n11202, n11363, n11362, n11364, n11204, n11461, n11460,
    n11462, n11205, n11245, n11244, n11246, n11206, n11479, n11208, n11291,
    n11212, n11213, n11215, n11218, n11217, n11220, n11219, n11225, n11224,
    n11236, n11233, n11231, n11230, n11232, n11234, n12499, n11235, n11238,
    n11237, n11243, n11242, n11255, n11248, n11247, n11250, n12448, n11253,
    n11252, n11254, n11257, n11256, n11259, n11258, n11261, n11260, n11264,
    n11263, n11266, n11265, n11271, n11269, n11268, n11270, n11274, n11601,
    n11286, n11279, n11278, n11281, n12868, n11284, n11283, n11285, n11288,
    n11287, n11290, n11289, n11295, n11294, n11298, n11297, n11313, n11303,
    n11307, n11306, n11309, n13284, n11311, n11310, n11312, n11315, n11314,
    n11317, n11320, n11318, n11334, n11321, n11330, n11325, n11323, n11324,
    n11326, n11328, n11329, n11332, n11331, n11333, n11336, n11335, n11338,
    n11337, n11340, n11339, n11355, n11343, n11347, n11345, n11346, n11353,
    n11350, n11351, n11352, n11354, n11358, n11357, n11361, n11360, n11368,
    n11366, n11365, n11367, n11369, n12090, n11376, n11374, n11373, n11375,
    n11388, n11646, n11379, n11387, n11380, n11384, n11383, n11385, n11386,
    n11412, n11392, n11397, n11396, n11411, n11402, n11401, n11406, n11404,
    n11403, n11405, n11409, n11408, n11410, n11413, n11415, n11414, n12205,
    n11417, n11424, n11422, n11420, n11421, n11423, n11431, n11427, n11429,
    n11430, n11432, n11434, n11433, n11436, n11438, n11437, n11440, n11439,
    n11445, n11444, n11452, n11450, n11449, n11451, n11454, n11453, n11457,
    n11456, n11459, n11458, n11464, n11463, n11471, n11469, n11468, n11470,
    n11472, n12329, n11476, n11474, n11475, n11478, n11477, n11483, n11482,
    n11490, n11488, n11487, n11489, n11491, n12845, n11494, n11493, n11496,
    n11495, n11500, n11498, n13504, n11499, n11514, n11502, n11506, n11505,
    n11512, n11509, n11510, n11511, n11513, n11516, n11515, n11518, n11517,
    n11521, n12149, n11520, n11523, n11522, n11985, n11545, n11774, n11536,
    n16854, n11538, n11543, n15559, n11999, n11541, n11542, n11896, n11544,
    n11547, n11546, n11551, n11555, n11559, n11558, n11561, n11565, n11564,
    n11566, n11593, n11576, n11579, n12680, n11577, n11578, n11591, n11589,
    n11590, n11592, n11595, n11861, n11594, n11608, n11599, n12150, n11602,
    n11604, n11606, n11605, n11607, n11614, n11611, n12159, n11612, n11613,
    n11620, n11617, n11616, n11619, n11618, n11622, n11621, n11624, n11623,
    n11625, n12191, n11627, n11635, n11633, n11631, n11632, n11634, n11639,
    n11637, n11638, n11640, n11642, n11641, n11645, n11739, n11652, n11650,
    n11648, n11647, n11649, n11651, n11656, n11657, n11673, n15691, n11931,
    n16238, n16158, n15816, n15103, n14669, n11665, n11664, n15637, n11666,
    n11671, n15533, n11913, n11669, n11670, n11676, n11672, n11678, n11677,
    n11702, n15703, n11925, n16237, n11930, n16242, n11680, n15680, n16245,
    n11815, n11681, n11690, n11928, n11682, n11685, n15687, n12478, n11688,
    n11687, n11689, n12479, n11699, n11691, n12041, n11694, n11692, n11693,
    n12472, n11697, n12482, n11695, n11696, n11698, n11700, n11703, n11701,
    n11705, n11704, n11709, n11711, n11710, n11713, n11712, n11716, n11715,
    n11718, n11717, n11721, n11720, n11730, n11728, n11725, n11726, n11727,
    n11729, n11732, n11731, n11734, n11733, n11736, n11735, n11738, n11737,
    n11743, n11741, n11740, n11742, n11750, n11746, n11748, n11749, n11771,
    n16479, n16489, n11772, n16853, n11753, n11752, n11758, n16411, n11756,
    n11755, n11757, n11765, n12724, n11762, n11764, n12729, n11766, n11769,
    n16431, n11768, n11899, n11770, n11799, n11776, n11775, n11778, n11777,
    n12135, n16850, n11790, n12131, n11780, n11779, n11781, n11785, n11783,
    n11782, n11784, n11794, n11788, n11787, n11789, n12136, n11792, n11791,
    n12251, n11793, n12253, n11795, n11797, n11796, n11893, n11798, n11801,
    n11800, n11803, n11802, n11806, n13828, n11805, n11808, n11807, n11828,
    n11842, n11810, n11809, n11826, n16063, n16160, n16159, n11813, n12043,
    n11844, n11824, n11816, n16064, n11817, n11821, n11819, n11818, n11820,
    n11823, n11822, n11846, n11825, n11829, n11827, n11831, n11830, n11839,
    n15660, n11837, n11836, n11838, n11851, n15074, n11849, n12477, n11845,
    n11847, n11848, n11850, n12545, n11857, n11871, n11869, n11862, n11866,
    n11865, n11867, n11868, n11870, n11879, n11877, n11878, n11880, n11882,
    n11881, n11895, n11894, n11898, n11897, n11901, n11900, n11905, n11907,
    n11906, n11909, n11908, n11917, n11912, n11914, n11915, n11916, n11921,
    n11919, n11920, n11940, n11948, n11924, n11923, n11938, n11927, n11926,
    n16161, n11950, n11936, n11929, n11935, n11933, n11932, n11934, n11952,
    n11937, n11941, n11939, n11943, n11942, n11945, n11944, n11947, n11946,
    n11957, n11955, n12952, n11951, n11953, n11954, n11956, n11959, n11958,
    n11961, n11960, n11964, n14449, n11963, n11966, n11965, n11968, n11967,
    n11977, n11972, n11973, n11975, n11974, n11976, n11979, n14167, n11978,
    n11981, n11980, n11983, n11992, n11996, n12307, n11994, n11993, n11995,
    n12003, n11998, n12000, n12001, n12002, n12008, n12031, n12013, n12017,
    n12016, n12018, n12027, n13021, n12024, n12025, n12026, n12029, n12028,
    n12030, n12033, n12032, n12063, n12037, n12035, n12034, n12036, n12059,
    n12039, n12042, n12040, n12062, n12057, n12343, n16067, n12366, n12215,
    n12044, n12236, n12066, n12049, n12047, n12046, n12048, n12053, n16244,
    n12051, n12052, n12067, n13560, n12054, n12055, n12056, n12058, n12061,
    n12060, n12072, n12065, n12064, n12070, n12068, n12069, n12073, n12071,
    n12075, n12074, n12077, n12076, n12081, n12083, n12082, n12097, n12087,
    n12095, n12089, n12088, n12093, n12091, n12092, n12094, n12096, n12102,
    n12120, n12103, n12963, n12105, n12104, n12106, n12118, n12111, n12112,
    n12115, n12114, n12116, n12117, n12119, n12128, n12126, n12127, n12145,
    n12129, n12287, n16849, n12285, n12130, n12275, n12132, n12134, n12133,
    n12140, n12286, n12300, n12138, n12137, n12139, n12303, n12142, n12141,
    n12143, n12146, n12144, n12148, n12147, n12171, n12154, n12153, n12157,
    n12156, n12168, n12163, n12162, n12166, n12165, n12167, n12169, n13526,
    n12170, n12173, n12172, n12175, n12174, n12178, n12177, n12180, n12179,
    n12183, n12182, n12185, n12184, n12188, n12196, n12190, n12189, n12194,
    n12192, n12193, n12195, n12198, n12197, n12200, n12202, n12210, n12204,
    n12203, n12208, n12206, n12207, n12209, n12212, n12211, n12214, n12213,
    n12216, n12338, n15730, n12341, n12337, n16254, n12218, n12447, n12362,
    n12242, n12219, n12223, n12221, n12220, n12222, n12269, n12234, n12224,
    n12226, n12225, n12263, n12230, n12228, n12227, n12229, n12232, n12231,
    n12233, n12244, n12237, n12342, n15742, n12239, n12241, n12240, n12363,
    n12262, n12918, n12243, n12250, n12248, n12246, n12245, n12247, n12249,
    n12609, n12252, n12254, n12259, n12257, n12256, n12258, n12261, n12260,
    n12271, n12267, n12265, n12264, n12266, n12268, n12270, n12274, n12273,
    n12295, n12277, n16510, n12276, n12278, n16855, n12394, n12279, n12280,
    n12284, n12282, n12281, n12283, n12290, n12288, n12401, n12663, n12289,
    n12668, n12291, n12293, n12292, n12296, n12294, n12298, n12297, n12299,
    n12305, n12302, n12304, n12306, n12309, n12308, n12311, n12310, n12314,
    n12313, n12318, n12317, n12320, n12319, n12336, n12321, n12437, n12323,
    n12325, n12326, n12334, n12328, n12327, n12332, n12330, n12331, n12333,
    n12335, n12358, n12340, n12339, n12347, n12706, n12345, n12344, n12346,
    n12716, n12355, n12717, n12353, n12351, n12350, n12352, n12354, n12356,
    n12357, n12361, n12360, n12387, n15759, n16077, n12580, n12379, n12368,
    n12369, n16166, n12585, n12588, n12374, n12377, n12376, n12378, n12384,
    n12697, n12382, n12380, n12693, n12381, n12383, n12385, n12386, n12390,
    n12389, n12412, n12393, n12617, n12395, n12399, n12397, n12396, n12398,
    n12406, n12616, n12404, n12403, n12607, n12794, n12405, n12799, n12408,
    n12410, n12409, n12413, n12411, n12415, n12414, n12419, n12423, n12422,
    n12428, n12426, n12425, n12427, n12433, n12431, n12432, n12436, n12438,
    n12443, n12441, n12442, n12444, n12457, n12446, n12445, n12455, n12453,
    n12451, n12450, n12452, n12454, n12456, n12460, n12464, n12462, n12461,
    n12463, n12466, n12469, n12468, n12471, n12470, n12476, n12474, n12473,
    n12475, n12489, n15653, n12487, n12481, n12483, n12485, n12486, n12488,
    n12495, n12493, n12492, n12494, n12498, n12497, n12505, n12503, n12501,
    n13502, n12500, n12502, n12504, n12512, n12508, n12510, n12511, n12514,
    n12513, n12526, n12519, n12520, n12523, n12522, n12524, n12525, n12527,
    n13415, n12534, n12532, n12533, n12542, n12540, n12541, n12544, n12543,
    n12555, n12546, n12553, n12549, n12551, n12552, n12554, n12557, n12556,
    n12559, n12563, n12562, n12570, n12566, n12568, n12567, n12569, n12577,
    n13482, n13481, n12574, n12573, n12575, n12576, n12603, n12893, n12578,
    n12579, n12581, n12634, n12584, n12583, n12601, n12739, n12586, n12591,
    n12589, n12590, n12595, n12593, n12592, n12594, n12597, n12598, n12633,
    n12599, n12600, n12602, n12606, n12605, n12608, n12774, n12642, n16423,
    n12613, n12611, n12610, n12612, n12628, n12625, n12615, n12614, n12624,
    n12619, n12618, n12764, n12620, n12622, n12621, n12623, n12646, n12626,
    n12627, n12630, n12629, n12632, n12631, n12641, n12639, n12635, n12637,
    n12638, n12640, n12648, n12644, n12643, n12645, n12647, n12651, n12650,
    n12656, n12655, n12658, n12657, n12661, n12660, n12667, n12665, n12664,
    n12666, n12670, n12669, n12672, n12674, n12679, n12677, n12676, n12678,
    n12681, n12683, n12682, n12686, n12685, n12690, n12692, n12691, n12703,
    n12695, n12701, n12699, n12698, n12700, n12702, n12705, n12704, n12715,
    n12709, n12708, n12711, n12710, n12713, n12712, n12714, n12721, n12719,
    n12718, n12720, n12723, n12722, n12728, n12726, n12725, n12727, n12731,
    n12730, n12732, n12737, n16218, n12735, n12734, n12736, n12757, n12738,
    n12896, n12741, n12743, n12742, n12745, n12890, n12919, n12754, n12907,
    n12906, n12748, n12930, n12752, n12750, n12749, n12751, n12753, n12755,
    n12756, n12760, n12759, n12781, n16861, n12763, n12767, n12766, n12812,
    n12768, n12773, n12771, n12770, n12772, n12777, n12775, n12804, n12824,
    n12776, n12826, n12779, n12778, n12780, n12784, n12783, n12787, n12786,
    n12789, n12788, n12792, n12791, n12798, n12796, n12795, n12797, n12801,
    n12800, n12803, n12802, n12809, n12807, n12805, n12984, n12806, n12808,
    n12823, n12811, n12813, n12993, n12815, n12819, n12817, n12816, n12818,
    n12821, n12820, n12822, n12833, n12828, n12827, n12829, n12831, n12832,
    n12835, n12834, n12838, n12840, n12844, n12842, n12841, n12843, n12846,
    n12849, n12848, n12852, n12851, n12854, n12856, n12855, n12865, n12859,
    n12863, n12861, n12860, n12862, n12864, n12867, n12866, n12878, n12869,
    n12876, n12874, n12881, n12880, n12885, n12884, n12886, n12914, n16177,
    n13063, n12905, n12894, n16083, n12895, n12898, n16075, n12897, n12899,
    n12902, n12901, n12903, n12908, n12951, n12910, n12909, n12911, n12917,
    n12916, n12928, n12922, n12921, n12926, n15083, n12924, n12923, n12925,
    n12927, n12934, n12932, n12931, n12933, n12936, n12935, n12943, n12991,
    n12937, n12941, n12940, n12942, n12946, n12945, n12948, n12947, n12950,
    n12949, n12960, n12958, n12954, n12956, n12957, n12959, n12962, n12961,
    n12973, n12964, n12971, n12967, n12969, n12970, n12975, n12974, n12977,
    n12980, n12979, n12983, n12982, n12989, n12987, n12985, n13102, n12986,
    n12988, n13005, n12992, n12995, n12996, n13001, n12999, n12998, n13000,
    n13003, n13002, n13004, n13009, n13012, n13014, n13020, n13018, n13017,
    n13019, n13022, n13025, n13024, n13028, n13027, n13033, n13051, n13035,
    n13034, n13036, n13049, n13042, n13043, n13046, n13045, n13047, n13048,
    n13050, n13059, n13057, n13058, n13072, n13070, n16181, n13062, n13140,
    n13068, n13187, n13098, n13075, n13074, n13149, n13077, n13079, n13195,
    n13083, n13081, n13080, n13085, n13084, n13086, n13095, n13090, n13091,
    n13246, n13093, n13092, n13094, n13096, n13097, n13100, n13099, n13107,
    n13105, n13330, n13104, n13106, n13118, n13108, n13318, n13109, n13110,
    n13114, n13112, n13111, n13113, n13116, n13117, n16962, n13121, n13126,
    n13136, n13130, n13134, n13133, n13135, n13139, n13138, n13146, n13142,
    n13144, n13172, n13145, n13155, n13148, n13147, n13150, n13151, n13160,
    n13158, n13157, n13159, n13161, n13164, n13167, n13166, n13168, n13178,
    n13171, n13173, n13181, n13185, n13209, n13188, n13191, n13194, n13549,
    n13198, n13197, n13199, n13201, n13203, n13220, n13204, n13205, n13212,
    n13218, n13216, n13229, n13225, n13223, n13222, n13224, n13228, n13237,
    n13231, n13240, n13249, n13242, n13252, n13254, n13253, n13266, n13259,
    n13260, n13263, n13262, n13777, n13264, n13265, n13267, n13342, n13274,
    n13766, n13272, n13273, n13282, n13790, n13280, n13281, n13285, n13287,
    n13286, n13297, n13291, n13294, n13299, n13304, n13306, n13311, n13310,
    n13312, n13338, n13317, n13316, n13321, n13319, n13323, n13377, n13324,
    n13329, n13327, n13326, n13328, n13361, n13331, n13334, n13339, n13341,
    n13345, n13343, n13344, n13355, n13347, n13351, n13350, n13352, n13358,
    n13357, n13371, n13359, n13363, n13365, n13636, n13366, n13369, n13368,
    n13385, n13373, n13372, n13374, n13379, n13647, n13384, n13386, n13388,
    n13394, n13392, n13391, n13396, n13405, n13399, n13398, n13403, n13436,
    n13401, n13404, n13408, n13414, n13412, n13411, n13413, n13416, n13417,
    n13421, n13420, n13428, n13423, n13422, n13426, n13424, n16801, n13427,
    n13440, n13433, n13432, n13438, n13435, n16933, n13439, n13448, n13443,
    n13451, n13455, n13457, n13463, n13462, n13464, n13467, n13475, n13471,
    n13774, n13473, n13472, n13474, n13476, n13478, n13498, n13486, n13485,
    n13495, n13489, n13493, n13492, n13494, n13496, n14114, n13500, n13499,
    n13516, n13505, n13507, n13506, n13514, n13510, n13518, n13535, n13531,
    n13527, n13529, n13528, n13530, n13532, n13538, n13537, n13540, n13539,
    n13566, n13543, n13542, n13564, n16185, n13567, n13551, n13569, n13555,
    n13554, n13556, n13608, n16187, n13687, n13691, n13572, n13576, n13577,
    n13578, n13590, n13582, n13586, n13584, n13583, n13585, n13587, n13593,
    n13591, n14024, n13592, n13602, n13598, n13597, n13599, n13613, n13606,
    n13605, n13616, n13630, n13623, n13621, n13620, n13622, n13633, n13638,
    n16874, n13729, n13640, n13639, n13659, n13642, n13641, n13643, n13649,
    n13716, n13655, n13662, n13654, n13656, n13660, n13668, n13665, n13671,
    n13676, n13675, n13677, n13681, n13684, n13689, n13799, n13806, n13696,
    n13695, n13697, n13701, n13702, n13705, n13709, n13707, n13706, n13708,
    n13710, n13864, n13721, n13951, n13724, n13723, n13725, n13856, n16456,
    n13855, n13959, n16386, n13732, n13735, n13738, n13742, n13748, n13747,
    n13749, n13755, n13761, n13764, n14026, n13770, n13788, n13772, n13771,
    n13773, n13786, n13778, n13780, n13783, n13782, n13784, n13785, n13787,
    n14033, n13794, n13795, n16229, n16230, n14185, n13911, n14180, n13807,
    n13913, n13916, n14186, n13812, n13811, n13813, n13815, n13818, n14212,
    n13823, n13821, n13820, n13822, n13831, n13829, n14137, n13830, n13850,
    n13836, n13838, n13837, n13848, n13844, n13846, n13845, n13847, n13849,
    n13852, n15586, n13851, n13853, n13858, n13857, n13861, n13860, n13862,
    n13873, n13872, n13874, n13878, n13884, n13883, n13885, n13893, n13890,
    n13896, n13899, n13908, n13904, n13902, n14707, n13903, n13906, n13905,
    n13907, n13909, n13918, n13917, n13919, n13923, n13924, n13928, n13932,
    n13930, n13929, n13931, n13945, n13948, n16650, n16651, n13953, n14070,
    n13956, n13955, n13957, n13961, n14084, n13964, n13967, n13970, n13975,
    n13974, n13979, n13978, n13980, n13992, n13995, n14002, n14001, n14003,
    n14007, n14895, n14006, n14008, n14011, n14010, n14023, n14016, n14017,
    n14020, n14019, n14586, n14021, n14022, n14025, n14575, n14030, n14031,
    n14599, n14038, n14046, n14045, n14052, n14050, n14048, n15188, n14049,
    n14051, n14053, n14067, n14065, n14061, n14466, n14063, n14062, n14064,
    n14066, n14068, n14073, n14077, n14274, n14081, n14080, n14082, n14085,
    n14283, n14086, n14091, n14094, n14099, n14097, n14098, n14103, n14102,
    n14104, n14127, n14126, n14122, n14120, n14115, n14118, n14117, n14119,
    n14121, n14123, n14144, n14142, n14138, n14140, n14139, n14141, n14143,
    n14145, n14151, n14423, n14150, n14152, n14159, n14891, n14158, n14160,
    n14166, n14174, n14170, n14168, n15274, n14169, n14172, n14171, n14228,
    n16192, n14183, n14188, n14206, n14189, n14236, n14191, n14193, n14214,
    n14243, n14199, n14197, n14196, n14198, n14200, n14208, n14216, n14215,
    n14217, n14222, n14225, n16106, n16196, n14234, n14399, n14403, n14240,
    n14245, n14247, n14250, n14249, n14251, n14258, n14264, n14263, n14266,
    n14265, n14267, n14276, n14362, n14279, n14278, n14280, n14290, n14293,
    n14297, n14302, n14301, n14303, n14308, n14316, n14319, n14326, n14325,
    n14332, n14330, n14328, n15399, n14327, n14329, n14339, n14338, n14346,
    n14349, n14353, n14354, n14358, n14568, n14357, n14359, n14364, n14488,
    n14367, n14366, n14368, n14370, n14380, n14494, n14383, n14382, n14393,
    n14396, n16198, n14548, n14407, n14406, n14408, n14410, n14416, n14415,
    n14417, n14424, n16906, n16926, n14427, n14430, n14431, n14446, n14442,
    n14440, n15120, n14441, n14443, n14469, n14454, n14452, n14456, n14455,
    n14465, n14461, n14459, n14463, n14462, n14464, n14470, n14478, n14477,
    n14484, n14482, n14480, n14479, n14481, n16888, n14490, n14497, n14648,
    n14499, n14498, n14500, n14504, n14508, n14519, n14522, n14532, n14535,
    n14538, n14541, n14818, n14549, n14822, n14551, n14553, n14563, n14559,
    n14558, n14560, n14569, n16912, n14571, n14709, n14581, n14580, n14582,
    n14595, n14588, n14589, n14592, n14591, n14697, n14593, n14716, n14619,
    n14615, n14613, n14612, n14614, n14616, n14633, n14629, n14627, n14626,
    n14628, n14630, n14639, n14772, n14643, n14642, n14646, n14651, n14653,
    n14664, n14667, n14673, n14672, n14682, n14680, n14683, n14690, n14688,
    n14691, n14694, n14693, n14706, n14699, n14700, n14703, n14702, n15191,
    n15178, n15207, n14745, n14741, n14739, n14738, n14740, n14742, n14751,
    n14749, n14753, n14752, n14759, n14757, n14761, n14764, n14768, n14774,
    n14776, n16892, n14845, n14777, n14798, n14783, n14853, n14788, n14795,
    n14799, n14802, n14807, n14806, n14814, n14812, n14813, n16117, n16202,
    n14820, n14930, n14898, n14841, n14839, n14842, n14990, n14848, n14847,
    n14867, n14851, n14856, n14858, n14857, n14870, n14868, n14871, n14876,
    n14875, n14889, n14882, n14893, n14896, n16011, n15072, n15071, n15656,
    n16038, n14901, n15640, n14976, n14902, n14903, n14910, n14913, n14912,
    n14916, n14915, n14917, n14920, n16204, n15055, n14933, n15059, n14937,
    n14936, n14938, n14961, n14942, n14947, n14946, n14956, n14964, n14962,
    n14965, n14972, n14969, n16037, n14975, n14977, n14987, n14985, n14988,
    n14993, n16753, n16901, n14996, n15002, n15000, n14999, n15006, n15247,
    n15021, n15009, n15012, n15011, n15024, n15022, n15025, n15034, n15032,
    n15035, n15040, n15041, n15049, n15044, n15043, n15047, n15046, n15048,
    n15050, n16299, n15056, n15307, n15062, n15314, n15064, n15111, n15076,
    n15075, n15084, n15157, n15156, n15098, n15093, n15092, n15096, n15095,
    n15097, n15099, n15113, n15116, n15114, n15117, n15121, n15131, n15129,
    n15124, n15133, n15145, n15144, n15152, n15442, n15147, n15173, n15169,
    n15168, n15171, n15170, n15172, n15174, n15280, n15186, n15185, n15187,
    n15203, n15193, n15194, n15197, n15196, n15257, n15200, n15210, n15217,
    n15216, n15224, n15220, n15231, n15453, n16910, n15232, n15444, n15233,
    n15236, n15243, n15245, n15250, n15248, n15451, n15261, n15259, n15258,
    n15262, n15263, n15264, n15266, n15270, n15275, n15276, n15295, n15293,
    n15296, n15305, n15303, n15313, n16212, n15487, n15316, n15478, n15417,
    n15331, n15340, n15339, n15349, n15345, n15357, n15356, n15359, n15358,
    n15362, n15379, n15387, n15391, n15390, n15392, n15397, n15402, n15400,
    n15401, n15403, n15421, n15419, n15422, n15434, n15432, n15431, n15433,
    n15435, n15440, n16894, n15551, n15448, n15454, n15471, n15458, n15462,
    n15461, n15474, n15472, n15475, n16128, n15481, n15635, n15490, n15645,
    n15544, n15493, n15503, n15505, n15512, n15531, n15529, n15523, n15522,
    n15543, n15547, n15545, n15548, n15553, n15555, n16340, n15624, n15566,
    n15567, n15569, n15570, n15581, n16782, n16353, n15620, n15587, n16808,
    n16397, n15592, n15597, n15610, n15608, n15606, n15605, n15607, n15609,
    n15631, n15629, n15632, n15636, n16370, n15638, n15644, n15642, n15641,
    n15650, n15647, n16366, n15652, n15651, n15668, n15666, n15664, n15665,
    n15672, n15671, n15676, n15675, n15677, n15678, n16001, n15682, n15681,
    n15689, n15686, n15685, n15702, n15688, n15706, n15692, n15693, n15699,
    n15695, n15694, n15717, n15697, n15698, n15700, n15713, n15704, n15705,
    n15710, n15708, n15709, n15711, n15712, n15719, n15716, n15718, n15729,
    n15721, n15720, n15728, n15727, n15725, n15724, n15726, n15737, n15735,
    n15733, n15732, n15734, n15736, n15745, n15741, n15740, n15743, n15744,
    n15749, n15747, n15746, n15748, n15768, n15753, n15752, n15769, n15757,
    n15766, n15755, n15756, n15765, n15758, n15763, n15760, n15761, n15762,
    n15764, n15783, n15767, n15771, n15770, n15775, n15774, n15785, n15779,
    n15778, n15784, n15780, n15787, n15786, n15794, n15791, n15790, n15795,
    n15793, n15799, n15797, n15798, n15809, n15801, n15800, n15808, n15807,
    n15805, n15804, n15806, n15815, n15813, n15811, n15810, n15812, n15814,
    n15825, n15818, n15817, n15824, n15822, n15821, n15823, n15848, n15846,
    n15827, n15828, n15834, n15831, n15832, n15844, n15838, n15837, n15842,
    n15841, n15854, n15843, n15845, n15847, n15859, n15852, n15851, n15862,
    n15857, n15856, n15858, n15868, n15861, n15860, n15866, n15864, n15865,
    n15870, n15869, n15871, n15877, n15872, n15875, n15874, n15876, n15879,
    n15878, n15894, n15881, n15884, n15892, n15886, n15890, n15889, n15891,
    n15906, n15897, n15899, n15903, n15914, n15907, n15909, n15911, n15922,
    n15918, n15917, n15920, n15926, n15924, n15931, n15929, n15928, n15941,
    n15934, n15939, n15938, n15947, n15945, n15957, n15950, n15955, n15954,
    n15963, n15961, n15960, n15967, n15966, n15974, n15971, n15970, n15979,
    n15977, n15976, n15992, n15981, n15980, n15990, n15993, n15995, n16004,
    n16000, n16003, n16005, n16016, n16010, n16009, n16012, n16030, n16024,
    n16022, n16138, n16023, n16031, n16035, n16025, n16032, n16042, n16317,
    n16208, n16043, n16148, n16046, n16145, n16052, n16053, n16057, n16096,
    n16281, n16279, n16066, n16068, n16069, n16070, n16071, n16072, n16074,
    n16080, n16084, n16079, n16264, n16082, n16081, n16087, n16086, n16265,
    n16090, n16268, n16089, n16091, n16092, n16093, n16094, n16095, n16097,
    n16098, n16100, n16102, n16103, n16104, n16105, n16123, n16108, n16114,
    n16118, n16119, n16127, n16147, n16223, n16151, n16153, n16157, n16163,
    n16162, n16165, n16167, n16169, n16171, n16172, n16174, n16176, n16178,
    n16180, n16182, n16184, n16186, n16188, n16191, n16193, n16195, n16197,
    n16199, n16203, n16216, n16217, n16225, n16327, n16305, n16231, n16234,
    n16233, n16288, n16241, n16239, n16240, n16243, n16247, n16246, n16251,
    n16250, n16253, n16255, n16258, n16257, n16262, n16261, n16263, n16267,
    n16266, n16269, n16273, n16272, n16275, n16277, n16278, n16280, n16284,
    n16283, n16285, n16287, n16290, n16292, n16293, n16295, n16298, n16302,
    n16329, n16338, n16336, n16334, n16335, n16337, n16341, n16399, n16344,
    n16350, n16391, n16351, n16355, n16406, n16374, n16375, n16380, n16379,
    n16385, n16384, n16394, n16392, n16395, n16402, n16802, n16903, n16418,
    n16422, n16414, n16413, n16417, n16420, n16435, n16436, n16443, n16440,
    n16445, n16448, n16447, n16450, n16449, n16452, n16451, n16455, n16464,
    n16463, n16469, n16468, n16483, n16474, n16473, n16481, n16478, n16477,
    n16488, n16480, n16484, n16491, n16490, n16493, n16492, n16500, n16498,
    n16497, n16499, n16591, n16509, n16508, n16515, n16511, n16530, n16519,
    n16518, n16528, n16521, n16520, n16534, n16526, n16525, n16524, n16527,
    n16529, n16532, n16531, n16537, n16535, n16536, n16538, n16547, n16541,
    n16545, n16543, n16544, n16546, n16559, n16549, n16552, n16563, n16557,
    n16555, n16569, n16561, n16562, n16567, n16565, n16566, n16581, n16572,
    n16579, n16577, n16578, n16580, n16590, n16583, n16588, n16585, n16596,
    n16593, n16595, n16599, n16598, n16600, n16601, n16602, n16606, n16612,
    n16609, n16611, n16613, n16618, n16635, n16629, n16632, n16641, n16639,
    n16643, n16638, n16649, n16644, n16646, n16655, n16653, n16652, n16684,
    n16656, n16683, n16670, n16664, n16663, n16674, n16667, n16672, n16671,
    n16673, n16688, n16678, n16677, n16690, n16682, n16681, n16685, n16692,
    n16691, n16701, n16694, n16693, n16698, n16697, n16713, n16705, n16704,
    n16710, n16717, n16716, n16719, n16729, n16722, n16725, n16739, n16733,
    n16732, n16736, n16742, n16750, n16751, n16758, n16756, n16755, n16765,
    n16764, n16762, n16761, n16772, n16770, n16768, n16767, n16771, n16789,
    n16777, n16776, n16781, n16780, n16787, n16785, n16784, n16793, n16807,
    n16794, n16805, n16799, n16816, n16803, n16815, n16811, n16810, n16823,
    n16827, n16840, n16838, n16839, n16844, n16846, n16852, n16858, n16856,
    n16857, n16860, n16862, n16864, n16865, n16867, n16869, n16871, n16873,
    n16876, n16877, n16879, n16881, n16883, n16885, n16893, n16942, n16919,
    n16955, n16932, n16950, n16938, n16937, n16945, n16941, n16953, n16951,
    n16954, n16959, n16965, n16963, n16964, n16966, n16969, n16968;
  assign n10912 = ~n10885 & ~n15426;
  assign n16383 = ~n11675 | ~n11674;
  assign n16378 = ~n11675 | ~n11661;
  assign n15414 = n16212 ^ ~n15487;
  assign n15532 = n16214 ^ n15645;
  assign n16419 = ~n11992 | ~n11990;
  assign P1_U3086 = ~P1_STATE_REG_SCAN_IN;
  assign n16358 = ~n9656 & ~n10958;
  assign n15323 = ~n11841 & ~n15654;
  assign n15670 = ~n10900 & ~n10899;
  assign n10299 = ~n10280 | ~n13522;
  assign n13348 = ~n10203 & ~n10202;
  assign n16702 = ~n10580 & ~n10579;
  assign n9283 = ~n10439 | ~n10440;
  assign n15388 = n9087 ^ P2_IR_REG_27__SCAN_IN;
  assign n9325 = ~n9023 | ~n9738;
  assign n9001 = ~n9000 & ~n10520;
  assign n11910 = ~n16236 & ~n16149;
  assign n9343 = ~n9339 & ~n10520;
  assign n10218 = ~n14426 | ~n8919;
  assign n16149 = n9014 ^ n9013;
  assign n8932 = ~n8931;
  assign n8931 = ~n9474;
  assign n14970 = ~n10969 | ~n8919;
  assign n9347 = ~n14355 | ~P2_IR_REG_31__SCAN_IN;
  assign n9087 = ~n9086 | ~P2_IR_REG_31__SCAN_IN;
  assign n9053 = ~n9048 & ~n9047;
  assign n8919 = ~n9043;
  assign n9493 = ~n9107 | ~n8974;
  assign n9043 = ~n9037;
  assign n13718 = ~n13716 | ~n13715;
  assign n10624 = ~n10622;
  assign n13314 = ~n12995 | ~n12994;
  assign n10280 = ~n13524 | ~n13521;
  assign n15674 = ~n15670;
  assign n9770 = n10121 | n10126;
  assign n8950 = n8949 | n8948;
  assign n8933 = ~n8931;
  assign n16453 = ~n10645 & ~n10644;
  assign n9012 = ~n9005 | ~n9006;
  assign n10297 = ~n10299;
  assign n10904 = ~n11843 | ~n9776;
  assign n10906 = ~n9770 & ~n11840;
  assign n11382 = ~P1_IR_REG_0__SCAN_IN;
  assign n15429 = ~n10866 | ~n10865;
  assign n10806 = ~n8920 | ~n15167;
  assign n14900 = n9018 ^ ~P1_IR_REG_27__SCAN_IN;
  assign n15602 = ~n9400 | ~n9399;
  assign n15338 = ~n10654 | ~n10653;
  assign n16936 = ~n16912;
  assign n15240 = ~n16419;
  assign n16442 = ~n16444;
  assign n16438 = ~n16439;
  assign n10958 = ~n9391 | ~P2_STATE_REG_SCAN_IN;
  assign n15516 = ~n11643 | ~n10137;
  assign n15999 = ~n10718 | ~n10717;
  assign n13672 = ~n13680;
  assign n9024 = ~n11891 | ~n9325;
  assign n10963 = ~n10961 | ~n11658;
  assign P2_U3151 = ~P2_STATE_REG_SCAN_IN;
  assign P1_U3973 = ~n10980 & ~P1_U3086;
  assign n8924 = ~n16322;
  assign n8928 = ~n8927;
  assign n10714 = n14156 | n9755;
  assign n9810 = ~n10730 & ~n8919;
  assign n10969 = ~n10730;
  assign n9430 = ~n12429 | ~n12430;
  assign n16045 = ~n16332 | ~n16322;
  assign n14804 = n10622 ^ n10623;
  assign n8918 = n9087 ^ P2_IR_REG_27__SCAN_IN;
  assign n14149 = ~n9359;
  assign n9957 = ~n10121 & ~n11843;
  assign n16446 = ~n16443 | ~n16442;
  assign n16441 = ~n16443 | ~n16438;
  assign n16430 = ~n16421 | ~n16420;
  assign n16222 = ~n16221 | ~n16220;
  assign n16421 = ~n16437 | ~n16419;
  assign n16352 = ~n16391 | ~n16419;
  assign n16221 = ~n16153 | ~n16236;
  assign n16220 = ~n16219 | ~n16218;
  assign n15571 = ~n15624 & ~n15569;
  assign n16219 = n16217 ^ ~n8924;
  assign n15628 = ~n15624 & ~n15623;
  assign n16326 = ~n16325 | ~n16324;
  assign n16144 = ~n16143 | ~n8924;
  assign n16921 = ~n16920 | ~n8922;
  assign n16944 = ~n16943 & ~n8925;
  assign n16920 = ~n16942 | ~n16919;
  assign n16943 = ~n16942 & ~n16941;
  assign n16429 = ~n16428 & ~n16427;
  assign n16343 = ~n16399;
  assign n15466 = ~n15459 | ~n15458;
  assign n16143 = ~n16142 | ~n16317;
  assign n15294 = ~n15295 | ~n16438;
  assign n16142 = ~n16141 | ~n16140;
  assign n16150 = ~n16148;
  assign n16041 = ~n16040 | ~n16208;
  assign n16342 = ~n16341 & ~n16900;
  assign n15297 = ~n15295 | ~n16442;
  assign n15558 = ~n15556 | ~n16340;
  assign n16428 = ~n16432 & ~n16423;
  assign n15507 = ~n15506 & ~n15505;
  assign n15326 = ~n15325 | ~n15324;
  assign n15459 = ~n15471 | ~n16419;
  assign n15622 = ~n15616 & ~n15615;
  assign n15491 = ~n15532 & ~n11663;
  assign n14689 = ~n14690 | ~n16438;
  assign n16432 = ~n16422;
  assign n16040 = ~n16036 | ~n16035;
  assign n16949 = ~n16948 & ~n16947;
  assign n14692 = ~n14690 | ~n16442;
  assign n15506 = ~n15532 & ~n15653;
  assign n16140 = ~n16320 & ~n16139;
  assign n16321 = ~n16319 & ~n16318;
  assign n15616 = ~n15620 & ~n15594;
  assign n15325 = ~n15417 | ~n13226;
  assign n16916 = ~n16911 | ~n16910;
  assign n16211 = ~n16210 & ~n16209;
  assign n15556 = ~n15554 | ~n16898;
  assign n15621 = ~n15620 | ~n15619;
  assign n16141 = ~n16137 | ~n16136;
  assign n15327 = ~n15313 & ~n15312;
  assign n15023 = ~n15024 | ~n16438;
  assign n16843 = ~n16842 | ~n16841;
  assign n16837 = ~n16842 & ~n16836;
  assign n16319 = ~n16316 & ~n16315;
  assign n16911 = ~n16909 & ~n16908;
  assign n16036 = ~n16317 | ~n16034;
  assign n15082 = ~n15069 & ~n15068;
  assign n16209 = ~n16208 | ~n16207;
  assign n16363 = ~n16362 & ~n16361;
  assign n15246 = ~n15289 & ~n15244;
  assign n15026 = ~n15024 | ~n16442;
  assign n16029 = ~n16028 | ~n16027;
  assign n16931 = ~n16930 & ~n16929;
  assign n16320 = ~n16208;
  assign n15016 = ~n15010 | ~n15009;
  assign n14539 = ~n14540 | ~n16442;
  assign n16316 = ~n16312 & ~n16311;
  assign n15053 = ~n15041 | ~n15511;
  assign n16930 = ~n16915 | ~n16914;
  assign n16909 = ~n16907 | ~n16934;
  assign n16832 = ~n16831 | ~n16830;
  assign n15177 = ~n15165 | ~n15511;
  assign n14574 = ~n16936 | ~n16424;
  assign n14979 = ~n14978 & ~n14977;
  assign n16027 = ~n16031 | ~n16026;
  assign n14542 = ~n14540 | ~n16438;
  assign n15289 = ~n15238 | ~n15237;
  assign n15312 = ~n15414 & ~n15653;
  assign n16362 = ~n16387 & ~n16356;
  assign n15483 = ~n15480 & ~n15479;
  assign n16210 = ~n16317 | ~n16154;
  assign n15365 = ~n15354 | ~n15596;
  assign n16814 = ~n16813 | ~n16812;
  assign n16946 = ~n16936 | ~n16935;
  assign n15069 = ~n15111 & ~n15323;
  assign n16136 = ~n16311 & ~n16135;
  assign n10941 = ~n10940 | ~n10939;
  assign n15415 = ~n15414 & ~n16365;
  assign n15450 = ~n15445 | ~n15557;
  assign n14963 = ~n14964 | ~n16381;
  assign n14953 = ~n14943 | ~n14942;
  assign n16915 = ~n16912 | ~n16933;
  assign n16907 = ~n16904 & ~n16903;
  assign n15081 = ~n15080 | ~n15079;
  assign n15102 = ~n15090 | ~n15511;
  assign n16908 = ~n16912 & ~n16933;
  assign n16312 = ~n16310 & ~n16309;
  assign n16835 = ~n16912 | ~n16591;
  assign n16311 = ~n16132 | ~n16131;
  assign n16836 = ~n16912 & ~n16925;
  assign n16039 = ~n16037;
  assign n15319 = ~n15317 | ~n15478;
  assign n16026 = ~n16035 | ~n16032;
  assign n10940 = ~n10922 | ~n10921;
  assign n15615 = ~n15614 | ~n15613;
  assign n15029 = ~n16037 & ~n15536;
  assign n14966 = ~n14964 | ~n16377;
  assign n15663 = ~n15662 | ~n15661;
  assign n15480 = ~n15482 & ~n15481;
  assign n14978 = ~n16037 & ~n15497;
  assign n14540 = ~n14537 | ~n14686;
  assign n15351 = ~n15337 | ~n15596;
  assign n14433 = ~n16926 | ~n16424;
  assign n14943 = ~n14961 | ~n13226;
  assign n16309 = ~n16308;
  assign n16904 = ~n16902 | ~n16901;
  assign n16372 = ~n16368 | ~n16367;
  assign n16315 = ~n16314 & ~n16313;
  assign n16131 = ~n16314 | ~n16313;
  assign n15662 = ~n16368 | ~n15659;
  assign n16137 = ~n16129 | ~n16308;
  assign n14905 = ~n14904 & ~n14903;
  assign n15614 = ~n15600 | ~n15599;
  assign n10922 = ~n10917;
  assign n15109 = ~n15104 | ~n15103;
  assign n15317 = ~n15315 & ~n15479;
  assign n15154 = ~n15143 | ~n15596;
  assign n10939 = ~n10938 & ~n10937;
  assign n14360 = ~n14352 | ~n14351;
  assign n16820 = ~n16816;
  assign n16826 = ~n16825 | ~n16824;
  assign n16829 = ~n16822 | ~n16821;
  assign n15066 = n15065 & n15064;
  assign n16804 = ~n16816 | ~n16803;
  assign n15067 = ~n15104 | ~n15057;
  assign n16028 = ~n16020 | ~n16019;
  assign n14537 = ~n16926 | ~n14685;
  assign n16015 = ~n16014 | ~n16013;
  assign n16139 = ~n16314 & ~n16138;
  assign n10937 = ~n10936 | ~n10935;
  assign n15315 = ~n16212 & ~n15316;
  assign n14923 = ~n14911 | ~n15511;
  assign n15619 = ~n15618 & ~n15617;
  assign n16434 = ~n16818 & ~n16433;
  assign n15416 = ~n15413 | ~n15412;
  assign n15304 = ~n15303 | ~n15302;
  assign n14570 = ~n14968 & ~n10218;
  assign n14904 = ~n16134 & ~n15497;
  assign n15226 = ~n15215 | ~n15596;
  assign n15158 = ~n15156 & ~n15155;
  assign n10357 = ~n14968 & ~n13123;
  assign n14840 = ~n14841 | ~n16377;
  assign n14869 = ~n14870 | ~n16442;
  assign n14800 = ~n14801 | ~n16438;
  assign n16427 = ~n16426 | ~n16425;
  assign n14803 = ~n14801 | ~n16442;
  assign n14982 = ~n16134 & ~n15536;
  assign n16934 = ~n16906 | ~n16905;
  assign n16902 = ~n16900 & ~n16899;
  assign n14887 = ~n14879 & ~n14878;
  assign n14952 = ~n14951 & ~n14950;
  assign n16314 = ~n16134;
  assign n14872 = ~n14870 | ~n16438;
  assign n15482 = ~n16214;
  assign n14843 = ~n14841 | ~n16381;
  assign n15065 = ~n15063 | ~n15314;
  assign n15465 = ~n15464 & ~n15463;
  assign n14793 = ~n14784 | ~n14783;
  assign n15594 = ~n15618 | ~n15593;
  assign n14862 = ~n14852 | ~n14851;
  assign n15412 = ~n15411 & ~n15410;
  assign n15541 = ~n15540 | ~n15539;
  assign n16818 = ~n16802;
  assign n16310 = ~n16307 & ~n16306;
  assign n16006 = ~n16008 & ~n16007;
  assign n14959 = ~n14954 & ~n16365;
  assign n15332 = ~n15328 & ~n15338;
  assign n15618 = n16900 ^ ~n15591;
  assign n16800 = ~n16802 & ~n16591;
  assign n16017 = ~n16010 | ~n16009;
  assign n15469 = ~n15467 & ~n16431;
  assign n15063 = ~n15060 & ~n15479;
  assign n14998 = ~n14996 | ~n15557;
  assign n14161 = ~n14155 | ~n14154;
  assign n14153 = ~n14155 | ~n14351;
  assign n16215 = n16018 ^ ~n16370;
  assign n15504 = ~n15501 | ~n15500;
  assign n15658 = ~n14973;
  assign n14968 = n10350 ^ ~n10349;
  assign n14801 = ~n14798 | ~n14797;
  assign n10935 = ~n10934 & ~n10933;
  assign n15302 = ~n15301 & ~n15300;
  assign n14941 = ~n14954 & ~n11663;
  assign n10350 = ~n10343 | ~n10342;
  assign n15301 = ~n15409 & ~n15074;
  assign n14973 = ~n16011 | ~n15656;
  assign n15079 = ~n15078 & ~n15077;
  assign n15500 = ~n15499 & ~n15498;
  assign n15060 = ~n15062 & ~n15061;
  assign n14886 = ~n14885 | ~n14884;
  assign n16361 = ~n16360 | ~n16359;
  assign n10920 = ~n10914 | ~n10913;
  assign n15108 = ~n15107 & ~n15106;
  assign n10910 = ~n10909 | ~n10908;
  assign n10933 = ~n10932 | ~n10931;
  assign n10905 = ~n10903 | ~n10902;
  assign n14877 = ~n14829 | ~n14828;
  assign n16792 = ~n16791 & ~n16790;
  assign n14425 = ~n14890 & ~n10218;
  assign n15411 = ~n15409 & ~n15534;
  assign n15539 = ~n15538 & ~n15537;
  assign n16398 = ~n16397;
  assign n16007 = ~n15676 & ~n15675;
  assign n10883 = ~n10882 | ~n10881;
  assign n16408 = ~n16407 & ~n16809;
  assign n16306 = ~n16305 & ~n16304;
  assign n16806 = ~n16795 | ~n16794;
  assign n15078 = ~n15105 & ~n15074;
  assign n16403 = ~n16400 | ~n8921;
  assign n10707 = ~n10706 & ~n10705;
  assign n14684 = ~n14682 | ~n16377;
  assign n15593 = n15592 & n15596;
  assign n14890 = n14148 ^ ~n14147;
  assign n16008 = ~n15672 | ~n15671;
  assign n14837 = ~n14880 | ~n15103;
  assign n16896 = ~n16894 | ~n16893;
  assign n16791 = ~n16777 | ~n16776;
  assign n14829 = ~n14880 | ~n15057;
  assign n14997 = ~n14993 | ~n14992;
  assign n14816 = ~n14805 | ~n15596;
  assign n15613 = ~n15612 & ~n15611;
  assign n15599 = ~n15598 & ~n15597;
  assign n15499 = ~n15535 & ~n15074;
  assign n15364 = ~n15363 & ~n15362;
  assign n15107 = ~n15105 & ~n15534;
  assign n15530 = ~n15529 & ~n15528;
  assign n15538 = ~n15535 & ~n15534;
  assign n15477 = ~n16049;
  assign n10902 = ~n15674 | ~n10901;
  assign n10908 = ~n15674 | ~n10907;
  assign n15409 = ~n15299 | ~n15496;
  assign n15061 = ~n16206;
  assign n14747 = ~n14734 | ~n15511;
  assign n14681 = ~n14682 | ~n16381;
  assign n15015 = ~n15014 & ~n15013;
  assign n14668 = ~n14666 | ~n16438;
  assign n14658 = ~n14647 | ~n14646;
  assign n15568 = ~n16773 & ~n15564;
  assign n10688 = ~n10687 & ~n15572;
  assign n16206 = ~n15975 | ~n16301;
  assign n10913 = ~n10725 | ~n10724;
  assign n16304 = ~n16303 & ~n16302;
  assign n15528 = ~n15527 | ~n15526;
  assign n15578 = ~n16898;
  assign n15623 = ~n16773 & ~n16433;
  assign n16407 = ~n16808;
  assign n16124 = ~n16123 & ~n16297;
  assign n16339 = ~n16773 | ~n16775;
  assign n16790 = ~n16781 & ~n16780;
  assign n14665 = ~n14666 | ~n16442;
  assign n10706 = ~n16773 & ~n15601;
  assign n14148 = ~n10338 | ~n10337;
  assign n15646 = ~n15669 | ~n15670;
  assign n14939 = ~n14934 | ~n15059;
  assign n16400 = ~n14894;
  assign n14934 = ~n14932 & ~n15479;
  assign n15019 = ~n15017 & ~n16431;
  assign n10721 = ~n15997 | ~n10901;
  assign n15552 = ~n15573 | ~n15575;
  assign n15975 = ~n16299;
  assign n15526 = ~n15525 & ~n15524;
  assign n15468 = ~n15573 & ~n16433;
  assign n14733 = ~n14728 & ~n14727;
  assign n14894 = n13998 ^ ~n13997;
  assign n15361 = ~n15573 & ~n15601;
  assign n15310 = ~n15309 & ~n15308;
  assign n15007 = ~n15017 & ~n15455;
  assign n10724 = ~n15997 | ~n10907;
  assign n15077 = ~n15076 | ~n15075;
  assign n14778 = ~n14845 | ~n14777;
  assign n14533 = ~n14534 | ~n16377;
  assign n15463 = ~n15462 | ~n15461;
  assign n14536 = ~n14534 | ~n16381;
  assign n14679 = ~n14670 | ~n14669;
  assign n16898 = n16778 ^ ~n16779;
  assign n14566 = ~n14565 & ~n14564;
  assign n15437 = ~n15436 | ~n15435;
  assign n13886 = ~n13880 | ~n14154;
  assign n13854 = ~n13880 | ~n14351;
  assign n16773 = ~n16778;
  assign n15153 = ~n15152 & ~n15151;
  assign n10861 = ~n10860 & ~n10859;
  assign n14621 = ~n14608 | ~n15511;
  assign n16783 = ~n15576 | ~n15575;
  assign n14728 = ~n14726 & ~n14725;
  assign n15588 = ~n15585 & ~n10218;
  assign n15573 = ~n15576;
  assign n14635 = ~n14625 | ~n15596;
  assign n14523 = ~n14521 | ~n16438;
  assign n14513 = ~n14505 | ~n14504;
  assign n14958 = ~n14957 | ~n14956;
  assign n14950 = ~n14949 | ~n14948;
  assign n15306 = ~n15429 & ~n15520;
  assign n14861 = ~n14860 & ~n14859;
  assign n14828 = ~n14827 & ~n14826;
  assign n14866 = ~n14865 & ~n14864;
  assign n15997 = ~n15519;
  assign n14932 = ~n14933 & ~n16204;
  assign n16301 = ~n15429 | ~n15308;
  assign n16227 = ~n15999 | ~n15519;
  assign n14534 = ~n14531 | ~n14530;
  assign n10622 = ~n10609 | ~n10608;
  assign n14565 = ~n14554 & ~n14553;
  assign n14520 = ~n14521 | ~n16442;
  assign n14860 = ~n14863 & ~n16356;
  assign n14827 = ~n14825 & ~n15479;
  assign n14317 = ~n14318 | ~n16377;
  assign n14531 = ~n14524 | ~n14669;
  assign n15054 = ~n16204;
  assign n15244 = ~n15243 | ~n15242;
  assign n14421 = ~n14420 & ~n14419;
  assign n13678 = ~n13672 | ~n14154;
  assign n14320 = ~n14318 | ~n16381;
  assign n14957 = ~n14955 | ~n16367;
  assign n15151 = ~n15150 | ~n15149;
  assign n14865 = ~n14863 & ~n16386;
  assign n9742 = ~n9737 & ~n13679;
  assign n14645 = ~n14640 & ~n11752;
  assign n15163 = ~n15162 & ~n15161;
  assign n13685 = ~n13682 & ~n13681;
  assign n14949 = ~n14955 | ~n15659;
  assign n15519 = ~n10720 & ~n10719;
  assign n15576 = ~n10685 | ~n10684;
  assign n10840 = ~n10839 & ~n10838;
  assign n14955 = n15072 & n14945;
  assign n14420 = ~n14411 & ~n14410;
  assign n14884 = ~n14883 & ~n14882;
  assign n15162 = ~n15160 & ~n15159;
  assign n10898 = ~n10328 | ~n10327;
  assign n15052 = ~n15051 & ~n15050;
  assign n10682 = ~n16759 & ~n10681;
  assign n14387 = ~n14371 | ~n14370;
  assign n10866 = ~n13459 | ~n9810;
  assign n14797 = ~n14796 & ~n14795;
  assign n15242 = ~n15241 & ~n15240;
  assign n14948 = ~n14947 & ~n14946;
  assign n14836 = ~n14835 & ~n14834;
  assign n14792 = ~n14791 & ~n14790;
  assign n14397 = ~n14395 | ~n16438;
  assign n10831 = ~n15161 & ~n10830;
  assign n14347 = ~n14348 | ~n16381;
  assign n14350 = ~n14348 | ~n16377;
  assign n14255 = ~n14254 & ~n14253;
  assign n10839 = ~n10835 & ~n15160;
  assign n10838 = ~n10837 & ~n15159;
  assign n10487 = ~n10469 & ~n15426;
  assign n14394 = ~n14395 | ~n16442;
  assign n15149 = ~n15148 & ~n15147;
  assign n13682 = ~n13680 & ~n13679;
  assign n14448 = ~n14438 | ~n15511;
  assign n16766 = ~n16448 & ~n16447;
  assign n14530 = ~n14529 & ~n14528;
  assign n15987 = ~n15971 & ~n15970;
  assign n14552 = ~n14550 | ~n15637;
  assign n14315 = ~n14307 | ~n14669;
  assign n14223 = ~n14224 | ~n16377;
  assign n15148 = ~n15442 & ~n15601;
  assign n14254 = ~n14248 & ~n14247;
  assign n14294 = ~n14292 | ~n16438;
  assign n14835 = ~n14881 & ~n15534;
  assign n14272 = ~n14259 | ~n14258;
  assign n14544 = ~n14402 & ~n14401;
  assign n14791 = ~n14794 & ~n16356;
  assign n14226 = ~n14224 | ~n16381;
  assign n15443 = ~n15446 | ~n15442;
  assign n10858 = ~n10856 | ~n10855;
  assign n15982 = ~n15972;
  assign n13680 = n10692 ^ n10691;
  assign n14503 = ~n14491 & ~n11752;
  assign n14306 = ~n14298 | ~n14297;
  assign n15161 = ~n10834 & ~n10833;
  assign n10837 = ~n10836;
  assign n10835 = ~n10836 & ~n10833;
  assign n14291 = ~n14292 | ~n16442;
  assign n14929 = ~n16202;
  assign n15350 = ~n15349 & ~n15348;
  assign n14796 = ~n14794 & ~n16386;
  assign n15051 = ~n15984 & ~n15518;
  assign n10664 = ~n10663 | ~n10662;
  assign n10692 = ~n10323 & ~n10322;
  assign n10662 = ~n15234 | ~n10661;
  assign n16121 = ~n15968 | ~n15983;
  assign n16054 = ~n15968 & ~n15983;
  assign n15176 = ~n15175 & ~n15174;
  assign n10657 = ~n10656 | ~n10655;
  assign n14345 = ~n14335 | ~n14669;
  assign n14662 = ~n14661 & ~n14660;
  assign n14881 = ~n14944 | ~n14831;
  assign n14995 = ~n16754;
  assign n15972 = ~n15968 & ~n15969;
  assign n10836 = ~n10832 & ~n15155;
  assign n14676 = ~n14675 | ~n14674;
  assign n15348 = ~n15347 | ~n15346;
  assign n15962 = ~n15961 & ~n15960;
  assign n13458 = ~n13456 & ~n13455;
  assign n14564 = ~n14563 | ~n14562;
  assign n14314 = ~n14313 & ~n14312;
  assign n10663 = ~n10659 | ~n10658;
  assign n14248 = ~n14313 & ~n14246;
  assign n14657 = ~n14656 & ~n14655;
  assign n14204 = ~n14203 & ~n14202;
  assign n14675 = ~n14671 | ~n16367;
  assign n10811 = ~n10810 | ~n10809;
  assign n15175 = ~n15166 & ~n15518;
  assign n14271 = ~n14270 & ~n14269;
  assign n13456 = ~n13453 & ~n13679;
  assign n9735 = ~n9734 | ~n9733;
  assign n15013 = ~n15012 | ~n15011;
  assign n15956 = ~n15959 & ~n15958;
  assign n14927 = ~n15166 & ~n15045;
  assign n15225 = ~n15224 & ~n15223;
  assign n15346 = n15345 & n15344;
  assign n14409 = ~n14405 | ~n15637;
  assign n14834 = ~n14833 | ~n14832;
  assign n14517 = ~n14516 & ~n14515;
  assign n14661 = ~n14659 & ~n16386;
  assign n15228 = ~n15234 & ~n15227;
  assign n14512 = ~n14511 & ~n14510;
  assign n14221 = ~n14220 & ~n14219;
  assign n14203 = ~n14194 & ~n14193;
  assign n14313 = ~n14241 | ~n14240;
  assign n14369 = ~n14365 & ~n11752;
  assign n14656 = ~n14659 & ~n16356;
  assign n15155 = ~n15088;
  assign n13993 = ~n13994 | ~n16381;
  assign n15166 = ~n15965;
  assign n14502 = ~n14501 | ~n14500;
  assign n13307 = ~n13305 & ~n13304;
  assign n10660 = ~n16454 | ~n15214;
  assign n14211 = ~n14260 & ~n11663;
  assign n15223 = ~n15222 | ~n15221;
  assign n14095 = ~n14093 | ~n16442;
  assign n16745 = ~n16746 & ~n16455;
  assign n16200 = ~n14819 | ~n14817;
  assign n14419 = ~n14418 | ~n14417;
  assign n14671 = n14557 & n14830;
  assign n14107 = ~n14099 | ~n14098;
  assign n14516 = ~n14514 & ~n16431;
  assign n14821 = ~n16050;
  assign n14859 = ~n14858 | ~n14857;
  assign n14286 = ~n14281 | ~n14280;
  assign n14220 = ~n14260 & ~n16365;
  assign n15959 = ~n15951 & ~n15950;
  assign n9734 = ~n9725 | ~n9724;
  assign n10679 = ~n13452 | ~n8921;
  assign n14528 = ~n14527 | ~n14526;
  assign n14344 = ~n14343 & ~n14342;
  assign n14241 = ~n14239 | ~n15637;
  assign n13996 = ~n13994 | ~n16377;
  assign n16895 = ~n14844 | ~n15004;
  assign n14146 = ~n14133 | ~n15511;
  assign n14815 = ~n14814 & ~n14813;
  assign n15227 = ~n15343;
  assign n16746 = ~n16452 | ~n16451;
  assign n14124 = ~n14111 | ~n15511;
  assign n15958 = ~n15955 | ~n15954;
  assign n14732 = ~n14731 | ~n14730;
  assign n16747 = ~n15338 & ~n14991;
  assign n14527 = ~n14525 | ~n16367;
  assign n15214 = ~n15329;
  assign n15965 = ~n10801 | ~n10800;
  assign n14844 = ~n16454 | ~n14991;
  assign n14281 = ~n14277 | ~n15557;
  assign n13949 = ~n13947 | ~n16381;
  assign n15005 = ~n15004;
  assign n14922 = ~n14921 & ~n14920;
  assign n16050 = ~n15948 & ~n15953;
  assign n14823 = ~n16115;
  assign n15101 = ~n15100 & ~n15099;
  assign n13946 = ~n13947 | ~n16377;
  assign n14562 = ~n14561 & ~n14560;
  assign n14343 = ~n14192 | ~n14191;
  assign n14674 = ~n14673 & ~n14672;
  assign n15221 = ~n15220 & ~n15219;
  assign n13305 = ~n13302 & ~n13679;
  assign n13936 = ~n13925 | ~n13924;
  assign n14238 = ~n14403 | ~n14237;
  assign n14391 = ~n14390 & ~n14389;
  assign n14386 = ~n14385 & ~n14384;
  assign n15948 = ~n15952;
  assign n14090 = ~n14089 & ~n14088;
  assign n14096 = ~n14083 & ~n14082;
  assign n13826 = ~n13825 & ~n13824;
  assign n14192 = ~n14190 | ~n15637;
  assign n14106 = ~n14105 & ~n14104;
  assign n13991 = ~n13984 | ~n14669;
  assign n14289 = ~n14288 & ~n14287;
  assign n13968 = ~n13969 | ~n16442;
  assign n13983 = ~n13975 | ~n13974;
  assign n14305 = ~n14304 & ~n14303;
  assign n14811 = ~n14810 | ~n14809;
  assign n10640 = ~n13301 | ~n8921;
  assign n10824 = ~n15952 & ~n9770;
  assign n14921 = ~n14918 | ~n14917;
  assign n14132 = ~n14128 & ~n14127;
  assign n10776 = ~n14730 | ~n14606;
  assign n15943 = ~n15935 & ~n15934;
  assign n14525 = ~n14556 & ~n14414;
  assign n14128 = ~n14126 & ~n14125;
  assign n14775 = ~n16735 | ~n16731;
  assign n14730 = ~n10779 | ~n10778;
  assign n14210 = ~n14209 | ~n14208;
  assign n13935 = ~n13934 & ~n13933;
  assign n13762 = ~n13763 | ~n16381;
  assign n13943 = ~n13942 & ~n13941;
  assign n13122 = ~n13120 & ~n16962;
  assign n14285 = ~n14299 & ~n15455;
  assign n14288 = ~n14299 & ~n16431;
  assign n14725 = ~n14607 | ~n14606;
  assign n14918 = ~n15932 | ~n15428;
  assign n10320 = ~n10303 & ~n15426;
  assign n14746 = ~n14745 & ~n14744;
  assign n14110 = ~n14127 & ~n14126;
  assign n13825 = ~n13816 & ~n13815;
  assign n14089 = ~n14100 & ~n16386;
  assign n14909 = ~n10794 & ~n10793;
  assign n14312 = ~n14311 | ~n14310;
  assign n14543 = ~n15932 & ~n15933;
  assign n16890 = ~n16718;
  assign n14083 = ~n14078 & ~n11752;
  assign n16728 = ~n16727 & ~n16726;
  assign n15287 = n15279 & n15278;
  assign n14105 = ~n14100 & ~n16356;
  assign n14634 = ~n14633 & ~n14632;
  assign n13128 = ~n13127 & ~n13126;
  assign n14390 = ~n14388 & ~n16386;
  assign n13713 = ~n13703 | ~n13702;
  assign n13765 = ~n13763 | ~n16377;
  assign n14385 = ~n14388 & ~n16356;
  assign n13629 = ~n13631 | ~n16381;
  assign n13972 = ~n13963 & ~n13962;
  assign n10815 = ~n13124 & ~n14967;
  assign n13632 = ~n13631 | ~n16377;
  assign n16112 = ~n15936 & ~n15933;
  assign n10645 = ~n13124 & ~n10218;
  assign n14311 = ~n14244 | ~n14412;
  assign n14632 = ~n14631 | ~n14630;
  assign n13922 = ~n13937 & ~n11663;
  assign n14545 = ~n15936 & ~n15937;
  assign n15932 = ~n15936;
  assign n15278 = ~n15277 & ~n15276;
  assign n16735 = ~n16730;
  assign n14555 = ~n15936 | ~n14413;
  assign n13990 = ~n13989 & ~n13988;
  assign n10638 = ~n9715 | ~n9714;
  assign n10778 = ~n10773 | ~n10772;
  assign n14607 = ~n14727;
  assign n14100 = ~n14087 & ~n14086;
  assign n16740 = ~n16730 | ~n16731;
  assign n14744 = ~n14743 | ~n14742;
  assign n10791 = ~n15936 & ~n9770;
  assign n14209 = ~n14207 | ~n15637;
  assign n13879 = ~n13877 & ~n13876;
  assign n13942 = ~n13937 & ~n16365;
  assign n15407 = ~n15406 & ~n15405;
  assign n13963 = ~n13958 | ~n13957;
  assign n13894 = ~n13891 | ~n13890;
  assign n14474 = ~n14473 & ~n14472;
  assign n14485 = ~n14484 & ~n14483;
  assign n10773 = ~n14736 | ~n10907;
  assign n15913 = ~n15912 & ~n15911;
  assign n14771 = ~n14770;
  assign n14786 = ~n16720 | ~n16721;
  assign n14284 = ~n14283 | ~n14375;
  assign n14620 = ~n14619 & ~n14618;
  assign n13759 = ~n13758 & ~n13757;
  assign n14436 = ~n14435 & ~n14434;
  assign n14310 = ~n14309 & ~n14308;
  assign n13989 = ~n13814 | ~n13813;
  assign n13712 = ~n13711 & ~n13710;
  assign n10259 = ~n10258 | ~n10257;
  assign n14087 = ~n14283;
  assign n14606 = ~n10775 | ~n10774;
  assign n10771 = ~n10770 & ~n10769;
  assign n15277 = ~n15273 & ~n15272;
  assign n14342 = ~n14341 | ~n14340;
  assign n10607 = ~n14622;
  assign n10606 = ~n14622 | ~n16724;
  assign n15405 = ~n15404 | ~n15403;
  assign n14770 = ~n16723 & ~n16721;
  assign n13589 = ~n13588 & ~n13587;
  assign n13891 = ~n13888 & ~n13887;
  assign n13628 = ~n13625 & ~n13624;
  assign n13615 = ~n16377 | ~n13614;
  assign n13814 = ~n13810 | ~n15637;
  assign n13900 = ~n10509 | ~n10508;
  assign n13700 = ~n13753 & ~n11663;
  assign n13966 = ~n13965 & ~n13964;
  assign n10642 = ~n9710 | ~n9709;
  assign n13612 = ~n16381 | ~n13614;
  assign n13737 = ~n13740 | ~n13734;
  assign n13579 = ~n13626 & ~n13577;
  assign n13565 = ~n13564 & ~n13563;
  assign n14341 = ~n14336 | ~n16367;
  assign n15272 = ~n15271 & ~n15270;
  assign n13661 = ~n13659 & ~n13658;
  assign n13758 = ~n13753 & ~n16365;
  assign n14401 = ~n14400 & ~n14914;
  assign n13875 = ~n13888 & ~n13874;
  assign n13921 = ~n13920 | ~n13919;
  assign n13958 = ~n13954 | ~n15557;
  assign n14736 = ~n14400;
  assign n14233 = ~n15919;
  assign n13982 = ~n13981 & ~n13980;
  assign n10774 = ~n10759 | ~n10758;
  assign n15404 = ~n15395 | ~n15394;
  assign n14472 = ~n10590 & ~n16703;
  assign n16720 = ~n16723;
  assign n14435 = ~n10740 & ~n10741;
  assign n15919 = ~n15915 & ~n15916;
  assign n13888 = ~n13868 | ~n13867;
  assign n13965 = ~n13976 & ~n16431;
  assign n13962 = ~n13976 & ~n15455;
  assign n14650 = ~n14649 & ~n16703;
  assign n14333 = ~n14332 & ~n14331;
  assign n13534 = ~n13533 & ~n13532;
  assign n10759 = ~n15915 | ~n10907;
  assign n14473 = ~n10589 & ~n14641;
  assign n13669 = ~n13666 | ~n13665;
  assign n10757 = ~n10756 & ~n10755;
  assign n14231 = ~n14230 & ~n14229;
  assign n15271 = ~n15269 & ~n15268;
  assign n15910 = ~n15915 & ~n14737;
  assign n14340 = ~n14339 & ~n14338;
  assign n12976 = n10611 ^ ~n10610;
  assign n13920 = ~n13916 | ~n13915;
  assign n13626 = ~n13575 | ~n13574;
  assign n14219 = ~n14218 | ~n14217;
  assign n13625 = ~n13617 & ~n16365;
  assign n14336 = ~n14243 & ~n14195;
  assign n14447 = ~n14446 & ~n14445;
  assign n14175 = ~n14174 & ~n14173;
  assign n13740 = ~n13726 & ~n13725;
  assign n13601 = ~n13600 & ~n13599;
  assign n13751 = ~n13750 & ~n13749;
  assign n15408 = ~n15372 | ~n15371;
  assign n14218 = ~n14261 | ~n16367;
  assign n13915 = ~n13914 & ~n15479;
  assign n15269 = ~n15384 & ~n15382;
  assign n13726 = ~n13722 & ~n11752;
  assign n13657 = ~n13663 & ~n13656;
  assign n16289 = ~n16101;
  assign n15393 = ~n15384 & ~n15383;
  assign n13610 = ~n13609 & ~n13608;
  assign n10741 = ~n10739 | ~n10738;
  assign n15213 = ~n15205 & ~n15204;
  assign n14649 = ~n16702;
  assign n13666 = ~n13663 & ~n13662;
  assign n13734 = ~n13733 & ~n13732;
  assign n16107 = ~n14337 & ~n15916;
  assign n16099 = ~n16155 | ~n16058;
  assign n16706 = ~n16702 | ~n16703;
  assign n13600 = ~n13596 & ~n15617;
  assign n13868 = ~n13863 & ~n13862;
  assign n13562 = ~n13608 & ~n13561;
  assign n13575 = ~n13580 | ~n15057;
  assign n10756 = ~n14337 & ~n9770;
  assign n13988 = ~n13987 | ~n13986;
  assign n10611 = ~n9705 | ~n9704;
  assign n10573 = ~n10572 | ~n16696;
  assign n13210 = ~n13207 | ~n13206;
  assign n14496 = ~n14495 | ~n16696;
  assign n10484 = ~n10483 & ~n10482;
  assign n15204 = ~n15203 | ~n15202;
  assign n13663 = ~n13652 | ~n13651;
  assign n13449 = ~n13446 | ~n13445;
  assign n10556 = ~n10555 | ~n16676;
  assign n15384 = ~n15260 & ~n15262;
  assign n10739 = ~n14262 | ~n10907;
  assign n15383 = ~n15382 & ~n15381;
  assign n13750 = ~n13745 & ~n16356;
  assign n13479 = ~n13477 & ~n13476;
  assign n10737 = ~n10736 & ~n10735;
  assign n13699 = ~n13698 | ~n13697;
  assign n15895 = ~n15882 & ~n15881;
  assign n9705 = ~n10593 | ~n10592;
  assign n10164 = ~n10139 | ~n10138;
  assign n13733 = ~n13745 & ~n16386;
  assign n16155 = ~n14187 | ~n15887;
  assign n14487 = ~n14495 & ~n14492;
  assign n14379 = ~n14378 & ~n14377;
  assign n16291 = ~n15908;
  assign n14261 = ~n14214 & ~n14213;
  assign n13519 = ~n13516 & ~n13515;
  assign n13561 = ~n13607 & ~n13560;
  assign n10555 = ~n14162;
  assign n13985 = ~n13818 & ~n14212;
  assign n14363 = ~n16675 | ~n16676;
  assign n14489 = ~n16695 & ~n16696;
  assign n13300 = ~n13297 & ~n13296;
  assign n15382 = ~n15265 & ~n15264;
  assign n10726 = n10467 & n10466;
  assign n14723 = ~n14715 & ~n14714;
  assign n15202 = ~n15201 | ~n15394;
  assign n15260 = ~n15265 & ~n15261;
  assign n14495 = ~n16695;
  assign n10736 = ~n15902 & ~n9770;
  assign n10593 = ~n9700 | ~n9699;
  assign n13652 = ~n13644 & ~n13643;
  assign n13698 = ~n13693 | ~n15637;
  assign n13477 = ~n13469 & ~n15617;
  assign n13446 = ~n13441;
  assign n14262 = ~n15902;
  assign n10461 = ~n10460 | ~n10459;
  assign n14373 = ~n14376 & ~n14372;
  assign n14378 = ~n14376 & ~n14375;
  assign n14179 = ~n14178 | ~n14177;
  assign n15286 = ~n15285 | ~n15371;
  assign n13609 = ~n13607 & ~n16365;
  assign n15406 = ~n15380 & ~n15379;
  assign n13207 = ~n13214 | ~n14669;
  assign n15370 = ~n15369 | ~n15368;
  assign n16689 = ~n16682 & ~n16681;
  assign n14227 = ~n15902 | ~n14610;
  assign n13441 = ~n13383 | ~n13382;
  assign n13574 = ~n13573 & ~n13572;
  assign n13941 = ~n13940 | ~n13939;
  assign n14181 = ~n15880 | ~n15883;
  assign n15368 = ~n15367 | ~n15366;
  assign n13214 = ~n13193 | ~n13192;
  assign n13354 = ~n13353 & ~n13352;
  assign n13397 = ~n13394 & ~n13393;
  assign n13515 = ~n13514 | ~n13513;
  assign n9700 = ~n10577 | ~n10575;
  assign n15201 = ~n15200 | ~n15256;
  assign n13250 = ~n13247 | ~n13246;
  assign n13353 = ~n13349 & ~n15617;
  assign n10437 = ~n10436 | ~n10435;
  assign n10577 = ~n9695 | ~n9694;
  assign n13573 = ~n13570 & ~n15479;
  assign n13664 = ~n13640 & ~n13639;
  assign n13247 = ~n13245 & ~n13244;
  assign n13445 = ~n13444 & ~n13443;
  assign n13558 = ~n13557 | ~n13556;
  assign n15366 = ~n15284 | ~n15283;
  assign n13383 = ~n13375 & ~n13374;
  assign n10412 = ~n10411 & ~n10410;
  assign n14708 = ~n14706 & ~n14705;
  assign n15205 = ~n15183 & ~n15182;
  assign n15279 = ~n15255 | ~n15378;
  assign n14705 = ~n14704 & ~n15268;
  assign n13692 = ~n13691 | ~n13690;
  assign n13557 = ~n13569 | ~n13553;
  assign n14605 = ~n14597 & ~n14596;
  assign n10402 = ~n10401 & ~n10400;
  assign n15283 = ~P2_REG1_REG_17__SCAN_IN | ~n15282;
  assign n13244 = ~n13243 | ~n13242;
  assign n13179 = ~n13176 | ~n13175;
  assign n10435 = ~n10434 | ~n10433;
  assign n10411 = ~n10406 & ~n10405;
  assign n10537 = ~n10536 | ~n16669;
  assign n15375 = ~n15374 | ~n15373;
  assign n10410 = ~n10409 & ~n14129;
  assign n10545 = ~n12176 | ~n8921;
  assign n13375 = ~n13442 & ~n15455;
  assign n13442 = ~n13367 & ~n13366;
  assign n13238 = ~n13235 | ~n13234;
  assign n13809 = ~n15887;
  assign n13206 = ~n13219 & ~n13205;
  assign n16882 = ~n14372 & ~n14282;
  assign n14375 = ~n14282;
  assign n13176 = ~n13154 & ~n13153;
  assign n13387 = ~n13333 | ~n13332;
  assign n10409 = ~n10407;
  assign n13803 = ~n14059 | ~n13808;
  assign n15284 = ~n15281 | ~n15280;
  assign n15140 = ~n15131 & ~n15130;
  assign n9692 = ~n9283 | ~n9282;
  assign n10434 = ~n14059 | ~n10907;
  assign n15195 = ~n15190 | ~n15189;
  assign n10432 = ~n10431 & ~n10430;
  assign n10406 = ~n10407 & ~n10408;
  assign n10401 = ~n14130 & ~n10408;
  assign n14040 = ~n14032 & ~n14031;
  assign n15212 = ~n15378 | ~n15211;
  assign n13333 = ~n13329 & ~n13328;
  assign n15253 = ~P2_REG2_REG_17__SCAN_IN | ~n15252;
  assign n13897 = ~n10518 & ~n14074;
  assign n14769 = ~n14767 & ~n14766;
  assign n13154 = ~n13148 | ~n13147;
  assign n13219 = ~n13200 | ~n13199;
  assign n13754 = ~n13817 & ~n13705;
  assign n15130 = ~n15129 | ~n15128;
  assign n16228 = ~n15888 & ~n13808;
  assign n13235 = ~n13232 & ~n13231;
  assign n10407 = ~n10404 & ~n14125;
  assign n14714 = ~n14713 & ~n15182;
  assign n10408 = ~n10386 | ~n10385;
  assign n13175 = ~n13174 & ~n13173;
  assign n16156 = ~n15873;
  assign n13137 = ~n13134 | ~n13133;
  assign n13817 = ~n13926;
  assign n14701 = ~n14696 | ~n14695;
  assign n15873 = ~n14135 & ~n14116;
  assign n13245 = ~n13087 | ~n13086;
  assign n13800 = ~n14135 | ~n14060;
  assign n13686 = ~n16056;
  assign n13898 = ~n10517 & ~n14079;
  assign n12915 = ~n12912 | ~n12911;
  assign n10384 = ~n10383 & ~n10382;
  assign n13232 = ~n13116 | ~n13115;
  assign n15128 = ~n15127 | ~n8934;
  assign n14722 = ~n14721 | ~n15378;
  assign n16056 = ~n13797 & ~n14060;
  assign n14597 = ~n14579 & ~n15182;
  assign n13611 = ~n13606 & ~n13605;
  assign n14765 = ~n14763 & ~n14762;
  assign n12912 = ~n12905 & ~n12955;
  assign n10403 = ~n10399 | ~n10398;
  assign n14135 = ~n13797;
  assign n9278 = ~n9275 | ~n10414;
  assign n15251 = ~n15210 | ~n15209;
  assign n14471 = ~n14469 & ~n14468;
  assign n16625 = ~n16620 & ~n16619;
  assign n14711 = ~P2_REG1_REG_15__SCAN_IN | ~n14710;
  assign n13865 = ~n16875;
  assign n10397 = ~n10396 & ~n10395;
  assign n13618 = ~n13704 & ~n13582;
  assign n14767 = ~n14753 & ~n14752;
  assign n14468 = ~n14467 | ~n14466;
  assign n16603 = ~n16460 & ~n16459;
  assign n14590 = ~n14585 | ~n14584;
  assign n13688 = ~n14113 & ~n14136;
  assign n10296 = ~n10298;
  assign n13952 = ~n16642 | ~n16645;
  assign n14763 = ~n14761 & ~n14760;
  assign n10508 = ~n10507 | ~n13960;
  assign n12944 = ~n12941 | ~n12940;
  assign n13131 = ~n13003 | ~n13002;
  assign n12758 = ~n12929 | ~n12755;
  assign n13522 = ~n10279 | ~n10278;
  assign n15125 = ~n15124 | ~n15123;
  assign n10263 = ~n10075 | ~n10074;
  assign n15135 = ~n15134 | ~n15133;
  assign n14467 = ~n14465 & ~n14464;
  assign n13603 = ~n13543 | ~n13542;
  assign n10373 = ~n11804 & ~n14967;
  assign n16875 = ~n16630 | ~n16456;
  assign n13544 = ~n16062;
  assign n14712 = ~n14717 | ~n14709;
  assign n14018 = ~n14013 | ~n14012;
  assign n10075 = ~n10077;
  assign n13548 = ~n16183;
  assign n10261 = ~n10077 | ~n10076;
  assign n13380 = ~n16872;
  assign n16062 = ~n13604 | ~n15850;
  assign n16624 = ~n16623 & ~n16622;
  assign n10295 = ~n10294 | ~n10293;
  assign n15134 = ~n14751 | ~n14750;
  assign n13078 = n16181 & n16270;
  assign n15863 = ~n13604 | ~n13571;
  assign n10279 = ~n10276;
  assign n13521 = ~n10276 | ~n10277;
  assign n15123 = ~n14759 | ~n14758;
  assign n10358 = ~n10301 | ~n10300;
  assign n10237 = ~n10236 | ~n16462;
  assign n16458 = ~n16628 & ~n13730;
  assign n15853 = ~n15849 | ~n15850;
  assign n14720 = ~n14717 | ~n14716;
  assign n16059 = ~n15849 | ~n13571;
  assign n10213 = ~n10212 | ~n13634;
  assign n10074 = ~n10076;
  assign n14758 = ~n14757 | ~n14756;
  assign n13581 = ~n15849 & ~n13541;
  assign n10277 = ~n10275 | ~n10274;
  assign n16872 = ~n13364 & ~n13645;
  assign n14750 = ~n14749 | ~n14748;
  assign n13715 = ~n16622;
  assign n10394 = ~n11714 & ~n14967;
  assign n13546 = ~n15835 & ~n15836;
  assign n14748 = ~n14454 | ~n14453;
  assign n14756 = ~n14461 | ~n14460;
  assign n13190 = ~n16276;
  assign n13781 = ~n13776 | ~n13775;
  assign n10076 = ~n10073 | ~n10072;
  assign n13637 = ~n13714 & ~n16462;
  assign n10071 = ~n10070 | ~n10069;
  assign n13728 = ~n13727;
  assign n13717 = ~n16465;
  assign n10273 = ~n10272 & ~n10271;
  assign n16622 = ~n13714 & ~n13859;
  assign n15830 = ~n15818 & ~n15817;
  assign n13186 = ~n15826 | ~n15829;
  assign n13184 = ~n9687 & ~n13007;
  assign n13727 = ~n16461 & ~n13859;
  assign n16274 = ~n15819 & ~n15829;
  assign n12929 = ~n12743 & ~n12742;
  assign n13202 = ~n15819 & ~n13143;
  assign n14453 = ~n14452 | ~n14451;
  assign n10286 = ~n11615 | ~n9810;
  assign n16465 = ~n16461 & ~n16462;
  assign n10252 = ~n11615 | ~n8921;
  assign n14460 = ~n14459 | ~n14458;
  assign n16276 = ~n15839 & ~n15836;
  assign n16061 = ~n15839 | ~n15836;
  assign n13645 = ~n13635 & ~n16466;
  assign n13648 = ~n13635 | ~n16466;
  assign n14451 = ~n13836 | ~n13835;
  assign n9687 = ~n13006 & ~n13008;
  assign n13261 = ~n13256 | ~n13255;
  assign n15562 = ~n15561 & ~n15560;
  assign n14572 = ~n14430 | ~n16425;
  assign n14458 = ~n13844 | ~n13843;
  assign n14029 = ~n14034 | ~n14026;
  assign n10050 = ~n10049 & ~n13508;
  assign n16415 = ~n16414 & ~n16413;
  assign n10270 = ~n11519 & ~n14967;
  assign n15449 = ~n15448 & ~n15447;
  assign n13008 = ~n9686 & ~n12688;
  assign n10210 = ~n11435 | ~n8921;
  assign n10047 = ~n13509 & ~n10048;
  assign n10062 = ~n11435 | ~n10842;
  assign n12814 = ~n12812 | ~n12811;
  assign n16349 = ~n16348 | ~n16347;
  assign n14686 = ~n16933 | ~n14428;
  assign n13508 = ~n10048;
  assign n10202 = ~n9646 & ~n16608;
  assign n16179 = ~n16088 | ~n16270;
  assign n14037 = ~n14034 | ~n14033;
  assign n13833 = ~P1_REG2_REG_15__SCAN_IN | ~n13484;
  assign n16809 = ~n15589;
  assign n15237 = ~n15236 & ~n15235;
  assign n16870 = ~n16594 & ~n13360;
  assign n13841 = ~P1_REG1_REG_15__SCAN_IN | ~n13491;
  assign n9686 = ~n12687 & ~n12689;
  assign n13044 = ~n13039 | ~n13038;
  assign n13039 = ~n12521 | ~n12520;
  assign n10048 = ~n10046 | ~n10045;
  assign n10200 = ~n9647 & ~n16605;
  assign n12858 = ~n9992 | ~n9991;
  assign n10044 = ~n10043 | ~n10042;
  assign n16775 = ~n16779;
  assign n16597 = ~n13360 & ~n13359;
  assign n16905 = ~n13403 | ~n13402;
  assign n16088 = ~n13089 | ~n13076;
  assign n13437 = n13436 & n13435;
  assign n13425 = n13436 & n13424;
  assign n15643 = ~n15642 & ~n15641;
  assign n16779 = ~n10701 | ~n10700;
  assign n13320 = ~n13319 & ~n13318;
  assign n10501 = n10500 & n10499;
  assign n16868 = ~n16592 | ~n16586;
  assign n12521 = ~n12516 | ~n12515;
  assign n15001 = ~n15000 & ~n14999;
  assign n9685 = ~n12416 & ~n12418;
  assign n15575 = ~n15572;
  assign n13360 = ~n16610 & ~n16608;
  assign n13089 = ~n13517;
  assign n15572 = ~n10495 | ~n10494;
  assign n13064 = ~n13293 | ~n13503;
  assign n13488 = ~n12561 | ~n12560;
  assign n10012 = ~n10011 & ~n10010;
  assign n10700 = n10699 & n10698;
  assign n9992 = ~n9988 | ~n9987;
  assign n16076 = ~n13293 & ~n15803;
  assign n16866 = ~n16582 & ~n16584;
  assign n12965 = ~n9608 | ~n9607;
  assign n13290 = ~n10014 & ~n10013;
  assign n13483 = ~n13481 & ~n13480;
  assign n12516 = ~n12113 | ~n12112;
  assign n13271 = ~n13276 | ~n13268;
  assign n13011 = ~n9584 & ~n12990;
  assign n16173 = ~n12578 & ~n16078;
  assign n15669 = ~n15673;
  assign n13268 = ~n13032 | ~n13031;
  assign n12113 = ~n12108 | ~n12107;
  assign n12560 = ~n12559 | ~n12558;
  assign n9684 = ~n12078 & ~n12080;
  assign n13409 = ~n13230;
  assign n14429 = ~P2_REG3_REG_28__SCAN_IN & ~n13400;
  assign n13390 = ~n16423;
  assign n15579 = ~n16423 | ~n13744;
  assign n15446 = ~n16759;
  assign n9639 = ~n11262 | ~n8921;
  assign n13293 = ~n15802;
  assign n10495 = n10491 & n10490;
  assign n16424 = ~n12307;
  assign n13279 = ~n13276 | ~n13275;
  assign n16582 = ~n16576;
  assign n15796 = ~n12889 | ~n12900;
  assign n12572 = ~n12155 | ~n12154;
  assign n9608 = ~n9605 | ~n13410;
  assign n14781 = ~n16454 & ~n15559;
  assign n15234 = ~n15334;
  assign n12108 = ~n12015 | ~n12014;
  assign n12558 = ~n12164 | ~n12163;
  assign n16570 = ~n12991 | ~n12997;
  assign n9989 = ~n9986 | ~n9985;
  assign n9984 = ~n9983 | ~n9982;
  assign n16573 = ~n13129 | ~n13410;
  assign n9683 = ~n11902 & ~n11904;
  assign n12889 = ~n15788;
  assign n15112 = ~n15999 | ~n15533;
  assign n15334 = ~n10635 | ~n10634;
  assign n16454 = ~n15338;
  assign n16078 = ~n15772 & ~n15777;
  assign n10001 = ~n11163 & ~n14967;
  assign n12155 = ~n12153 & ~n12152;
  assign n16574 = ~n13016 | ~n12990;
  assign n10896 = ~n15495 | ~n8920;
  assign n12164 = ~n12162 & ~n12161;
  assign n13275 = ~n13056 | ~n13055;
  assign n15308 = ~n15520;
  assign n16018 = ~n10930 | ~n10929;
  assign n13029 = ~n12531 | ~n12530;
  assign n12837 = ~n9940 | ~n9939;
  assign n12015 = ~n12010 | ~n12009;
  assign n16734 = ~n10621 | ~n10620;
  assign n12530 = ~P2_REG1_REG_9__SCAN_IN | ~n12529;
  assign n12010 = ~n11864 | ~n11863;
  assign n10930 = ~n15655 | ~n8920;
  assign n12161 = ~n12160 & ~n12159;
  assign n15045 = ~n15964;
  assign n12836 = ~n9937 | ~n9938;
  assign n12152 = ~n12151 & ~n12150;
  assign n15969 = ~n15983;
  assign n16439 = ~n11892 | ~n11891;
  assign n15520 = ~n10873 | ~n10872;
  assign n15495 = ~n10889 & ~n15655;
  assign n15964 = ~n10808 | ~n10807;
  assign n16721 = ~n16724;
  assign n10620 = n10619 & n10618;
  assign n14826 = ~n15953 & ~n15639;
  assign n10889 = ~n10888 & ~P1_REG3_REG_28__SCAN_IN;
  assign n10872 = n10871 & n10870;
  assign n10718 = ~n15517 | ~n8920;
  assign n11864 = ~n11859 | ~n11858;
  assign n10828 = ~n15953 & ~n10827;
  assign n16444 = ~n11989 | ~n11535;
  assign n12531 = ~n12536 | ~n12528;
  assign n11892 = ~n11890 | ~n11889;
  assign n9682 = ~n11706 & ~n11708;
  assign n16703 = ~n14641;
  assign n10871 = ~n8920 | ~n15430;
  assign n10888 = ~n10887 & ~n10886;
  assign n16560 = ~n12810 | ~n13015;
  assign n11598 = ~n11597 & ~n11596;
  assign n11610 = ~n11504 | ~n11503;
  assign n10807 = n10806 & n10805;
  assign n9394 = ~n9393 & ~n9392;
  assign n11889 = ~n11888 | ~n11887;
  assign n15953 = ~n15949;
  assign n12440 = ~n9914 & ~n9913;
  assign n9938 = ~n9936 | ~n9935;
  assign n11987 = ~n11983 | ~n11982;
  assign n15497 = ~n15660;
  assign n11859 = ~n11563 | ~n11562;
  assign n11070 = ~n9567 | ~n9566;
  assign n12538 = ~P2_REG2_REG_9__SCAN_IN | ~n12537;
  assign n15659 = ~n15074;
  assign n14547 = ~n15323 & ~n12952;
  assign n10849 = ~n8920 | ~n15042;
  assign n15439 = ~n15515;
  assign n11986 = ~n11985 | ~n11984;
  assign n11534 = ~n11985 | ~n11531;
  assign n15937 = ~n15933;
  assign n16851 = ~n12392 | ~n12391;
  assign n15601 = ~n15342;
  assign n16553 = ~n12762 | ~n12769;
  assign n10887 = ~n10869 | ~P1_REG3_REG_26__SCAN_IN;
  assign n14641 = ~n10588 | ~n10587;
  assign n16696 = ~n14492;
  assign n11563 = ~n11630 | ~n11629;
  assign n11596 = ~n11509 | ~n11508;
  assign n12539 = ~n12536 | ~n12535;
  assign n12100 = ~n12099 | ~n12098;
  assign n11503 = ~n11502 | ~n11501;
  assign n15518 = ~n15428;
  assign n9681 = ~n11548 & ~n11550;
  assign n12535 = ~n12125 | ~n12124;
  assign n10869 = n10847 & P1_REG3_REG_25__SCAN_IN;
  assign n10821 = n10820 & n10819;
  assign n16259 = ~n12447 & ~n12847;
  assign n11630 = ~n11557 | ~n11556;
  assign n15511 = ~n15426;
  assign n11643 = ~n10129 | ~n10128;
  assign n11644 = ~n11653 & ~n10132;
  assign n15428 = ~n10142 | ~n14874;
  assign n15933 = ~n10789 | ~n10788;
  assign n15094 = ~n10146 | ~n11686;
  assign n16548 = ~n12765 | ~n12761;
  assign n12364 = ~n12447 & ~n12375;
  assign n15167 = ~n14873;
  assign n11886 = ~n9388 & ~n9387;
  assign n11550 = ~n9680 & ~n11390;
  assign n9399 = ~n9398 & ~n9397;
  assign n11533 = ~n11984 | ~n11532;
  assign n11508 = ~n11296 | ~n11295;
  assign n11501 = ~n11305 | ~n11304;
  assign n15342 = ~n9657 | ~n11990;
  assign n9398 = ~n11888 & ~n9395;
  assign n11557 = ~n11553 | ~n11552;
  assign n16631 = ~n13730;
  assign n11296 = ~n11294 & ~n11293;
  assign n12435 = ~n9891 & ~n9890;
  assign n14611 = ~n10768 | ~n10767;
  assign n9649 = ~n9390 | ~n9650;
  assign n11890 = ~n11885 | ~n11884;
  assign n11304 = ~n11303 & ~n11302;
  assign n12006 = ~P2_REG1_REG_7__SCAN_IN | ~n12005;
  assign n16542 = ~n12675 & ~n12407;
  assign n10788 = n10787 & n10786;
  assign n15455 = ~n16410;
  assign n15426 = ~n10144 | ~n10123;
  assign n9680 = ~n11389 & ~n11391;
  assign n10847 = n10804 & P1_REG3_REG_24__SCAN_IN;
  assign n11834 = ~n11833 | ~n11832;
  assign n11391 = ~n9679 & ~n9678;
  assign n11990 = ~n16358;
  assign n11302 = ~n11301 & ~n11300;
  assign n15028 = ~n16038 & ~n15640;
  assign n12007 = ~n12020 | ~n12004;
  assign P1_U3085 = ~n9020 | ~P1_STATE_REG_SCAN_IN;
  assign n11553 = ~n11428 & ~n9168;
  assign n11293 = ~n11292 & ~n11291;
  assign n14610 = ~n15901;
  assign n11786 = ~n16475 | ~n16479;
  assign n9364 = ~n11888 | ~n16960;
  assign n16540 = ~n12793 & ~n12467;
  assign n16482 = ~n16475;
  assign n16665 = ~n10534 | ~n10533;
  assign n9527 = ~n9513 | ~n8921;
  assign n11884 = ~n11883 | ~n11997;
  assign n13730 = ~n10180 & ~n10179;
  assign n10767 = n10766 & n10765;
  assign n14737 = ~n15916;
  assign n10804 = n10818 & P1_REG3_REG_23__SCAN_IN;
  assign n9389 = ~n11524 | ~n11531;
  assign n13101 = ~n9363 & ~n9362;
  assign n13694 = ~n14136;
  assign n10818 = n10785 & P1_REG3_REG_22__SCAN_IN;
  assign n13023 = ~n9604 & ~n9603;
  assign n16960 = ~n11997 & ~n10958;
  assign n15916 = ~n10754 | ~n10753;
  assign n16065 = ~n15715 & ~n12038;
  assign n11763 = ~n11762 & ~n11761;
  assign n12900 = ~n15789;
  assign n11301 = ~n11193 | ~n11277;
  assign n15836 = ~n15840;
  assign n11292 = ~n11210 & ~n11209;
  assign n9383 = ~n9382 | ~n9384;
  assign n9387 = ~n9650 & ~n9386;
  assign n13571 = ~n15850;
  assign n9678 = ~n11172 & ~n11171;
  assign n14079 = ~n10172 | ~n10171;
  assign n15564 = ~n13871 | ~n14685;
  assign n12022 = ~P2_REG2_REG_7__SCAN_IN | ~n12021;
  assign n11835 = ~n11655 | ~n11660;
  assign n11883 = ~n9650;
  assign n11661 = ~n11674;
  assign n15557 = ~n11752;
  assign n15901 = ~n10477 | ~n10476;
  assign n11832 = ~n10984 & ~n11674;
  assign n11428 = ~n11426 & ~n11425;
  assign n11172 = ~n9677 & ~n9676;
  assign n12023 = ~n12020 | ~n12019;
  assign n16133 = ~n11081 | ~n11080;
  assign n11209 = ~n11273 & ~n11272;
  assign n11982 = ~n11984 & ~n16591;
  assign n11426 = ~n9160 | ~n9159;
  assign n16313 = ~n11105 & ~n11104;
  assign n13808 = ~n10429 | ~n10428;
  assign n10546 = ~n10527 | ~n14047;
  assign n14177 = ~n10458 & ~n10457;
  assign n15850 = ~n10292 | ~n10291;
  assign n10123 = ~n10984 & ~n10131;
  assign n13283 = ~n10041 & ~n10040;
  assign n10785 = n10764 & P1_REG3_REG_21__SCAN_IN;
  assign n12407 = ~n9498 & ~n9497;
  assign n11855 = ~n11854 | ~n11853;
  assign n11277 = ~n11275 | ~n11276;
  assign n15654 = ~n14874;
  assign n10827 = ~n10906;
  assign n10653 = ~n10652 & ~n10651;
  assign n10634 = ~n10633 & ~n10632;
  assign n10604 = ~n10603 & ~n10602;
  assign n10587 = ~n10586 & ~n10585;
  assign n10561 = ~n10560 | ~n10559;
  assign n10569 = ~n10568 & ~n10567;
  assign n10674 = ~n10673 & ~n10672;
  assign n10552 = ~n10551 & ~n10550;
  assign n10525 = ~n10524 | ~n10523;
  assign n10527 = ~P2_REG3_REG_16__SCAN_IN & ~n10488;
  assign n10533 = ~n10532 & ~n10531;
  assign n10515 = ~n10514 | ~n10513;
  assign n10171 = ~n10170 & ~n10169;
  assign n10192 = ~n10191 | ~n10190;
  assign n10224 = ~n10223 | ~n10222;
  assign n9638 = ~n9637 & ~n9636;
  assign n10764 = n10747 & P1_REG3_REG_20__SCAN_IN;
  assign n11984 = ~n11531;
  assign n14874 = ~n11658 | ~n11654;
  assign n11272 = ~n11481 | ~n11208;
  assign n15182 = ~n15371;
  assign n9676 = ~n11077 & ~n11076;
  assign n11275 = ~n11486 | ~n11192;
  assign n11077 = ~n9675 & ~n9674;
  assign n11891 = ~n10958;
  assign n10747 = n10711 & P1_REG3_REG_19__SCAN_IN;
  assign n16345 = ~n16411;
  assign n10251 = ~n10250 & ~n10249;
  assign n13769 = ~P2_REG1_REG_12__SCAN_IN | ~n13789;
  assign n10488 = ~n10184 | ~n10166;
  assign n11574 = ~P2_REG1_REG_5__SCAN_IN | ~n11626;
  assign n10544 = ~n10543 & ~n10542;
  assign n15371 = ~n11322 & ~n15386;
  assign n9385 = ~n11751;
  assign n11875 = ~n11874 | ~n11873;
  assign n10131 = ~n15536 | ~n11667;
  assign n11873 = ~n11588 | ~n11587;
  assign n13276 = ~n13258;
  assign n10579 = ~n8933 & ~n10578;
  assign n10269 = ~n10268 | ~n10267;
  assign n10595 = ~n8933 & ~n10594;
  assign n10421 = ~n10420 | ~n10419;
  assign n11575 = ~n11585 | ~n11573;
  assign n16346 = ~n15559;
  assign n10711 = ~n10470 & ~n10478;
  assign n11322 = ~n9101 | ~n9089;
  assign n16365 = ~n15103;
  assign n10613 = ~n8933 & ~n10612;
  assign n10733 = ~n10732 | ~n10731;
  assign n9674 = ~n11025 & ~n11024;
  assign n10644 = ~n8933 & ~n10643;
  assign n10028 = ~n10027 & ~n10026;
  assign n15536 = ~n16369;
  assign n10393 = ~n10392 | ~n10391;
  assign n13789 = ~n13779;
  assign n11025 = ~n9673 | ~n9672;
  assign n11573 = ~n11572 | ~n11571;
  assign n10228 = ~n10165 | ~n13470;
  assign n8925 = ~n16918;
  assign n10470 = ~n10452 | ~P1_REG3_REG_17__SCAN_IN;
  assign n11754 = ~n11539;
  assign n10285 = ~n10284 & ~n10283;
  assign n10671 = ~n13431;
  assign n13258 = ~n9634 & ~n9633;
  assign n9089 = ~n9098 & ~P2_U3151;
  assign n11587 = ~P2_REG2_REG_5__SCAN_IN | ~n11636;
  assign n16367 = ~n15534;
  assign n8927 = ~n10005;
  assign n10061 = ~n10060 & ~n10059;
  assign n11662 = ~n10904;
  assign n9973 = ~n9972 & ~n9971;
  assign n15479 = ~n15637;
  assign n15584 = ~n8921;
  assign n10450 = ~n10449 & ~n10448;
  assign n10962 = ~n10116 & ~n10114;
  assign n11588 = ~n11585 | ~n11586;
  assign n10116 = ~n13460;
  assign n11554 = ~n9170 | ~n9169;
  assign n16146 = ~n11667;
  assign n11560 = ~n11559 | ~n11558;
  assign n12517 = ~n12115 | ~n12114;
  assign n11572 = ~n11569 | ~n11568;
  assign n13040 = ~n12523 | ~n12522;
  assign n12109 = ~n12017 | ~n12016;
  assign n9755 = ~n14005;
  assign n10452 = n10425 & P1_REG3_REG_16__SCAN_IN;
  assign n12011 = ~n11866 | ~n11865;
  assign n11860 = ~n11565 | ~n11564;
  assign n9633 = ~n9632 & ~n9631;
  assign n11569 = ~n9137 | ~n9136;
  assign n10966 = ~n9671 & ~n9670;
  assign n11537 = ~n14685 & ~n16591;
  assign n10425 = ~n10375 & ~n10374;
  assign n11586 = ~n11584 | ~n11583;
  assign n10226 = ~n9368 | ~n9367;
  assign n9002 = ~n9322 | ~n9738;
  assign n9323 = ~n9322 & ~n9738;
  assign n14685 = ~n16433;
  assign n12101 = ~P2_REG1_REG_8__SCAN_IN | ~n12121;
  assign n10239 = ~n9249 & ~n9250;
  assign n9261 = ~n9260;
  assign n9242 = ~n9241;
  assign n9137 = ~n11416 | ~P2_REG1_REG_3__SCAN_IN;
  assign n10024 = ~n10022 | ~P1_IR_REG_31__SCAN_IN;
  assign n9564 = ~n9197 | ~n9196;
  assign n10375 = ~n10151 | ~P1_REG3_REG_13__SCAN_IN;
  assign n9271 = ~n9270;
  assign n9628 = ~n9221 & ~n9223;
  assign n9251 = ~n9250;
  assign n11584 = ~n11581 | ~n11580;
  assign n12125 = ~P2_REG2_REG_8__SCAN_IN | ~n12121;
  assign n9224 = ~n9223;
  assign n10053 = ~n9231 & ~n9232;
  assign n16956 = ~n13119;
  assign n9620 = ~n9616 | ~n9615;
  assign n9733 = ~n10321 | ~n9732;
  assign n9610 = ~n9213 | ~n9212;
  assign n9233 = ~n9232;
  assign n9196 = ~n9195 | ~SI_8_;
  assign n12121 = ~n12110;
  assign n9384 = ~n16961;
  assign n9380 = ~n9366 | ~n9365;
  assign n10151 = ~n10150 & ~n10149;
  assign n10322 = ~n10321;
  assign n9223 = ~n9220 & ~SI_11_;
  assign n9212 = ~n9211 | ~SI_10_;
  assign n9136 = ~n9135 | ~n9450;
  assign n11581 = ~n9150 | ~n9149;
  assign n9232 = ~n9230 & ~SI_12_;
  assign n11211 = ~n11299;
  assign n9616 = ~n9614 | ~P2_IR_REG_10__SCAN_IN;
  assign n12536 = ~n12518;
  assign n10955 = ~n9669 & ~n9668;
  assign n11856 = ~P2_REG1_REG_6__SCAN_IN | ~n11872;
  assign n9065 = ~n9064 | ~SI_3_;
  assign n11876 = ~P2_REG2_REG_6__SCAN_IN | ~n11872;
  assign n9724 = ~n9723 | ~SI_25_;
  assign n9184 = ~n9183 | ~SI_6_;
  assign n9709 = ~n9708 | ~SI_22_;
  assign n9920 = ~n9919 | ~P1_IR_REG_31__SCAN_IN;
  assign n9731 = ~n9730;
  assign n9203 = ~n9202 | ~SI_9_;
  assign n9179 = ~n9178 | ~SI_5_;
  assign n9197 = ~n9194 | ~n9193;
  assign n9150 = ~n11419 | ~P2_REG2_REG_3__SCAN_IN;
  assign n9189 = ~n9188 | ~SI_7_;
  assign n9719 = ~n9718 | ~SI_24_;
  assign n9135 = ~n9133 | ~n9132;
  assign n10021 = ~n9997 | ~P1_IR_REG_31__SCAN_IN;
  assign n9070 = ~n9069 | ~SI_4_;
  assign n9258 = ~n9257;
  assign n9231 = ~n9229 & ~n9228;
  assign n9230 = ~n9229;
  assign n9619 = ~n9617;
  assign n9249 = ~n9247 & ~n9246;
  assign n10332 = ~n10331 | ~SI_28_;
  assign n9268 = ~n9267;
  assign n9694 = ~n9693 | ~SI_19_;
  assign n9239 = ~n9238;
  assign n9248 = ~n9247;
  assign n10150 = ~n10035 | ~P1_REG3_REG_11__SCAN_IN;
  assign n9240 = ~n9238 & ~n9237;
  assign n10414 = n9276 ^ SI_17_;
  assign n9221 = ~n9219 & ~n9218;
  assign n10337 = ~n10336 | ~SI_29_;
  assign n9699 = ~n9698 | ~SI_20_;
  assign n9133 = ~n9131 | ~n9130;
  assign n9229 = ~n9227 & ~n9226;
  assign n9219 = ~n9217 & ~n9216;
  assign n9149 = ~n9148 | ~n9450;
  assign n9188 = ~n9187 | ~n9186;
  assign n10035 = ~n10032 & ~n11308;
  assign n9194 = ~n9192 & ~n9191;
  assign n9183 = ~n9182 | ~n9181;
  assign n9178 = ~n9045 | ~n9044;
  assign n11872 = ~n9523 | ~n9590;
  assign n9997 = ~n9996 | ~n9995;
  assign n9523 = ~n9519 | ~n9518;
  assign n9727 = ~n10345 & ~n13461;
  assign n9728 = n10345 & P1_DATAO_REG_26__SCAN_IN;
  assign n9356 = ~n9598 & ~P2_REG3_REG_9__SCAN_IN;
  assign n9569 = ~n9590 & ~P2_IR_REG_7__SCAN_IN;
  assign n9996 = ~n9968 & ~P1_IR_REG_8__SCAN_IN;
  assign n9696 = ~n10345 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n14154 = ~n13123;
  assign n13679 = ~n10345 | ~P2_U3151;
  assign n9544 = ~n9590 | ~P2_IR_REG_31__SCAN_IN;
  assign n9217 = ~n10345 & ~n10025;
  assign n9284 = ~n10345 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n9273 = ~n10345 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n9148 = ~n9147 | ~n9146;
  assign n11568 = ~n11567;
  assign n9131 = ~n9095 | ~n9094;
  assign n13683 = ~n14356;
  assign n11583 = ~n11582 | ~P2_REG2_REG_4__SCAN_IN;
  assign n9264 = ~n10345 & ~n9263;
  assign n10388 = ~n10281 | ~P1_IR_REG_31__SCAN_IN;
  assign n11571 = ~n11582 | ~P2_REG1_REG_4__SCAN_IN;
  assign n10324 = ~n10345 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n9598 = ~n9551 | ~n9354;
  assign n9280 = ~n10344 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n13123 = ~n10344 | ~P1_U3086;
  assign n10002 = ~n9975 & ~n11280;
  assign n9707 = ~n10344 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n9590 = ~n9522 | ~n9521;
  assign n9761 = ~n9287 | ~n8951;
  assign n9067 = ~n9043 | ~P2_DATAO_REG_4__SCAN_IN;
  assign n9968 = ~n9943 | ~n9942;
  assign n9702 = ~n10344 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n9712 = ~n10344 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n9519 = ~n9517 | ~P2_IR_REG_6__SCAN_IN;
  assign n9717 = ~n10344 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n9054 = ~n9043 & ~n9431;
  assign n9285 = ~n10344 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n9697 = ~n10344 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n9943 = ~n9893 & ~P1_IR_REG_5__SCAN_IN;
  assign n9551 = ~n9552 & ~P2_REG3_REG_7__SCAN_IN;
  assign n9287 = ~n10265 & ~n8950;
  assign n9132 = ~n11002 | ~P2_REG1_REG_2__SCAN_IN;
  assign n9975 = ~n9950 | ~P1_REG3_REG_7__SCAN_IN;
  assign n11344 = ~n9092 | ~n9094;
  assign n9520 = ~n9516 | ~n9515;
  assign n9552 = ~n9501 | ~n9353;
  assign n9950 = ~n9925 & ~n11249;
  assign n9925 = ~n9898 | ~P1_REG3_REG_5__SCAN_IN;
  assign n9031 = ~n9026 & ~P2_ADDR_REG_19__SCAN_IN;
  assign n9501 = ~n9502 & ~P2_REG3_REG_5__SCAN_IN;
  assign n9336 = ~n9335 | ~n9334;
  assign n9749 = ~n9748 | ~P1_IR_REG_31__SCAN_IN;
  assign n9008 = ~n10417 & ~P1_IR_REG_21__SCAN_IN;
  assign n8990 = ~n8989 | ~n8993;
  assign n8995 = ~n8994 | ~n8993;
  assign n8961 = ~n8963 | ~P1_IR_REG_31__SCAN_IN;
  assign n9502 = ~n9352 | ~n12301;
  assign n9078 = ~P2_IR_REG_22__SCAN_IN;
  assign n10374 = ~P1_REG3_REG_14__SCAN_IN | ~P1_REG3_REG_15__SCAN_IN;
  assign n10478 = ~P1_REG3_REG_18__SCAN_IN;
  assign n10417 = ~P1_IR_REG_31__SCAN_IN;
  assign n8951 = ~P1_IR_REG_19__SCAN_IN;
  assign n10445 = ~P1_IR_REG_18__SCAN_IN;
  assign n9084 = ~P2_IR_REG_26__SCAN_IN;
  assign n10520 = ~P2_IR_REG_31__SCAN_IN;
  assign n10282 = ~P2_DATAO_REG_14__SCAN_IN;
  assign n10489 = ~P2_REG3_REG_19__SCAN_IN;
  assign n14047 = ~P2_REG3_REG_17__SCAN_IN;
  assign n10166 = ~P2_REG3_REG_15__SCAN_IN;
  assign n9662 = ~P1_ADDR_REG_19__SCAN_IN;
  assign n8954 = ~P1_IR_REG_23__SCAN_IN;
  assign n8964 = ~P1_IR_REG_19__SCAN_IN & ~P1_IR_REG_25__SCAN_IN;
  assign n9025 = ~P1_RD_REG_SCAN_IN;
  assign n9631 = ~P2_IR_REG_11__SCAN_IN;
  assign n9882 = ~P1_REG3_REG_4__SCAN_IN | ~P1_REG3_REG_3__SCAN_IN;
  assign n9618 = ~P2_IR_REG_10__SCAN_IN;
  assign n9027 = ~P2_RD_REG_SCAN_IN;
  assign n8984 = ~P2_IR_REG_17__SCAN_IN & ~P2_IR_REG_16__SCAN_IN;
  assign n8983 = ~P2_IR_REG_14__SCAN_IN & ~P2_IR_REG_15__SCAN_IN;
  assign n8985 = ~P2_IR_REG_19__SCAN_IN & ~P2_IR_REG_18__SCAN_IN;
  assign n9028 = ~P2_ADDR_REG_19__SCAN_IN;
  assign n9006 = ~P1_IR_REG_21__SCAN_IN;
  assign n11267 = ~P2_DATAO_REG_12__SCAN_IN;
  assign n16967 = ~n16957 | ~n16956;
  assign n16957 = ~n16955 | ~n16954;
  assign n16393 = ~n16394 | ~n16438;
  assign n16922 = ~n16848 | ~n16847;
  assign n16364 = ~n16352 | ~n16351;
  assign n16396 = ~n16394 | ~n16442;
  assign n15633 = ~n15631 | ~n16442;
  assign n16848 = n16846 ^ ~n16845;
  assign n15630 = ~n15631 | ~n16438;
  assign n16437 = ~n16418 & ~n16417;
  assign n15667 = ~n15666 & ~n15665;
  assign n15508 = ~n15494 | ~n15493;
  assign n15549 = ~n15547 | ~n16381;
  assign n15546 = ~n15547 | ~n16377;
  assign n16152 = ~n16044 & ~n16043;
  assign n16376 = ~n15650 & ~n15649;
  assign n15563 = ~n15558 | ~n15557;
  assign n16404 = ~n16399 | ~n16398;
  assign n15494 = ~n15544 | ~n13226;
  assign n15476 = ~n15474 | ~n16442;
  assign n16952 = ~n16951 | ~n8925;
  assign n16325 = n16323 ^ ~n8924;
  assign n15473 = ~n15474 | ~n16438;
  assign n15514 = ~n15512 | ~n15511;
  assign n16833 = ~n16828;
  assign n16213 = ~n16212 | ~n16211;
  assign n15420 = ~n15421 | ~n16381;
  assign n16323 = ~n16321 & ~n16320;
  assign n15423 = ~n15421 | ~n16377;
  assign n15513 = ~n15510 & ~n15509;
  assign n15085 = ~n15082 & ~n15081;
  assign n15118 = ~n15116 | ~n16377;
  assign n15441 = ~n15438 & ~n15437;
  assign n16828 = ~n16815 | ~n16814;
  assign n16416 = ~n16422 | ~n16410;
  assign n15648 = ~n15647 | ~n15646;
  assign n15115 = ~n15116 | ~n16381;
  assign n15542 = ~n15532 & ~n16365;
  assign n15033 = ~n15034 | ~n16377;
  assign n15492 = ~n15486 | ~n15485;
  assign n15036 = ~n15034 | ~n16381;
  assign n15457 = ~n15450 | ~n15449;
  assign n16390 = ~n16389 & ~n16388;
  assign n15292 = ~n15289 & ~n15288;
  assign n15438 = ~n15427 & ~n15426;
  assign n15418 = ~n15416 & ~n15415;
  assign n15486 = ~n15483 | ~n15635;
  assign n16842 = ~n16835 | ~n16834;
  assign n14986 = ~n14987 | ~n16381;
  assign n16389 = ~n16387 & ~n16386;
  assign n14687 = ~n16936 | ~n14685;
  assign n16034 = ~n16033 | ~n16032;
  assign n14989 = ~n14987 | ~n16377;
  assign n15031 = ~n15027 | ~n16367;
  assign n14980 = ~n15027 | ~n15659;
  assign n15030 = ~n15029 & ~n15028;
  assign n15010 = ~n15021 | ~n16419;
  assign n15320 = ~n15414 & ~n11663;
  assign n15321 = ~n15319 | ~n15318;
  assign n16409 = ~n16406 & ~n16900;
  assign n16841 = ~n16912 | ~n16925;
  assign n16797 = ~n16807;
  assign n16813 = ~n16807 | ~n16806;
  assign n15110 = ~n15109 | ~n15108;
  assign n16929 = ~n16928 | ~n16927;
  assign n15238 = ~n15233 | ~n15557;
  assign n16033 = ~n16031;
  assign n16373 = ~n16372 | ~n16371;
  assign n16830 = ~n16820 | ~n16819;
  assign n16831 = ~n16829;
  assign n14983 = ~n14982 & ~n15028;
  assign n14984 = ~n14981 | ~n16367;
  assign n15008 = ~n15002 | ~n15001;
  assign n15080 = ~n15104 | ~n15070;
  assign n14888 = ~n14887 & ~n14886;
  assign n15164 = ~n15158 & ~n15157;
  assign n14906 = ~n14981 | ~n15659;
  assign n16914 = ~n16926 | ~n16913;
  assign n15627 = ~n15626 | ~n15625;
  assign n16928 = ~n16926 | ~n16925;
  assign n15580 = ~n15626 | ~n15579;
  assign n16935 = ~n16934 | ~n16933;
  assign n15600 = ~n15618;
  assign n15470 = ~n15469 & ~n15468;
  assign n16368 = ~n15658 & ~n15657;
  assign n15089 = ~n15157 & ~n15156;
  assign n15336 = ~n15332 & ~n15331;
  assign n14960 = ~n14959 & ~n14958;
  assign n10917 = n10911 ^ n10910;
  assign n16308 = ~n16128 & ~n16127;
  assign n16822 = ~n16906 | ~n16798;
  assign n16923 = ~n16818 | ~n16801;
  assign n14974 = ~n16134 | ~n15658;
  assign n16819 = ~n16818 | ~n16817;
  assign n16899 = ~n16898 | ~n16897;
  assign n10911 = n10905 ^ ~n10904;
  assign n10915 = ~n10920 | ~n15511;
  assign n16214 = ~n15477 | ~n15634;
  assign n15464 = ~n15467 & ~n16423;
  assign n15456 = ~n15467 & ~n15455;
  assign n14852 = ~n14867 | ~n16419;
  assign n16927 = ~n16802 | ~n16817;
  assign n10921 = ~n10920 & ~n15426;
  assign n14784 = ~n14798 | ~n16419;
  assign n16426 = ~n16802 | ~n16424;
  assign n15661 = ~n16370 | ~n15660;
  assign n14951 = ~n14954 & ~n15653;
  assign n16132 = ~n16130 | ~n16370;
  assign n14879 = ~n14877 & ~n15323;
  assign n16371 = ~n16370 | ~n16369;
  assign n16788 = ~n16787 | ~n16786;
  assign n15577 = ~n15574 | ~n16782;
  assign n16897 = ~n16896 & ~n16895;
  assign n15657 = ~n15656 & ~n16011;
  assign n14838 = ~n14837 | ~n14836;
  assign n15634 = ~n16128;
  assign n16226 = ~n16049 & ~n16048;
  assign n14009 = ~n16400 | ~n14154;
  assign n15424 = n10879 ^ n10880;
  assign n16786 = ~n16785 | ~n16784;
  assign n15996 = ~n15679 | ~n15678;
  assign n15978 = ~n15977 | ~n15976;
  assign n14940 = ~n14939 | ~n14938;
  assign n14850 = ~n14846 & ~n11752;
  assign n16769 = ~n16768 | ~n16767;
  assign n16812 = ~n16811 | ~n16810;
  assign n15291 = ~n15290 | ~n15625;
  assign n16360 = ~n16407 | ~n16424;
  assign n14782 = ~n14780 | ~n14779;
  assign n16207 = ~n16206 & ~n16205;
  assign n10932 = ~n15674 | ~n15428;
  assign n10914 = n10723 ^ ~n10904;
  assign n15249 = ~n15290 | ~n15579;
  assign n14004 = ~n16400 | ~n14351;
  assign n14885 = ~n14880 | ~n15070;
  assign n15299 = ~n15997 | ~n15298;
  assign n15498 = ~n15670 & ~n15497;
  assign n15537 = ~n15670 & ~n15536;
  assign n15598 = ~n15595;
  assign n16049 = ~n15673 & ~n15670;
  assign n10879 = n10876 ^ ~n10904;
  assign n15590 = ~n16808 & ~n16809;
  assign n16388 = ~n16808 & ~n16433;
  assign n10723 = ~n10722 | ~n10721;
  assign n14897 = ~n14894 & ~n14967;
  assign n15105 = ~n15298 | ~n15073;
  assign n14780 = ~n14778 | ~n15557;
  assign n15994 = ~n15999 & ~n16001;
  assign n15020 = ~n15019 & ~n15018;
  assign n16002 = ~n16047 | ~n16000;
  assign n15612 = ~n16808 & ~n15601;
  assign n15014 = ~n15017 & ~n16423;
  assign n16354 = ~n16778 | ~n16775;
  assign n14647 = ~n14663 | ~n16419;
  assign n15106 = ~n15309 & ~n15536;
  assign n14666 = ~n14663 | ~n14662;
  assign n15037 = ~n10862 & ~n10861;
  assign n14567 = ~n14670 | ~n14547;
  assign n15496 = ~n15519 | ~n15071;
  assign n16047 = ~n15998 | ~n15997;
  assign n15488 = ~n15999 | ~n15997;
  assign n10880 = ~n10878 | ~n10877;
  assign n10876 = ~n10875 | ~n10874;
  assign n15550 = ~n15576 | ~n15572;
  assign n15073 = ~n15429 | ~n15072;
  assign n13998 = ~n10333 | ~n10332;
  assign n15525 = ~n15519 & ~n15518;
  assign n15489 = ~n15998 | ~n15519;
  assign n15436 = ~n15429 | ~n15428;
  assign n15410 = ~n15519 & ~n15536;
  assign n15300 = ~n15519 & ~n15497;
  assign n10878 = ~n15429 | ~n10907;
  assign n10875 = ~n15429 | ~n10901;
  assign n14663 = ~n14645 & ~n14644;
  assign n16297 = ~n16122 | ~n16121;
  assign n14521 = ~n14518 | ~n14517;
  assign n14554 = ~n14677 & ~n15323;
  assign n10862 = ~n10857 & ~n10858;
  assign n15452 = ~n16910;
  assign n14422 = ~n14524 | ~n14547;
  assign n14505 = ~n14518 | ~n16419;
  assign n15989 = ~n15988 | ~n15987;
  assign n14678 = ~n14677 & ~n14676;
  assign n16205 = ~n16204 | ~n16203;
  assign n14546 = ~n14544 & ~n14543;
  assign n15988 = ~n15986 | ~n15985;
  assign n14486 = ~n14476 | ~n15596;
  assign n16122 = ~n16120 | ~n16119;
  assign n14931 = ~n14930 | ~n14929;
  assign n16296 = ~n16120 | ~n16055;
  assign n14318 = ~n14315 | ~n14314;
  assign n13465 = ~n13459 | ~n14154;
  assign n14677 = ~n14552 | ~n14551;
  assign n10857 = n10854 ^ ~n10904;
  assign n15973 = ~n15987 & ~n15972;
  assign n14518 = ~n14503 & ~n14502;
  assign n10854 = ~n10853 | ~n10852;
  assign n15986 = ~n15984 & ~n15983;
  assign n15288 = ~n15442 & ~n16433;
  assign n15058 = ~n16054;
  assign n16752 = ~n16450 | ~n16449;
  assign n14411 = ~n14529 & ~n15323;
  assign n14371 = ~n14392 | ~n16419;
  assign n14256 = ~n14307 | ~n14547;
  assign n14883 = ~n14881 & ~n15074;
  assign n14348 = ~n14345 | ~n14344;
  assign n15241 = ~n15442 & ~n15564;
  assign n15230 = ~n16759 & ~n15442;
  assign n14395 = ~n14392 | ~n14391;
  assign n15985 = ~n15981 | ~n15980;
  assign n16120 = ~n16054 & ~n16053;
  assign n10856 = ~n15968 | ~n10907;
  assign n14205 = ~n14335 | ~n14547;
  assign n10853 = ~n15968 | ~n10901;
  assign n16744 = ~n16743 | ~n16742;
  assign n14224 = ~n14257 | ~n14221;
  assign n14259 = ~n14257 | ~n13226;
  assign n14945 = ~n14944 | ~n15968;
  assign n15984 = ~n15968;
  assign n14292 = ~n14295 | ~n14289;
  assign n14392 = ~n14369 & ~n14368;
  assign n14824 = ~n14822 | ~n14821;
  assign n14298 = ~n14295 | ~n16419;
  assign n14529 = ~n14409 | ~n14408;
  assign n14334 = ~n14324 | ~n15596;
  assign n10656 = ~n15334 | ~n15333;
  assign n10832 = ~n15086;
  assign n10659 = ~n15334 | ~n10660;
  assign n16754 = ~n15334 | ~n15227;
  assign n15159 = ~n10813 | ~n10812;
  assign n15968 = ~n10844 | ~n10843;
  assign n16760 = ~n10679 | ~n10678;
  assign n15018 = ~n15227 & ~n16433;
  assign n16749 = ~n16748 & ~n16747;
  assign n16201 = ~n16200 | ~n16199;
  assign n14295 = ~n14286 & ~n14285;
  assign n10729 = ~n10727 | ~n10726;
  assign n10830 = ~n15086 & ~n15088;
  assign n16743 = ~n16739 | ~n16738;
  assign n16051 = ~n15166 | ~n15964;
  assign n14257 = ~n14211 & ~n14210;
  assign n14092 = ~n14093 | ~n16438;
  assign n15344 = ~n15343 | ~n15342;
  assign n14833 = ~n15965 | ~n16369;
  assign n14831 = ~n15965 | ~n14830;
  assign n14176 = ~n14165 | ~n15596;
  assign n13453 = ~n13452;
  assign n10844 = ~n13452 | ~n10842;
  assign n14925 = ~n15965 & ~n15964;
  assign n10813 = ~n15965 | ~n10907;
  assign n16748 = ~n16746;
  assign n13313 = ~n13452 | ~n14154;
  assign n14511 = ~n14514 & ~n16423;
  assign n14270 = ~n14260 & ~n15653;
  assign n14184 = ~n14183 | ~n14227;
  assign n15086 = n10825 ^ ~n10904;
  assign n14194 = ~n14343 & ~n15323;
  assign n10810 = ~n15965 | ~n10901;
  assign n14817 = ~n15948 | ~n15949;
  assign n13994 = ~n13991 | ~n13990;
  assign n16738 = ~n16737 | ~n16736;
  assign n14418 = ~n14525 | ~n15659;
  assign n14557 = ~n15948 | ~n14555;
  assign n14232 = ~n14228 | ~n14227;
  assign n15940 = ~n15943 | ~n15942;
  assign n14093 = ~n14096 | ~n14090;
  assign n10655 = ~n15329 | ~n15338;
  assign n14069 = ~n14057 | ~n15511;
  assign n14785 = ~n14651 & ~n14650;
  assign n15951 = ~n15948 & ~n16021;
  assign n14501 = ~n14506 | ~n16410;
  assign n15088 = ~n10829 & ~n10828;
  assign n10825 = ~n10824 & ~n10823;
  assign n16115 = ~n15952 & ~n15949;
  assign n13302 = ~n13301;
  assign n13827 = ~n13984 | ~n14547;
  assign n15219 = ~n16453 & ~n15601;
  assign n14790 = ~n14789 | ~n14788;
  assign n14731 = ~n14729;
  assign n10801 = ~n13301 | ~n9810;
  assign n15100 = ~n15952 & ~n15518;
  assign n13925 = ~n13944 | ~n13226;
  assign n14819 = ~n15952 | ~n15953;
  assign n14054 = ~n14044 | ~n15596;
  assign n14404 = ~n14403 | ~n16055;
  assign n14830 = ~n15952 | ~n14556;
  assign n10677 = ~n9720 | ~n9719;
  assign n14246 = ~n14245 | ~n13226;
  assign n13971 = ~n13969 | ~n16438;
  assign n14991 = ~n16453;
  assign n15004 = ~n15338 | ~n16453;
  assign n13947 = ~n13944 | ~n13943;
  assign n14561 = ~n15952 & ~n15497;
  assign n14864 = ~n16453 & ~n16433;
  assign n14809 = ~n16735 | ~n15342;
  assign n15942 = ~n15939 | ~n15938;
  assign n13301 = n10638 ^ ~n10637;
  assign n15925 = ~n15924 & ~n15923;
  assign n14526 = ~n15932 | ~n16369;
  assign n13944 = ~n13922 & ~n13921;
  assign n14182 = ~n14180 | ~n14179;
  assign n15935 = ~n15932 & ~n16021;
  assign n13969 = ~n13972 | ~n13966;
  assign n14304 = ~n14299 & ~n16423;
  assign n14729 = ~n10779 & ~n10778;
  assign n16741 = ~n16733 | ~n16732;
  assign n15930 = ~n15929 & ~n15928;
  assign n10792 = ~n10791 & ~n10790;
  assign n14789 = ~n16735 | ~n16424;
  assign n13120 = ~n13124 & ~n13679;
  assign n14854 = ~n16730 | ~n16734;
  assign n16718 = ~n14636 & ~n14770;
  assign n13895 = ~n16442 | ~n13894;
  assign n13816 = ~n13989 & ~n15323;
  assign n10608 = ~n10607 | ~n16721;
  assign n13763 = ~n13760 | ~n13759;
  assign n13910 = ~n13901 | ~n15596;
  assign n13934 = ~n13937 & ~n15653;
  assign n13127 = ~n13124 & ~n13123;
  assign n16727 = ~n16722 & ~n16721;
  assign n14414 = ~n15936 & ~n14413;
  assign n16055 = ~n16106 & ~n15910;
  assign n16294 = ~n15936 | ~n15933;
  assign n15905 = ~n15904 | ~n15903;
  assign n13703 = ~n13760 | ~n13226;
  assign n13892 = ~n16438 | ~n13894;
  assign n14727 = ~n10775 & ~n10774;
  assign n13631 = ~n13628 | ~n13627;
  assign n14743 = ~n14736 | ~n15428;
  assign n14631 = ~n16720 | ~n15342;
  assign n13876 = ~n13875 & ~n15240;
  assign n9715 = ~n10642 | ~n10641;
  assign n14244 = ~n14242 & ~n15534;
  assign n16194 = ~n14237 | ~n14235;
  assign n16712 = ~n16711 | ~n16710;
  assign n13739 = ~n13737 | ~n16438;
  assign n14202 = ~n14201 | ~n14200;
  assign n16726 = ~n16725 & ~n16724;
  assign n13736 = ~n13737 | ~n16442;
  assign n13760 = ~n13700 & ~n13699;
  assign n13804 = ~n13911 | ~n13802;
  assign n13711 = ~n13753 & ~n15653;
  assign n13670 = ~n16442 | ~n13669;
  assign n14434 = ~n10743 & ~n10742;
  assign n10770 = ~n14400 & ~n9770;
  assign n13667 = ~n16438 | ~n13669;
  assign n10258 = ~n10256 | ~n15596;
  assign n14309 = ~n14400 & ~n15536;
  assign n14412 = ~n14400 | ~n14243;
  assign n14242 = ~n14400 & ~n14243;
  assign n12978 = ~n12976 & ~n13679;
  assign n14773 = ~n16723 | ~n16721;
  assign n15927 = ~n14400 & ~n14611;
  assign n14660 = ~n16723 & ~n16433;
  assign n10614 = ~n12976 & ~n10218;
  assign n10782 = ~n12976 & ~n14967;
  assign n15898 = ~n15896 | ~n16228;
  assign n13981 = ~n13976 & ~n16423;
  assign n13658 = ~n13657 & ~n15240;
  assign n15912 = ~n16107 & ~n15907;
  assign n13614 = ~n13611 | ~n13610;
  assign n16715 = ~n16705 | ~n16704;
  assign n13563 = ~n15323 & ~n13562;
  assign n14374 = ~n14085 & ~n16660;
  assign n13588 = ~n13617 & ~n15653;
  assign n13801 = ~n13799 | ~n13798;
  assign n16687 = ~n16686 & ~n16685;
  assign n15915 = ~n14337;
  assign n10761 = ~n12785 & ~n14967;
  assign n14230 = ~n14337 & ~n14737;
  assign n16686 = ~n16690 & ~n16689;
  assign n14195 = ~n14337 & ~n14214;
  assign n16286 = ~n16058 | ~n16057;
  assign n13533 = ~n13525 & ~n15426;
  assign n15896 = ~n15895;
  assign n10596 = ~n12785 & ~n10218;
  assign n14515 = ~n16702 & ~n16433;
  assign n16714 = ~n16702 & ~n16703;
  assign n16708 = ~n16694 | ~n16693;
  assign n16707 = ~n16698 | ~n16697;
  assign n14337 = ~n10746 & ~n10745;
  assign n16101 = ~n14262 | ~n14610;
  assign n13877 = ~n13889 & ~n16423;
  assign n10571 = ~n14321 | ~n14492;
  assign n13863 = ~n13889 & ~n15455;
  assign n13914 = ~n13913 & ~n13912;
  assign n13867 = ~n13866 | ~n15557;
  assign n13559 = ~n13607 & ~n11663;
  assign n13889 = ~n13858 & ~n13857;
  assign n10554 = ~n14162 | ~n16680;
  assign n12652 = ~n12490;
  assign n14493 = ~n16695 | ~n14492;
  assign n14287 = ~n16675 & ~n16433;
  assign n10580 = ~n12490 & ~n10218;
  assign n14389 = ~n16695 & ~n16433;
  assign n10139 = ~n10124 | ~n15511;
  assign n14377 = ~n16675 & ~n16680;
  assign n15882 = ~n16230 & ~n16021;
  assign n10746 = ~n12490 & ~n14967;
  assign n14229 = ~n15902 & ~n14610;
  assign n14213 = ~n15902 & ~n14212;
  assign n14187 = ~n16230;
  assign n15908 = ~n15902 | ~n15901;
  assign n13644 = ~n13664 & ~n15455;
  assign n10460 = ~n15880 | ~n10901;
  assign n14178 = ~n15880;
  assign n13296 = ~n13295 | ~n13294;
  assign n10467 = ~n15880 | ~n10907;
  assign n16675 = ~n16679;
  assign n13568 = ~n13567 | ~n15863;
  assign n14361 = ~n16679 | ~n16680;
  assign n14376 = ~n16679 & ~n16676;
  assign n13295 = ~n13292 | ~n15511;
  assign n13513 = ~n13512 | ~n15511;
  assign n13651 = ~n13650 | ~n15557;
  assign n10734 = ~n12315 & ~n14967;
  assign n15256 = ~n15199 | ~n15198;
  assign n15377 = ~n15376 | ~n15375;
  assign n10562 = ~n12315 & ~n10218;
  assign n13912 = ~n13809 & ~n16228;
  assign n10451 = ~n12176 | ~n10842;
  assign n13547 = ~n13191 & ~n13548;
  assign n15199 = ~n15195 | ~n15194;
  assign n13444 = ~n13442 & ~n16431;
  assign n13511 = ~n10019 | ~n13289;
  assign n14273 = ~n16659 | ~n16665;
  assign n16654 = ~n16653 | ~n16652;
  assign n13243 = ~n13241 | ~n14669;
  assign n12176 = n10441 ^ ~n10440;
  assign n15373 = ~n15254 | ~n15253;
  assign n10405 = ~n14130;
  assign n13553 = ~n13552 & ~n15479;
  assign n13805 = ~n13686 | ~n16156;
  assign n10535 = ~n14041 | ~n16665;
  assign n15887 = ~n15888 | ~n13808;
  assign n15190 = ~n14701 | ~n14700;
  assign n10431 = ~n15888 & ~n9770;
  assign n14088 = ~n16658 & ~n16433;
  assign n10441 = ~n10439;
  assign n13552 = ~n13551 & ~n16185;
  assign n13927 = ~n15888 | ~n13817;
  assign n14372 = n16658 & n16665;
  assign n14282 = ~n16658 & ~n16665;
  assign n16880 = ~n16650 | ~n16651;
  assign n14275 = ~n16658 | ~n16669;
  assign n13189 = ~n13187 | ~n13186;
  assign n13802 = ~n15888 | ~n15885;
  assign n14130 = n10384 ^ n10904;
  assign n14059 = ~n15888;
  assign n13174 = ~n13170 & ~n16365;
  assign n10386 = ~n14135 | ~n10907;
  assign n14072 = ~n14071 | ~n14079;
  assign n15180 = ~n15179 | ~n15178;
  assign n10404 = ~n14108;
  assign n10400 = ~n14108 & ~n10403;
  assign n15254 = ~n15281 | ~n15251;
  assign n13200 = ~n13196 | ~n15637;
  assign n10383 = ~n13797 & ~n9770;
  assign n13798 = ~n13797 | ~n14116;
  assign n10422 = ~n11962 & ~n14967;
  assign n13550 = ~n13549 | ~n13548;
  assign n14696 = ~n14590 | ~n14589;
  assign n13087 = ~n13083 | ~n13082;
  assign n13926 = ~n13797 | ~n13704;
  assign n16626 = ~n16625 & ~n16624;
  assign n16627 = ~n16603 & ~n16602;
  assign n14076 = ~n14075 | ~n14074;
  assign n15209 = ~n15208 | ~n15207;
  assign n16636 = ~n16642 | ~n13960;
  assign n10505 = n10507 ^ n13960;
  assign n10399 = ~n14113 | ~n10907;
  assign n16060 = ~n14113 | ~n13694;
  assign n16634 = ~n16633 | ~n16632;
  assign n13065 = ~n13063 | ~n13062;
  assign n12968 = ~n12966 & ~n12965;
  assign n16642 = ~n16637;
  assign n13704 = n13619 & n13581;
  assign n10396 = ~n13619 & ~n9770;
  assign n16282 = ~n13619 | ~n14136;
  assign n16633 = ~n16630 | ~n16629;
  assign n13950 = ~n16637 | ~n13960;
  assign n14113 = ~n13619;
  assign n14585 = ~n14018 | ~n14017;
  assign n13719 = ~n13870 | ~n13730;
  assign n13887 = ~n13870 & ~n16433;
  assign n13545 = ~n16059;
  assign n14719 = ~P2_REG2_REG_15__SCAN_IN | ~n14718;
  assign n16617 = ~n16469 | ~n16468;
  assign n10254 = ~n10253 | ~n13730;
  assign n13595 = n10253 ^ n13730;
  assign n10301 = ~n15849 | ~n10907;
  assign n13720 = ~n16628 | ~n16631;
  assign n14577 = ~n14576 | ~n14575;
  assign n16620 = ~n16621 & ~n16465;
  assign n16183 = ~n16061 | ~n13190;
  assign n13604 = ~n15849;
  assign n10294 = ~n15849 | ~n10901;
  assign n14013 = ~n13781 | ~n13780;
  assign n10193 = ~n11714 & ~n15584;
  assign n12891 = ~n12890 | ~n15796;
  assign n10212 = ~n13346;
  assign n10211 = ~n13346 | ~n16466;
  assign n13541 = ~n15839 | ~n13202;
  assign n13061 = ~n16271;
  assign n10275 = ~n15835 | ~n10907;
  assign n13364 = ~n13648;
  assign n16615 = ~n16467 | ~n16466;
  assign n16621 = ~n16464 | ~n16463;
  assign n12746 = ~n12744 & ~n16173;
  assign n10272 = ~n15839 & ~n9770;
  assign n14028 = ~P2_REG1_REG_13__SCAN_IN | ~n14027;
  assign n16467 = ~n13635;
  assign n16604 = ~n13635 | ~n13634;
  assign n16271 = ~n15819 | ~n15829;
  assign n14601 = ~n14600 | ~n14599;
  assign n13776 = ~n13261 | ~n13260;
  assign n12744 = ~n12582 | ~n12581;
  assign n15781 = ~n15771 & ~n15770;
  assign n10225 = ~n11519 & ~n15584;
  assign n10049 = ~n13509;
  assign n13256 = ~n13044 | ~n13043;
  assign n13073 = ~n12898 | ~n12897;
  assign n16834 = ~n16925 | ~n16798;
  assign n13835 = ~n13834 | ~n13833;
  assign n13843 = ~n13842 | ~n13841;
  assign n15560 = ~n16809 & ~n15559;
  assign n12582 = ~n12580 | ~n12579;
  assign n14036 = ~P2_REG2_REG_13__SCAN_IN | ~n14035;
  assign n15447 = ~n16775 & ~n15559;
  assign n13768 = ~n13767 | ~n13766;
  assign n10056 = ~n10055 | ~n10054;
  assign n12365 = ~n12363 & ~n12362;
  assign n9646 = ~n9647;
  assign n13066 = ~n13089 | ~n13283;
  assign n12689 = ~n9685 & ~n12417;
  assign n15561 = ~n15575 & ~n16411;
  assign n15235 = ~n15575 & ~n15559;
  assign n10017 = ~n10016;
  assign n13376 = ~n16607 & ~n16608;
  assign n13143 = ~n13089 | ~n13088;
  assign n13839 = ~n13489 | ~n13488;
  assign n10046 = ~n13517 | ~n10907;
  assign n13832 = ~n13483 & ~n13482;
  assign n13402 = n13436 & n13401;
  assign n10057 = ~n10052 | ~n10053;
  assign n12888 = ~n16085;
  assign n10043 = ~n13517 | ~n10901;
  assign n13792 = ~n13791 | ~n13790;
  assign n13378 = ~n16610 & ~n16605;
  assign n16270 = ~n13517 | ~n13283;
  assign n16607 = ~n16610;
  assign n13362 = ~n16610 | ~n16608;
  assign n9991 = ~n9990 | ~n9989;
  assign n13270 = ~P2_REG1_REG_11__SCAN_IN | ~n13269;
  assign n16592 = ~n13409 | ~n13101;
  assign n16539 = ~n16530 | ~n16529;
  assign n12418 = ~n9684 & ~n12079;
  assign n16085 = ~n13293 | ~n15803;
  assign n16356 = ~n15579;
  assign n16425 = ~n16358 | ~n14429;
  assign n13407 = n9625 ^ n13101;
  assign n9626 = ~n9625 | ~n13101;
  assign n10029 = ~n11262 | ~n9810;
  assign n10011 = ~n15802 & ~n9770;
  assign n13480 = ~n12573 | ~n12572;
  assign n9609 = ~n9608;
  assign n9625 = n13230 ^ n15591;
  assign n13278 = ~P2_REG2_REG_11__SCAN_IN | ~n13277;
  assign n12373 = ~n12372 | ~n16256;
  assign n15413 = ~n15673 | ~n15533;
  assign n16586 = ~n13230 | ~n13325;
  assign n12080 = ~n9683 & ~n11903;
  assign n16759 = ~n10675 | ~n10674;
  assign n12372 = ~n12370 | ~n16168;
  assign n12747 = ~n15776 | ~n12597;
  assign n16514 = ~n16500 | ~n16499;
  assign n12424 = ~P2_STATE_REG_SCAN_IN | ~n14167;
  assign n15540 = ~n16018 | ~n15533;
  assign n12238 = ~n12236 | ~n12235;
  assign n13031 = ~n13030 | ~n13029;
  assign n13010 = ~n9583 & ~n12997;
  assign n9960 = ~n9959 | ~n9958;
  assign n10874 = ~n15520 | ~n10907;
  assign n10855 = ~n15969 | ~n10906;
  assign n9624 = ~n11163 & ~n15584;
  assign n10877 = ~n15520 | ~n10906;
  assign n10852 = ~n15969 | ~n10907;
  assign n15485 = ~n15999 | ~n15484;
  assign n15792 = ~n15788 | ~n15789;
  assign n12370 = ~n12367 | ~n16164;
  assign n10722 = ~n15999 | ~n10907;
  assign n16576 = ~n13315 | ~n13023;
  assign n12994 = ~n13016 | ~n12997;
  assign n15772 = ~n9949 | ~n9948;
  assign n12547 = ~n9561 | ~n9560;
  assign n16170 = ~n12587 | ~n16260;
  assign n12045 = ~n12043 & ~n16160;
  assign n16513 = ~n16512 & ~n16511;
  assign n11904 = ~n9682 & ~n11707;
  assign n16494 = ~n16491 | ~n16503;
  assign n12367 = ~n12050 | ~n16248;
  assign n13055 = ~n13054 | ~n13053;
  assign n12160 = ~n11611 | ~n11610;
  assign n16512 = ~n16505 & ~n16504;
  assign n14779 = ~n16724 | ~n16345;
  assign n9949 = ~n11070 | ~n10842;
  assign n13053 = ~n12539 | ~n12538;
  assign n11988 = ~n11987 | ~n11986;
  assign n9911 = ~n12439 | ~n9910;
  assign n15655 = n10888 & P1_REG3_REG_28__SCAN_IN;
  assign n12151 = ~n11599 & ~n11598;
  assign n12050 = ~n16064 | ~n16244;
  assign n11708 = ~n9681 & ~n11549;
  assign n15502 = ~n13226 | ~n15533;
  assign n12528 = ~n12101 | ~n12100;
  assign n11535 = ~n11534 | ~n11533;
  assign n15068 = ~n13226 & ~P1_REG2_REG_26__SCAN_IN;
  assign n11722 = ~n9802 | ~n9801;
  assign n14878 = ~n13226 & ~P1_REG2_REG_24__SCAN_IN;
  assign n16505 = ~n16487 | ~n16486;
  assign n10850 = ~n10849 | ~n10848;
  assign n9934 = ~n9933 | ~n9932;
  assign n9561 = ~n9558 | ~n13015;
  assign n9204 = ~n9587 | ~n9586;
  assign n15617 = ~n15596;
  assign n11814 = ~n11811 & ~n16159;
  assign n15754 = ~n15750;
  assign n9914 = n9907 ^ n11662;
  assign n9393 = ~n11886 & ~n11885;
  assign n15521 = ~n15094;
  assign n16381 = ~n16383;
  assign n9801 = ~n9800 | ~n9799;
  assign n16377 = ~n16378;
  assign n15324 = ~n15323 | ~n15322;
  assign n16487 = ~n16481 | ~n16480;
  assign n12810 = ~n16551;
  assign n16486 = ~n16485 | ~n16484;
  assign n9913 = ~n9909 & ~n9908;
  assign n15146 = ~n15604;
  assign n12459 = n9488 ^ n16522;
  assign n12187 = n9508 ^ n12467;
  assign n9653 = ~n9649 | ~n11891;
  assign n12762 = ~n12765;
  assign n16551 = ~n9548 | ~n9547;
  assign n14914 = ~n14611;
  assign n16501 = ~n16493 | ~n16492;
  assign n12235 = ~n16249 | ~n12366;
  assign n12098 = ~n12007 | ~n12006;
  assign n16235 = ~n11679 | ~n16237;
  assign n11811 = ~n11685 | ~n11684;
  assign n12322 = n9889 ^ n10904;
  assign n9889 = ~n9888 | ~n9887;
  assign n11532 = ~n11529 | ~n11528;
  assign n12765 = ~n9527 | ~n9526;
  assign n12400 = ~n16855;
  assign n11724 = ~n9796 | ~n9795;
  assign n10646 = ~n15591;
  assign n11679 = ~n15703 | ~n11925;
  assign n9924 = ~n11039 | ~n10842;
  assign n12124 = ~n12123 | ~n12122;
  assign n10553 = ~n14300 | ~n8930;
  assign n13634 = ~n16466;
  assign n12122 = ~n12023 | ~n12022;
  assign n15731 = ~n15738 | ~n12217;
  assign n11529 = ~n9383 | ~n9403;
  assign n12420 = ~n16471;
  assign n11526 = ~n11525 | ~n11891;
  assign n12675 = ~n12467;
  assign n11659 = ~n11658 | ~n11657;
  assign n9020 = ~n9019 | ~n10969;
  assign n14450 = ~n11196 | ~n13881;
  assign n11530 = ~n13871 | ~n16947;
  assign n13503 = ~n15803;
  assign n15777 = ~n15773;
  assign n13731 = ~n16431;
  assign n12004 = ~n11856 | ~n11855;
  assign n16475 = ~n9417 & ~n9416;
  assign n16608 = ~n9645 & ~n9644;
  assign n16466 = ~n9375 | ~n9374;
  assign n13859 = ~n10234 | ~n10233;
  assign n15883 = ~n14177;
  assign n12997 = ~n9582 | ~n9581;
  assign n10179 = ~n10178 | ~n10177;
  assign n13960 = ~n10199 & ~n10198;
  assign n13015 = ~n9557 | ~n9556;
  assign n10534 = ~n14101 | ~n8930;
  assign n12769 = ~n9535 | ~n9534;
  assign n15820 = ~n10068 | ~n10067;
  assign n10476 = ~n10475 & ~n10474;
  assign n12375 = ~n9904 | ~n9903;
  assign n15803 = ~n10009 & ~n10008;
  assign n14060 = ~n10381 | ~n10380;
  assign n15789 = ~n9981 | ~n9980;
  assign n14136 = ~n10312 | ~n10311;
  assign n15751 = ~n9931 | ~n9930;
  assign n15840 = ~n10158 & ~n10157;
  assign n15773 = ~n9956 | ~n9955;
  assign n11655 = ~n10113 | ~n10112;
  assign n10199 = ~n10195 | ~n10194;
  assign n11524 = ~n9405;
  assign n9603 = ~n9602 | ~n9601;
  assign n11997 = ~n11759 | ~n8925;
  assign n16516 = ~n16507;
  assign n10172 = ~n13977 | ~n8930;
  assign n9362 = ~n9361 | ~n9360;
  assign n9425 = ~n9424 | ~n9423;
  assign n16496 = ~n12255;
  assign n9645 = ~n9641 | ~n9640;
  assign n9656 = ~n11767 | ~n14685;
  assign n13871 = ~n11767;
  assign n9019 = ~n9015 | ~n10135;
  assign n9331 = ~n11984 | ~n9405;
  assign n9832 = n9827 & n9826;
  assign n15394 = ~n15268;
  assign n11812 = ~n12480;
  assign n10157 = ~n10156 | ~n10155;
  assign n10158 = ~n10148 | ~n10147;
  assign n16847 = ~n8922;
  assign n11528 = ~n9385 | ~n16939;
  assign n11853 = ~n11575 | ~n11574;
  assign n12019 = ~n11876 | ~n11875;
  assign n10209 = n10208 & n10207;
  assign n9791 = ~n9770 & ~n15684;
  assign n10458 = ~n10454 | ~n10453;
  assign n10112 = ~n10961;
  assign n16507 = ~n9462 | ~n9461;
  assign n11759 = ~n8922 & ~n16798;
  assign n10115 = ~n10961 & ~P1_D_REG_1__SCAN_IN;
  assign n11663 = ~n11949 | ~n8924;
  assign n9623 = ~n9622 | ~n9621;
  assign n9411 = ~n9407 | ~n9406;
  assign n9512 = ~n9180 | ~n9179;
  assign n9015 = ~n10133 | ~n11667;
  assign n11761 = ~n8922 & ~n11760;
  assign n10851 = ~n10846 | ~n10845;
  assign n10119 = ~n10961 & ~P1_D_REG_0__SCAN_IN;
  assign n10560 = ~n16401 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n10926 = ~n8923;
  assign n10180 = ~n10174 | ~n10173;
  assign n10524 = ~n16401 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n15268 = ~P2_U3893 | ~n16958;
  assign n15398 = n9101 & n9100;
  assign n10639 = ~n16401 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n10678 = ~n16401 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n10684 = ~n16401 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n10693 = ~n16401 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n10191 = ~n16401 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n10223 = ~n16401 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n11949 = ~n11911 & ~n11662;
  assign n10514 = ~n16401 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n10198 = ~n10197 | ~n10196;
  assign n10111 = ~n10110 | ~n10109;
  assign n9324 = ~n9325 & ~P2_D_REG_1__SCAN_IN;
  assign n10549 = ~n13434;
  assign n16845 = n8926 ^ ~n16591;
  assign n10372 = ~n10371 | ~n10370;
  assign n9841 = ~n11044 | ~n10842;
  assign n11751 = ~n8926 | ~n9384;
  assign n10000 = ~n9999 | ~n9998;
  assign n15639 = ~n15484;
  assign n10118 = ~n10117 & ~n10116;
  assign n14935 = ~n15533;
  assign n10110 = ~n10107 | ~P1_B_REG_SCAN_IN;
  assign n11101 = ~n9756 & ~n9755;
  assign n11833 = ~n16146 | ~n10130;
  assign n10420 = ~n10864 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n9463 = ~n14149 & ~n13999;
  assign n13779 = n10206 ^ n10205;
  assign n10865 = ~n10864 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n10268 = ~n10864 | ~P2_DATAO_REG_13__SCAN_IN;
  assign n9101 = ~n9021 | ~n13119;
  assign n15484 = n16146 & n11686;
  assign n10843 = ~n10864 | ~P2_DATAO_REG_25__SCAN_IN;
  assign n16333 = ~n16328;
  assign n9813 = ~n10864 | ~P2_DATAO_REG_2__SCAN_IN;
  assign n8926 = n16918;
  assign n9342 = ~n9340 & ~n10520;
  assign n8920 = n9781;
  assign n10745 = ~n14970 & ~n12491;
  assign n15369 = ~P2_REG1_REG_18__SCAN_IN | ~n15381;
  assign n10005 = ~n9756 & ~n14005;
  assign n14971 = ~n14970 & ~n14969;
  assign n10781 = ~n14970 & ~n12883;
  assign n10864 = ~n14970;
  assign n14892 = ~n14970 & ~n14891;
  assign n9023 = ~n9022 | ~n13454;
  assign n10719 = ~n14970 & ~n13674;
  assign n10899 = ~n14970 & ~n13882;
  assign n10814 = ~n14970 & ~n13125;
  assign n10206 = ~n10204 | ~P2_IR_REG_31__SCAN_IN;
  assign n9098 = ~n9088 | ~n14426;
  assign n13454 = ~n9322;
  assign n14967 = ~n9810;
  assign n9756 = ~n14156;
  assign n15281 = ~n15184;
  assign n10120 = ~n10135 | ~P1_STATE_REG_SCAN_IN;
  assign n10204 = ~n9632 | ~n9631;
  assign n15381 = n10541 ^ P2_IR_REG_18__SCAN_IN;
  assign n9088 = ~n16591 | ~n13119;
  assign n10216 = ~n10215;
  assign n10240 = ~n10239;
  assign n10188 = ~n10187;
  assign n10363 = ~n10362;
  assign n8921 = ~n10218;
  assign n9474 = ~n14426 | ~n9043;
  assign n9329 = ~n13303 | ~n9328;
  assign n9344 = ~n11319 | ~n15386;
  assign n14156 = n9745 ^ ~P1_IR_REG_30__SCAN_IN;
  assign n9632 = ~n9630 | ~P2_IR_REG_31__SCAN_IN;
  assign n9752 = ~n9750 | ~n9749;
  assign n15386 = ~n15388;
  assign n13303 = n9001 ^ ~P2_IR_REG_24__SCAN_IN;
  assign n14426 = ~n16958 | ~n8918;
  assign n8968 = ~n8962 | ~n8961;
  assign n8953 = ~n8952 | ~P1_IR_REG_31__SCAN_IN;
  assign n10135 = n8973 ^ ~P1_IR_REG_23__SCAN_IN;
  assign n9322 = n8992 ^ P2_IR_REG_25__SCAN_IN;
  assign n9750 = ~n9747 | ~P1_IR_REG_29__SCAN_IN;
  assign n9286 = ~n9691;
  assign n10576 = ~n10575;
  assign n9011 = ~n9009 & ~n9008;
  assign n9630 = ~n9619 | ~n9618;
  assign n9732 = ~n9731 | ~SI_26_;
  assign n8973 = ~n8972 & ~n10417;
  assign n8962 = ~n8960 | ~P1_IR_REG_26__SCAN_IN;
  assign n14598 = ~n14587;
  assign n13119 = n9004 ^ P2_IR_REG_23__SCAN_IN;
  assign n9328 = ~n9738;
  assign n14717 = ~n14698;
  assign n16433 = ~n16961 | ~n16939;
  assign n9459 = n9064 ^ ~SI_3_;
  assign n9259 = ~n9257 & ~n9256;
  assign n9269 = ~n9267 & ~n9266;
  assign n10327 = ~n10326 | ~SI_27_;
  assign n9747 = ~n9746 | ~P1_IR_REG_31__SCAN_IN;
  assign n9213 = ~n9210 | ~n9209;
  assign n9408 = n9053 ^ ~n9051;
  assign n8960 = ~n8959 | ~P1_IR_REG_31__SCAN_IN;
  assign n10676 = n9723 ^ SI_25_;
  assign n9014 = ~n9012 | ~P1_IR_REG_31__SCAN_IN;
  assign n9511 = n9183 ^ SI_6_;
  assign n10342 = ~n10341 | ~SI_30_;
  assign n9379 = ~n9356 | ~n9355;
  assign n9069 = ~n9068 | ~n9067;
  assign n9210 = ~n9208 & ~n9207;
  assign n10341 = ~n10340 | ~n10339;
  assign n8970 = ~n8969 & ~n10417;
  assign n9202 = ~n9201 | ~n9200;
  assign n16939 = n9081 ^ P2_IR_REG_21__SCAN_IN;
  assign n10336 = ~n10335 | ~n10334;
  assign n9969 = ~n9996 & ~n10417;
  assign n9079 = ~n9077 & ~n10520;
  assign n8959 = ~n8969 | ~n8958;
  assign n9617 = ~n9613 | ~n9612;
  assign n14351 = ~n13679;
  assign n9591 = ~n9613 & ~n10520;
  assign n14157 = ~n13309;
  assign n9052 = ~n9051;
  assign n9570 = ~n9569 & ~n10520;
  assign n9721 = ~n10345 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n9245 = n8919 & P1_DATAO_REG_14__SCAN_IN;
  assign n9068 = ~n8919 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n9235 = ~n10345 & ~n9234;
  assign n9208 = ~n8919 & ~n9205;
  assign n9254 = ~n10345 & ~n9253;
  assign n9226 = ~n8919 & ~n11267;
  assign n9201 = ~n8919 | ~P1_DATAO_REG_9__SCAN_IN;
  assign n9244 = ~n10345 & ~n10282;
  assign n14034 = ~n14015;
  assign n16322 = n9288 ^ P1_IR_REG_19__SCAN_IN;
  assign n9182 = ~n8919 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n10032 = ~n10002 | ~P1_REG3_REG_9__SCAN_IN;
  assign n9192 = ~n8919 & ~n11054;
  assign n9706 = ~n10345 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n9279 = ~n8919 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n10247 = ~n9333 & ~P2_IR_REG_14__SCAN_IN;
  assign n9187 = ~n8919 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n9711 = ~n10345 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n9186 = ~n9043 | ~P2_DATAO_REG_7__SCAN_IN;
  assign n9274 = ~n10344 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n9181 = ~n9043 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n9044 = ~n9043 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n9058 = ~n9043 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n9200 = ~n10344 | ~P2_DATAO_REG_9__SCAN_IN;
  assign n9916 = ~n9943 & ~n10417;
  assign n9207 = ~n9043 & ~n9206;
  assign n9191 = ~n9043 & ~n9568;
  assign n9722 = ~n10344 | ~P2_DATAO_REG_25__SCAN_IN;
  assign n9216 = ~n10344 & ~n9635;
  assign n9517 = ~n9520 | ~P2_IR_REG_31__SCAN_IN;
  assign n10265 = ~n8944 | ~n9859;
  assign n9139 = ~n9138 & ~n10520;
  assign n9494 = ~n9516 & ~n10520;
  assign n10219 = ~n8982 | ~n8981;
  assign n8981 = ~n8980 & ~n9589;
  assign n9030 = ~n9029 & ~n9028;
  assign n9138 = ~n9493 & ~P2_IR_REG_3__SCAN_IN;
  assign n9516 = ~n9493 & ~n9492;
  assign n8997 = ~n8995 & ~P2_IR_REG_21__SCAN_IN;
  assign n9134 = ~n9493 | ~P2_IR_REG_31__SCAN_IN;
  assign n9096 = ~n9107 & ~n10520;
  assign n8965 = ~n8964 | ~n8963;
  assign n8986 = ~n8985 | ~n9341;
  assign n8987 = ~n8984 | ~n8983;
  assign n8949 = ~n8946 | ~n8945;
  assign n9518 = ~n9521 | ~P2_IR_REG_31__SCAN_IN;
  assign n8943 = ~n9833 | ~n8942;
  assign n9026 = ~n9025 | ~n9662;
  assign n8974 = ~P2_IR_REG_2__SCAN_IN;
  assign n9543 = ~P2_IR_REG_7__SCAN_IN;
  assign n8996 = ~P2_IR_REG_24__SCAN_IN & ~P2_IR_REG_22__SCAN_IN;
  assign n9491 = ~P2_IR_REG_4__SCAN_IN & ~P2_IR_REG_3__SCAN_IN;
  assign n9038 = ~SI_0_ | ~P2_DATAO_REG_0__SCAN_IN;
  assign n9046 = ~SI_0_ | ~P1_DATAO_REG_0__SCAN_IN;
  assign n9334 = ~P2_IR_REG_15__SCAN_IN;
  assign n9335 = ~P2_IR_REG_16__SCAN_IN;
  assign n9341 = ~P2_IR_REG_20__SCAN_IN;
  assign n9107 = ~P2_IR_REG_1__SCAN_IN & ~P2_IR_REG_0__SCAN_IN;
  assign n8975 = ~P2_IR_REG_9__SCAN_IN & ~P2_IR_REG_10__SCAN_IN;
  assign n8963 = ~P1_IR_REG_26__SCAN_IN;
  assign n9743 = ~P1_IR_REG_28__SCAN_IN;
  assign n8979 = ~P2_IR_REG_8__SCAN_IN;
  assign n9748 = ~P1_IR_REG_29__SCAN_IN;
  assign n9729 = ~SI_26_;
  assign n10364 = ~n9262 | ~n9261;
  assign n16134 = ~n14893 & ~n14892;
  assign n16900 = ~n16397 & ~n15590;
  assign n13431 = ~n9359 & ~n13999;
  assign n8922 = n16940;
  assign n16940 = n9342 ^ ~n9341;
  assign n9405 = ~n9330 | ~n9329;
  assign n11100 = ~n10714;
  assign n8923 = n11101;
  assign n16918 = n9343 ^ P2_IR_REG_19__SCAN_IN;
  assign n16774 = ~n16961 & ~n16939;
  assign n16044 = ~n16042 & ~n16041;
  assign n8929 = ~n9463;
  assign n8930 = ~n8929;
  assign n10730 = ~n11686 & ~n14900;
  assign n16958 = n9083 ^ P2_IR_REG_28__SCAN_IN;
  assign n10826 = ~n9957;
  assign n9428 = n15591 ^ n16476;
  assign n9446 = n15591 ^ n12255;
  assign n15591 = ~n9405 & ~n9404;
  assign n9037 = ~n9031 & ~n9030;
  assign n9726 = ~n9199;
  assign n9199 = ~n9037;
  assign n15087 = ~n10799 | ~n14907;
  assign n13103 = ~n13102 & ~n16584;
  assign n10795 = ~n10780 & ~n14729;
  assign n10777 = ~n14724 & ~n14727;
  assign n13346 = n13635 ^ n15591;
  assign n9367 = ~P2_REG3_REG_12__SCAN_IN;
  assign n9368 = ~n9380;
  assign n9355 = ~P2_REG3_REG_10__SCAN_IN;
  assign n16533 = ~n16525 | ~n16524;
  assign n16661 = ~n16683 | ~n16659;
  assign n11773 = ~n11772;
  assign n10015 = ~n9994 & ~n9993;
  assign n9993 = ~n9992;
  assign n9964 = n9960 ^ ~n11662;
  assign n9959 = ~n15772 | ~n10901;
  assign n11683 = ~n11928;
  assign n9263 = ~P2_DATAO_REG_16__SCAN_IN;
  assign n9206 = ~P1_DATAO_REG_10__SCAN_IN;
  assign n14074 = ~n14079;
  assign n10517 = n14075 ^ ~n15591;
  assign n10589 = n16702 ^ ~n15591;
  assign n9509 = ~n9508 | ~n12467;
  assign n9361 = ~n8930 | ~n13419;
  assign n11556 = ~n11555 | ~n11570;
  assign n12020 = ~n12012;
  assign n10667 = P2_REG3_REG_24__SCAN_IN | n10627;
  assign n10627 = n10647 | P2_REG3_REG_23__SCAN_IN;
  assign n13322 = ~n13409 | ~n13325;
  assign n10222 = ~n10558 | ~n14015;
  assign n9492 = ~n9491;
  assign n10433 = ~n13808 | ~n10906;
  assign n10833 = ~n15159;
  assign n9872 = ~n9871 | ~n9870;
  assign n12872 = ~n9962 | ~n9961;
  assign n10276 = n10273 ^ ~n11662;
  assign n10274 = ~n15836 | ~n10906;
  assign n10796 = n10792 ^ ~n11662;
  assign n10907 = ~n10826;
  assign n14237 = ~n15910;
  assign n13067 = ~n13517 | ~n13076;
  assign n10800 = ~n10864 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n9220 = ~n9219;
  assign n9478 = n9069 ^ SI_4_;
  assign n9641 = ~n8930 | ~n13395;
  assign n14041 = n16658 ^ ~n15591;
  assign n9354 = ~P2_REG3_REG_8__SCAN_IN;
  assign n10572 = ~n14321;
  assign n9371 = ~n8930 | ~n13356;
  assign n10208 = ~n13779 | ~n10558;
  assign n9366 = ~n9379;
  assign n13389 = n13331 ^ n16870;
  assign n13233 = n16868 ^ ~n13330;
  assign n9521 = ~P2_IR_REG_6__SCAN_IN;
  assign n10742 = ~n10741;
  assign n10743 = ~n10740;
  assign n15998 = ~n15999;
  assign n9998 = ~n10730 | ~n11507;
  assign n15132 = n10446 ^ n10445;
  assign n16485 = ~n16488 | ~n16482;
  assign n16503 = ~n16490 | ~n16489;
  assign n16614 = ~n16604;
  assign n15944 = ~n15943;
  assign n16232 = ~n16157 | ~n16156;
  assign n16795 = ~n16808 | ~n16798;
  assign n9536 = ~n12671 | ~n12769;
  assign n9431 = ~P1_DATAO_REG_2__SCAN_IN;
  assign n10016 = n10012 ^ ~n11662;
  assign n10045 = ~n13076 | ~n10906;
  assign n9246 = ~SI_14_;
  assign n10661 = ~n10660;
  assign n10658 = ~n15333;
  assign n10686 = n15576 ^ ~n15591;
  assign n10253 = n16628 ^ ~n15591;
  assign n16917 = ~n16939;
  assign n9485 = ~n8930 | ~n12659;
  assign n9094 = ~n9107 | ~P2_REG1_REG_0__SCAN_IN;
  assign n9146 = ~n11002 | ~P2_REG2_REG_2__SCAN_IN;
  assign n9147 = ~n9145 | ~n9144;
  assign n12014 = ~n12013 | ~n12012;
  assign n12123 = P2_REG2_REG_8__SCAN_IN ^ ~n12110;
  assign n13470 = ~P2_REG3_REG_13__SCAN_IN;
  assign n10647 = P2_REG3_REG_22__SCAN_IN | n10617;
  assign n10617 = n10598 | P2_REG3_REG_21__SCAN_IN;
  assign n9450 = ~n11418;
  assign n16347 = ~n16801 | ~n16346;
  assign n14846 = n16895 ^ n14990;
  assign n16884 = n16679 ^ n16680;
  assign n9622 = ~n16401 | ~P1_DATAO_REG_10__SCAN_IN;
  assign n16863 = n13016 ^ ~n12990;
  assign n16859 = ~n16553 | ~n16548;
  assign n9939 = ~n9938;
  assign n10882 = ~n10879;
  assign n10298 = n10295 ^ n10904;
  assign n10293 = ~n15850 | ~n10907;
  assign n10740 = n10737 ^ n10904;
  assign n10738 = ~n15901 | ~n10906;
  assign n10725 = ~n15999 | ~n10906;
  assign n10775 = n10757 ^ n10904;
  assign n10758 = ~n15916 | ~n10906;
  assign n10779 = n10771 ^ n10904;
  assign n10772 = ~n14611 | ~n10906;
  assign n10077 = n10071 ^ n11662;
  assign n10069 = ~n15820 | ~n10907;
  assign n12217 = ~n15739;
  assign n10834 = n10811 ^ ~n11662;
  assign n10809 = ~n15964 | ~n10907;
  assign n9988 = n9984 ^ ~n11662;
  assign n9982 = ~n15789 | ~n10907;
  assign n9986 = ~n15788 | ~n10907;
  assign n13509 = n10044 ^ n11662;
  assign n10042 = ~n13076 | ~n10907;
  assign n9874 = ~n9873 | ~n9872;
  assign n14108 = n10397 ^ ~n11662;
  assign n10454 = ~n8920 | ~n13819;
  assign n10453 = ~n8928 | ~P1_REG1_REG_18__SCAN_IN;
  assign n10147 = ~n8928 | ~P1_REG1_REG_13__SCAN_IN;
  assign n10148 = ~n11100 | ~P1_REG2_REG_13__SCAN_IN;
  assign n10156 = ~n8920 | ~n13520;
  assign n11486 = ~n11485 | ~n11484;
  assign n15535 = n15670 ^ n15496;
  assign n15311 = ~n15307 & ~n15306;
  assign n14928 = ~n14926 & ~n14925;
  assign n14405 = n16198 ^ n14548;
  assign n13152 = ~n13150 | ~n15637;
  assign n11684 = ~n15687;
  assign n10440 = n9281 ^ SI_18_;
  assign n10416 = ~n10368 | ~n10367;
  assign n9266 = ~SI_16_;
  assign n9256 = ~SI_15_;
  assign n10387 = ~P1_IR_REG_14__SCAN_IN;
  assign n9237 = ~SI_13_;
  assign n9211 = ~n9210;
  assign n9193 = ~SI_8_;
  assign n9860 = ~P1_IR_REG_4__SCAN_IN;
  assign n9056 = ~SI_2_;
  assign n12990 = ~n12997;
  assign n16462 = ~n13859;
  assign n15328 = n15330 ^ n15214;
  assign n9640 = ~n13431 | ~P2_REG1_REG_11__SCAN_IN;
  assign n9601 = ~n13430 | ~P2_REG0_REG_9__SCAN_IN;
  assign n10598 = P2_REG3_REG_20__SCAN_IN | n10581;
  assign n14622 = n16723 ^ ~n15591;
  assign n10518 = ~n10517;
  assign n16669 = ~n16665;
  assign n15333 = n15343 ^ n15591;
  assign n15329 = n16453 ^ n10646;
  assign n10590 = ~n10589;
  assign n16676 = ~n16680;
  assign n9353 = ~P2_REG3_REG_6__SCAN_IN;
  assign n10681 = ~n10680;
  assign n15352 = n10686 ^ n15572;
  assign n10586 = ~n10583 | ~n10582;
  assign n10550 = ~n10549 & ~n14296;
  assign n10169 = ~n10549 & ~n13973;
  assign n10197 = ~n13430 | ~P2_REG0_REG_15__SCAN_IN;
  assign n10174 = ~n13430 | ~P2_REG0_REG_14__SCAN_IN;
  assign n10229 = ~n13431 | ~P2_REG1_REG_13__SCAN_IN;
  assign n9370 = ~n13431 | ~P2_REG1_REG_12__SCAN_IN;
  assign n9363 = ~n9351 | ~n9350;
  assign n9440 = ~n13431 | ~P2_REG1_REG_2__SCAN_IN;
  assign n13430 = ~n10631;
  assign n9145 = n9157 ^ ~P2_REG2_REG_2__SCAN_IN;
  assign n9155 = ~n9119 | ~n9118;
  assign n9130 = n9157 ^ ~P2_REG1_REG_2__SCAN_IN;
  assign n11580 = n11570 ^ ~P2_REG2_REG_4__SCAN_IN;
  assign n11552 = n11554 ^ ~n11570;
  assign n11567 = n11570 ^ P2_REG1_REG_4__SCAN_IN;
  assign n11626 = n11628 ^ ~n11573;
  assign n11636 = n11628 ^ ~n11586;
  assign n11562 = ~n11561 | ~n11628;
  assign n12005 = n12012 ^ ~n12004;
  assign n12021 = n12012 ^ ~n12019;
  assign n12099 = P2_REG1_REG_8__SCAN_IN ^ ~n12110;
  assign n13793 = ~P2_REG2_REG_12__SCAN_IN | ~n13789;
  assign n14602 = ~P2_REG2_REG_14__SCAN_IN | ~n14598;
  assign n15267 = ~n15269 | ~P2_U3893;
  assign n16357 = P2_REG3_REG_28__SCAN_IN ^ ~n13400;
  assign n15239 = n10667 ^ n10666;
  assign n15341 = P2_REG3_REG_24__SCAN_IN ^ ~n10627;
  assign n15218 = P2_REG3_REG_23__SCAN_IN ^ ~n10647;
  assign n14808 = P2_REG3_REG_22__SCAN_IN ^ ~n10617;
  assign n14507 = P2_REG3_REG_20__SCAN_IN ^ ~n10581;
  assign n14381 = P2_REG3_REG_19__SCAN_IN ^ n10563;
  assign n14300 = P2_REG3_REG_18__SCAN_IN ^ ~n10546;
  assign n13746 = n10184 ^ P2_REG3_REG_15__SCAN_IN;
  assign n13356 = ~n10226 | ~n9369;
  assign n13367 = ~n13636;
  assign n14659 = n16890 ^ n14785;
  assign n14644 = ~n14643 | ~n14642;
  assign n14514 = ~n14506;
  assign n14388 = n16886 ^ n14494;
  assign n10559 = ~n10558 | ~n8926;
  assign n10526 = ~n11962 & ~n15584;
  assign n10523 = ~n10558 | ~n15184;
  assign n10513 = ~n10558 | ~n15192;
  assign n10190 = ~n10558 | ~n14698;
  assign n12939 = n16863 ^ ~n12984;
  assign n12830 = ~n12777 | ~n12776;
  assign n9497 = ~n9496 | ~n9495;
  assign n9480 = ~n9476 | ~n9475;
  assign n16476 = ~n9411 & ~n9410;
  assign n9522 = ~n9520;
  assign n10909 = ~n15673 | ~n10906;
  assign n12873 = ~n12871 | ~n12870;
  assign n14726 = ~n14724;
  assign n15885 = ~n13808;
  assign n15160 = ~n10834;
  assign n10812 = ~n15964 | ~n10906;
  assign n10797 = ~n10796;
  assign n14125 = ~n10403;
  assign n10786 = ~n8923 | ~P1_REG0_REG_22__SCAN_IN;
  assign n10783 = ~n8928 | ~P1_REG1_REG_22__SCAN_IN;
  assign n10765 = ~n8923 | ~P1_REG0_REG_21__SCAN_IN;
  assign n10762 = ~n8928 | ~P1_REG1_REG_21__SCAN_IN;
  assign n10427 = ~n8920 | ~n14058;
  assign n10040 = ~n10039 | ~n10038;
  assign n10041 = ~n10031 | ~n10030;
  assign n9852 = ~n8928 | ~P1_REG1_REG_4__SCAN_IN;
  assign n9807 = ~n8920 | ~P1_REG3_REG_2__SCAN_IN;
  assign n9754 = ~n8920 | ~P1_REG3_REG_0__SCAN_IN;
  assign n13834 = ~n13840 | ~n13832;
  assign n13842 = ~n13840 | ~n13839;
  assign n14760 = ~n15123 | ~n8934;
  assign n15517 = n10886 ^ n10887;
  assign n10419 = ~n10730 | ~n14755;
  assign n13617 = ~n13580;
  assign n10267 = ~n10730 | ~n12571;
  assign n13213 = ~n10375 | ~n10154;
  assign n13241 = n16181 ^ ~n13187;
  assign n9923 = ~n9922 & ~n9921;
  assign n15649 = ~n16366 & ~n11663;
  assign n14550 = n16200 ^ ~n14822;
  assign n14190 = n16194 ^ ~n14236;
  assign n14260 = n16192 ^ n14228;
  assign n13937 = n13912 ^ n13911;
  assign n13753 = n13805 ^ ~n13799;
  assign n13756 = ~n13754 | ~n16367;
  assign n12636 = ~n12595 | ~n12594;
  assign n12694 = ~n12379 & ~n12378;
  assign n12696 = n16170 ^ ~n12580;
  assign n9691 = n9693 ^ SI_19_;
  assign n9222 = ~n9629;
  assign n9228 = ~SI_12_;
  assign n9995 = ~P1_IR_REG_9__SCAN_IN;
  assign n10020 = ~P1_IR_REG_10__SCAN_IN;
  assign n9563 = ~n9565 & ~n9564;
  assign n10344 = ~n9037;
  assign n10705 = ~n10704 | ~n10703;
  assign n10503 = ~n15604 | ~n15589;
  assign n13026 = ~n9578 | ~n9598;
  assign n13349 = n13348 ^ ~n13347;
  assign n13977 = P2_REG3_REG_16__SCAN_IN ^ ~n10488;
  assign n13469 = n13468 ^ ~n13467;
  assign n9659 = ~n9654 | ~n15596;
  assign n9654 = n10201 ^ ~n9648;
  assign n15354 = n15353 ^ ~n15352;
  assign n15360 = ~n15359 | ~n15358;
  assign n16605 = ~n16608;
  assign n13410 = ~n13023;
  assign n14035 = n14034 ^ n14033;
  assign n14032 = ~n14025 | ~n14024;
  assign n14718 = n14717 ^ n14716;
  assign n14579 = P2_REG1_REG_15__SCAN_IN ^ n14710;
  assign n14596 = ~n14595 | ~n14594;
  assign n14594 = ~n14593 | ~n15394;
  assign n14713 = n15178 ^ n15179;
  assign n14715 = ~n14708 | ~n14707;
  assign n15252 = n15281 ^ n15251;
  assign n15183 = P2_REG1_REG_17__SCAN_IN ^ n15282;
  assign n14654 = ~n16720 | ~n16424;
  assign n14509 = ~n14649 | ~n16424;
  assign n13743 = ~n13740 | ~n16419;
  assign n13395 = ~n9381 | ~n9380;
  assign n13336 = ~n13335 | ~n13334;
  assign n13335 = ~n13389 | ~n13731;
  assign n13234 = ~n13233 | ~n13731;
  assign n14352 = ~n14968;
  assign n9737 = ~n13459;
  assign n14439 = P1_REG3_REG_19__SCAN_IN ^ n10711;
  assign n10936 = ~n15495 | ~n15516;
  assign n13525 = n13524 ^ ~n13523;
  assign n13523 = ~n13522 | ~n13521;
  assign n13819 = P1_REG3_REG_18__SCAN_IN ^ ~n10470;
  assign n10469 = n10468 ^ ~n10726;
  assign n15136 = n15135 ^ ~P1_REG2_REG_19__SCAN_IN;
  assign n15127 = n8924 ^ ~n15126;
  assign n14307 = n16196 ^ n14399;
  assign n14252 = ~n14736 | ~n15660;
  assign n14268 = ~n14261 | ~n15659;
  assign n13984 = n14185 ^ ~n14180;
  assign n13217 = ~n13216 | ~n13215;
  assign n13215 = ~n13214 | ~n14547;
  assign n13156 = ~n13155 | ~n13176;
  assign n10637 = ~n10636;
  assign n16504 = ~n16503 | ~n16502;
  assign n16502 = ~n16501;
  assign n16558 = ~n16557 | ~n16556;
  assign n16556 = ~n16560 | ~n16555;
  assign n16568 = ~n16567 | ~n16566;
  assign n16571 = ~n16570;
  assign n16589 = ~n16588 | ~n16587;
  assign n16587 = ~n16586 | ~n16585;
  assign n15782 = ~n15781 & ~n15780;
  assign n16619 = ~n16618 | ~n16617;
  assign n16616 = ~n16614 & ~n16613;
  assign n16459 = ~n16458 & ~n16774;
  assign n16460 = ~n16457 & ~n16798;
  assign n16457 = ~n16456;
  assign n16640 = ~n16639 | ~n16638;
  assign n16648 = ~n16647 | ~n16646;
  assign n16647 = ~n16644 | ~n16643;
  assign n15833 = ~n15832 & ~n16021;
  assign n15855 = ~n15838 & ~n15837;
  assign n16668 = ~n16667 | ~n16666;
  assign n16662 = ~n16661 | ~n16660;
  assign n15867 = ~n15866 | ~n15865;
  assign n16711 = ~n16715 | ~n16706;
  assign n16709 = ~n16707;
  assign n16700 = ~n16699 | ~n16707;
  assign n15893 = ~n15892 | ~n15891;
  assign n15904 = ~n15900 | ~n15899;
  assign n15900 = ~n15898 | ~n15897;
  assign n16737 = ~n16741;
  assign n15921 = ~n15920 & ~n15919;
  assign n15923 = ~n16106 & ~n16021;
  assign n15946 = ~n15945 | ~n15944;
  assign n16757 = ~n16756 | ~n16755;
  assign n16763 = ~n16762 & ~n16761;
  assign n15991 = ~n15990 | ~n15989;
  assign n15679 = ~n16227 | ~n15677;
  assign n16190 = ~n16189 | ~n16188;
  assign n16189 = ~n16286;
  assign n16116 = ~n16114 & ~n16113;
  assign n16111 = ~n16110 | ~n16109;
  assign n16110 = ~n16108 | ~n16107;
  assign n16796 = ~n16806;
  assign n16891 = ~n16890 | ~n16889;
  assign n16889 = ~n16888 & ~n16887;
  assign n16887 = ~n16886 | ~n16885;
  assign n16020 = ~n16017;
  assign n16019 = ~n16018 | ~n16370;
  assign n16013 = ~n16017 | ~n16012;
  assign n16014 = ~n16008 | ~n16007;
  assign n16058 = ~n16229;
  assign n16252 = ~n15731 | ~n12366;
  assign n16817 = ~n16801;
  assign n16821 = ~n16913 | ~n16591;
  assign n14637 = ~n16706;
  assign n16303 = ~n16300 & ~n16299;
  assign n16300 = ~n16298 & ~n16297;
  assign n16129 = ~n16226 | ~n16126;
  assign n16126 = ~n16227 | ~n16125;
  assign n16125 = ~n16124 & ~n16299;
  assign n16135 = ~n16134 & ~n16133;
  assign n16109 = ~n15927;
  assign n16164 = ~n16252;
  assign n16168 = ~n16259 & ~n12369;
  assign n16256 = ~n16166;
  assign n16073 = ~n15754 & ~n15751;
  assign n9205 = ~P2_DATAO_REG_10__SCAN_IN;
  assign n9583 = n13016 ^ n15591;
  assign n9605 = n13315 ^ n15591;
  assign n16825 = ~n16906 | ~n16591;
  assign n16824 = ~n16913 | ~n16798;
  assign n16925 = ~n16933;
  assign n13257 = ~n13046 | ~n13045;
  assign n14014 = ~n13783 | ~n13782;
  assign n16630 = ~n16458;
  assign n16924 = ~n16409 & ~n16408;
  assign n16913 = ~n16905;
  assign n14992 = ~n16747;
  assign n16731 = ~n16734;
  assign n16666 = ~n16650;
  assign n16660 = ~n16651;
  assign n9635 = ~P1_DATAO_REG_11__SCAN_IN;
  assign n16584 = ~n16573;
  assign n9937 = n9934 ^ n11662;
  assign n9933 = ~n15750 | ~n10901;
  assign n9932 = ~n15751 | ~n9957;
  assign n9798 = ~n11378;
  assign n16307 = ~n16226;
  assign n16154 = n16314 ^ n16313;
  assign n14924 = ~n16121;
  assign n16113 = ~n16294;
  assign n10732 = ~n10864 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n13690 = ~n16187;
  assign n16260 = ~n16073;
  assign n16248 = ~n16063;
  assign n16249 = ~n16067;
  assign n10330 = ~n10344 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n10329 = ~n8919 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n10325 = ~n10344 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n9253 = ~P2_DATAO_REG_15__SCAN_IN;
  assign n9234 = ~P2_DATAO_REG_13__SCAN_IN;
  assign n9209 = ~SI_10_;
  assign n9568 = ~P1_DATAO_REG_8__SCAN_IN;
  assign n9029 = ~n9027 | ~P1_ADDR_REG_19__SCAN_IN;
  assign n9060 = ~n9437;
  assign n13013 = ~n12550 & ~n9562;
  assign n9488 = n15591 ^ n16523;
  assign n9508 = n15591 ^ n12407;
  assign n10623 = n16730 ^ ~n15591;
  assign n9647 = n16610 ^ n15591;
  assign n12671 = n12765 ^ n15591;
  assign n10680 = n16760 ^ ~n15591;
  assign n10194 = ~n13434 | ~P2_REG2_REG_15__SCAN_IN;
  assign n10196 = ~n13431 | ~P2_REG1_REG_15__SCAN_IN;
  assign n10177 = ~n13434 | ~P2_REG2_REG_14__SCAN_IN;
  assign n10173 = ~n13431 | ~P2_REG1_REG_14__SCAN_IN;
  assign n9360 = ~n13430 | ~P2_REG0_REG_10__SCAN_IN;
  assign n9156 = ~n9121 | ~n9120;
  assign n11419 = n9148 ^ n9450;
  assign n9167 = ~n9165 | ~n9450;
  assign n11629 = n11560 ^ n11585;
  assign n11854 = P2_REG1_REG_6__SCAN_IN ^ n11872;
  assign n11863 = ~n11862 | ~n11861;
  assign n12009 = n12011 ^ n12020;
  assign n12107 = n12109 ^ n12121;
  assign n12515 = n12517 ^ n12536;
  assign n13038 = n13040 ^ n13052;
  assign n13255 = n13257 ^ ~n13258;
  assign n13775 = n13779 ^ ~n13777;
  assign n13032 = ~P2_REG1_REG_10__SCAN_IN | ~n13052;
  assign n14012 = n14014 ^ n14034;
  assign n14584 = n14586 ^ n14598;
  assign n14695 = n14697 ^ n14717;
  assign n14578 = ~P2_REG1_REG_14__SCAN_IN | ~n14598;
  assign n15189 = n15191 ^ ~n15192;
  assign n15198 = n15257 ^ n15281;
  assign n15265 = ~n15256;
  assign n15181 = ~P2_REG1_REG_16__SCAN_IN | ~n15206;
  assign n15565 = P2_REG3_REG_27__SCAN_IN ^ ~n10697;
  assign n10498 = n10667 | P2_REG3_REG_25__SCAN_IN;
  assign n10207 = ~n16401 | ~P1_DATAO_REG_12__SCAN_IN;
  assign n12392 = ~n16542;
  assign n12391 = ~n16540;
  assign n11760 = ~n16798 | ~n16917;
  assign n9382 = ~n16847 | ~n16939;
  assign n16412 = ~n16346 | ~n14427;
  assign n15574 = ~n15454 & ~n15453;
  assign n15445 = n16894 ^ n15551;
  assign n14994 = ~n16753;
  assign n15003 = ~n14856 & ~n14855;
  assign n14855 = ~n14854;
  assign n14640 = n16890 ^ ~n14772;
  assign n14506 = n16888 ^ n14648;
  assign n14491 = n16888 ^ n14638;
  assign n16886 = n16695 ^ ~n16696;
  assign n14365 = n16886 ^ ~n14488;
  assign n14277 = n16884 ^ ~n14362;
  assign n14078 = n16882 ^ ~n14274;
  assign n13954 = n16880 ^ n14070;
  assign n16878 = n16637 ^ n16645;
  assign n13722 = n16878 ^ n13951;
  assign n9476 = ~n16401 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n9388 = ~n11529;
  assign n11527 = ~n9321 & ~n9325;
  assign n9327 = ~n9325;
  assign n9326 = ~P2_D_REG_0__SCAN_IN;
  assign n8994 = ~P2_IR_REG_25__SCAN_IN;
  assign n8993 = ~P2_IR_REG_23__SCAN_IN;
  assign n8989 = ~P2_IR_REG_24__SCAN_IN;
  assign n9515 = ~P2_IR_REG_5__SCAN_IN;
  assign n12839 = ~n9915 & ~n12440;
  assign n9915 = ~n9912 & ~n9911;
  assign n10903 = ~n15673 | ~n10907;
  assign n10436 = n10432 ^ n10904;
  assign n9965 = ~n9964;
  assign n9966 = ~n9963;
  assign n10464 = n10461 ^ n11662;
  assign n10459 = ~n15883 | ~n10907;
  assign n11480 = ~n11246 | ~n11206;
  assign n11485 = ~n11241 | ~n11191;
  assign n11481 = ~n11480 | ~n11479;
  assign n11280 = ~P1_REG3_REG_8__SCAN_IN;
  assign n11305 = n11507 ^ P1_REG1_REG_10__SCAN_IN;
  assign n10149 = ~P1_REG3_REG_12__SCAN_IN;
  assign n13484 = n13490 ^ ~n13832;
  assign n13491 = n13490 ^ ~n13839;
  assign n14899 = ~n15496;
  assign n15298 = ~n15071;
  assign n14944 = ~n14898;
  assign n10848 = ~n8923 | ~P1_REG0_REG_25__SCAN_IN;
  assign n10845 = ~n8928 | ~P1_REG1_REG_25__SCAN_IN;
  assign n14413 = ~n14412;
  assign n14556 = ~n14555;
  assign n10371 = ~n10864 | ~P2_DATAO_REG_16__SCAN_IN;
  assign n10392 = ~n10864 | ~P2_DATAO_REG_15__SCAN_IN;
  assign n11308 = ~P1_REG3_REG_10__SCAN_IN;
  assign n9896 = ~n9895 | ~n9894;
  assign n12596 = ~n12224 | ~n12371;
  assign n12348 = ~n12041 | ~n12040;
  assign n15309 = ~n15429;
  assign n14825 = n16202 ^ ~n14930;
  assign n14207 = n16192 ^ n14206;
  assign n13810 = n14185 ^ n14186;
  assign n13693 = n13805 ^ ~n13806;
  assign n13580 = n16187 ^ n13687;
  assign n13570 = n16187 ^ n13691;
  assign n13196 = n16183 ^ ~n13549;
  assign n13082 = ~n13081 | ~n13080;
  assign n13088 = ~n13141;
  assign n13141 = ~n15802 | ~n12907;
  assign n9999 = ~n10864 | ~P2_DATAO_REG_10__SCAN_IN;
  assign n16175 = n12889 ^ n12900;
  assign n12740 = ~n12896 | ~n12893;
  assign n15057 = ~n11663;
  assign n9814 = ~n9813 | ~n9812;
  assign n11653 = ~n11833;
  assign n11660 = ~n10115 & ~n10962;
  assign n10107 = ~n13165 | ~n13308;
  assign n14147 = n10341 ^ SI_30_;
  assign n13997 = n10336 ^ SI_29_;
  assign n10897 = n10331 ^ SI_28_;
  assign n10690 = n10326 ^ SI_27_;
  assign n10610 = n9708 ^ SI_22_;
  assign n10592 = n9703 ^ SI_21_;
  assign n10575 = n9698 ^ SI_20_;
  assign n10415 = ~n9272 | ~n9271;
  assign n9272 = ~n10364 | ~n10362;
  assign n11615 = n10241 ^ n10240;
  assign n9218 = ~SI_11_;
  assign n9629 = ~n9215 & ~n9214;
  assign n9214 = ~n9213;
  assign n9215 = ~n9611 & ~n9610;
  assign n9587 = ~n9563 & ~n9198;
  assign n9198 = ~n9197;
  assign n9586 = n9202 ^ SI_9_;
  assign n9021 = ~n9002 & ~n13303;
  assign n9548 = ~n11039 | ~n8921;
  assign n12550 = ~n12548 & ~n12547;
  assign n12199 = n15591 ^ n16507;
  assign n14321 = n16695 ^ ~n15591;
  assign n15595 = n15591 ^ ~n16778;
  assign n15583 = ~n10689 & ~n10688;
  assign n15582 = n15595 ^ n16779;
  assign n14624 = ~n10591 & ~n14472;
  assign n15142 = ~n10665 & ~n10664;
  assign n15141 = n16759 ^ n10680;
  assign n9352 = ~P2_REG3_REG_4__SCAN_IN;
  assign n10165 = ~n10226;
  assign n15603 = ~n15355;
  assign n13714 = ~n16461;
  assign n13466 = n16461 ^ ~n15591;
  assign n13468 = ~n10214 | ~n10213;
  assign n10214 = ~n13348 | ~n10211;
  assign n9365 = ~P2_REG3_REG_11__SCAN_IN;
  assign n14162 = n16679 ^ n15591;
  assign n14164 = ~n10538 | ~n10537;
  assign n10538 = ~n14043 | ~n10535;
  assign n10536 = ~n14041;
  assign n9392 = ~n9391 | ~n9649;
  assign n9395 = ~n16960;
  assign n15604 = ~n9364 & ~n11754;
  assign n9657 = ~n11885 | ~n9655;
  assign n16948 = ~n16946;
  assign n10698 = ~n13434 | ~P2_REG2_REG_27__SCAN_IN;
  assign n10490 = ~n13431 | ~P2_REG1_REG_26__SCAN_IN;
  assign n10673 = ~n10669 | ~n10668;
  assign n10633 = ~n10629 | ~n10628;
  assign n10652 = ~n10649 | ~n10648;
  assign n10618 = ~n13431 | ~P2_REG1_REG_22__SCAN_IN;
  assign n10603 = ~n10600 | ~n10599;
  assign n10568 = ~n10565 | ~n10564;
  assign n10532 = ~n10529 | ~n10528;
  assign n9486 = ~n9485 | ~n9484;
  assign n9464 = ~n13430 | ~P2_REG0_REG_3__SCAN_IN;
  assign n9144 = ~n9108 | ~n11348;
  assign n9095 = ~n9093 | ~P2_REG1_REG_1__SCAN_IN;
  assign n11416 = n9135 ^ n9450;
  assign n11858 = n11860 ^ n11872;
  assign n11874 = P2_REG2_REG_6__SCAN_IN ^ n11872;
  assign n11319 = ~n16958;
  assign n12529 = n12536 ^ n12528;
  assign n13030 = P2_REG1_REG_10__SCAN_IN ^ n13052;
  assign n13269 = n13276 ^ n13268;
  assign n13056 = ~P2_REG2_REG_10__SCAN_IN | ~n13052;
  assign n13767 = P2_REG1_REG_12__SCAN_IN ^ ~n13779;
  assign n14027 = n14034 ^ n14026;
  assign n14576 = P2_REG1_REG_14__SCAN_IN ^ n14598;
  assign n14710 = n14717 ^ n14709;
  assign n15179 = P2_REG1_REG_16__SCAN_IN ^ n15206;
  assign n14704 = n15190 ^ n15189;
  assign n15282 = n15281 ^ n15280;
  assign n15374 = P2_REG2_REG_18__SCAN_IN ^ n15381;
  assign n15389 = n8926 ^ P2_REG1_REG_19__SCAN_IN;
  assign n15367 = n15381 ^ P2_REG1_REG_18__SCAN_IN;
  assign n15385 = n8926 ^ ~P2_REG2_REG_19__SCAN_IN;
  assign n15376 = ~P2_REG2_REG_18__SCAN_IN | ~n15381;
  assign n15460 = P2_REG3_REG_26__SCAN_IN ^ ~n10498;
  assign n16659 = ~n16658;
  assign n14101 = P2_REG3_REG_17__SCAN_IN ^ n10527;
  assign n14071 = ~n14075;
  assign n12662 = ~n16523;
  assign n9438 = ~n8921 | ~n11007;
  assign n9439 = ~n9433 & ~n9432;
  assign n9417 = ~n9413 | ~n9412;
  assign n9413 = ~n13430 | ~P2_REG0_REG_1__SCAN_IN;
  assign n11525 = n11524 ^ n11531;
  assign n16387 = n16900 ^ ~n16406;
  assign n16348 = ~n16779 | ~n16345;
  assign n15467 = n16894 ^ n15574;
  assign n15017 = n16901 ^ n15247;
  assign n14863 = n16895 ^ ~n15003;
  assign n14849 = ~n14848 | ~n14847;
  assign n14794 = n16892 ^ ~n14853;
  assign n16723 = ~n10596 & ~n10595;
  assign n14299 = n14284 ^ ~n16884;
  assign n13976 = n16880 ^ ~n14084;
  assign n13745 = n16878 ^ n13959;
  assign n13866 = n13865 ^ ~n13864;
  assign n13650 = n16874 ^ ~n13716;
  assign n13332 = ~n13389 | ~n16410;
  assign n9621 = ~n10558 | ~n13041;
  assign n13129 = ~n13315;
  assign n13132 = n16866 ^ n13102;
  assign n11887 = ~n11886;
  assign n9391 = ~n9021 & ~n16956;
  assign n9346 = ~P2_IR_REG_29__SCAN_IN;
  assign n8988 = ~n8987 & ~n8986;
  assign n9338 = ~P2_IR_REG_17__SCAN_IN;
  assign n15184 = n10522 ^ P2_IR_REG_17__SCAN_IN;
  assign n15192 = n10512 ^ P2_IR_REG_16__SCAN_IN;
  assign n14698 = n10510 ^ P2_IR_REG_15__SCAN_IN;
  assign n14015 = n10221 ^ n10220;
  assign n10205 = ~P2_IR_REG_12__SCAN_IN;
  assign n9614 = ~n9617 | ~P2_IR_REG_31__SCAN_IN;
  assign n11628 = n9494 ^ P2_IR_REG_5__SCAN_IN;
  assign n9157 = n9096 ^ P2_IR_REG_2__SCAN_IN;
  assign n15509 = ~n10884 | ~n10883;
  assign n10881 = ~n10880;
  assign n15510 = n10914 ^ ~n10913;
  assign n10841 = ~n15087 | ~n10831;
  assign n10859 = ~n10858;
  assign n10860 = ~n10857;
  assign n15738 = ~n12349;
  assign n12434 = ~n12437 | ~n12325;
  assign n14056 = n10436 ^ n10435;
  assign n9898 = ~n9882;
  assign n12086 = n9873 ^ n9872;
  assign n9990 = ~n9988;
  assign n10146 = n10144 & n10143;
  assign n14724 = ~n10744 & ~n14434;
  assign n10744 = ~n14437 & ~n14435;
  assign n10278 = ~n10277;
  assign n10025 = ~P2_DATAO_REG_11__SCAN_IN;
  assign n15829 = ~n15820;
  assign n13512 = n13511 ^ ~n13510;
  assign n9803 = ~n11723 | ~n11724;
  assign n11744 = ~n9822 | ~n9821;
  assign n11745 = ~n9824 | ~n9823;
  assign n10727 = ~n10465 | ~n10464;
  assign n10144 = ~n11835 & ~n11661;
  assign n12439 = ~n9914 | ~n9913;
  assign n16318 = ~n16317;
  assign n16224 = ~n16324;
  assign n16331 = ~n11658 | ~n11911;
  assign n10894 = ~n10891 | ~n10890;
  assign n10805 = ~n8923 | ~P1_REG0_REG_24__SCAN_IN;
  assign n10819 = ~n8923 | ~P1_REG0_REG_23__SCAN_IN;
  assign n10752 = ~n10749 | ~n10748;
  assign n10457 = ~n10456 | ~n10455;
  assign n10155 = ~n8923 | ~P1_REG0_REG_13__SCAN_IN;
  assign n11241 = ~n11240 | ~n11239;
  assign n11300 = n11211 ^ P1_REG1_REG_9__SCAN_IN;
  assign n11597 = P1_REG2_REG_11__SCAN_IN ^ ~n11609;
  assign n11504 = P1_REG1_REG_11__SCAN_IN ^ n11609;
  assign n12561 = n12564 ^ ~P1_REG1_REG_14__SCAN_IN;
  assign n11197 = ~n10972 | ~n10980;
  assign n15126 = P1_REG1_REG_19__SCAN_IN ^ n15125;
  assign n10716 = ~n10713 | ~n10712;
  assign n15104 = n15061 ^ n15307;
  assign n15430 = P1_REG3_REG_26__SCAN_IN ^ n10869;
  assign n15042 = P1_REG3_REG_25__SCAN_IN ^ n10847;
  assign n15070 = ~n15653;
  assign n15091 = P1_REG3_REG_23__SCAN_IN ^ n10818;
  assign n15952 = ~n10815 & ~n10814;
  assign n14398 = ~n16112;
  assign n15936 = ~n10782 & ~n10781;
  assign n13938 = n13928 & n13927;
  assign n14116 = ~n14060;
  assign n13607 = n16185 ^ n13567;
  assign n15826 = ~n15819;
  assign n12953 = n16177 ^ n13063;
  assign n11841 = ~n11835 & ~n11834;
  assign n15684 = ~n9790 & ~n9789;
  assign n15318 = ~n15520 | ~n15484;
  assign n14954 = n15054 ^ n15055;
  assign n14832 = ~n15969 | ~n15533;
  assign n14880 = n16202 ^ ~n14926;
  assign n14239 = n14238 ^ n16196;
  assign n13987 = ~n13985 | ~n16367;
  assign n13986 = ~n15880 | ~n16369;
  assign n13940 = ~n13938 | ~n16367;
  assign n13939 = ~n14059 | ~n16369;
  assign n13192 = ~n13191 | ~n13548;
  assign n13193 = ~n13547;
  assign n13170 = n16179 ^ ~n13140;
  assign n13153 = ~n13152 | ~n13151;
  assign n12955 = ~n12904 | ~n12903;
  assign n12904 = ~n12899 | ~n15637;
  assign n12892 = ~n14669;
  assign n12038 = ~n15714;
  assign n11675 = ~n11660 & ~n11659;
  assign n10961 = ~n10111 | ~n10116;
  assign n11674 = ~n10119 & ~n10118;
  assign n10984 = ~n11658;
  assign n15585 = n10898 ^ ~n10897;
  assign n10691 = ~n10690;
  assign n8958 = ~P1_IR_REG_25__SCAN_IN;
  assign n10114 = n8970 ^ P1_IR_REG_25__SCAN_IN;
  assign n9720 = ~n10638 | ~n10636;
  assign n10636 = n9718 ^ SI_24_;
  assign n9710 = ~n10611 | ~n10610;
  assign n10641 = n9713 ^ SI_23_;
  assign n16236 = ~n9011 & ~n9010;
  assign n9010 = ~n9012;
  assign n12785 = n10593 ^ ~n10592;
  assign n12181 = ~n12176;
  assign n14755 = n10418 ^ P1_IR_REG_17__SCAN_IN;
  assign n11962 = n10415 ^ n10414;
  assign n14457 = n10369 ^ ~P1_IR_REG_16__SCAN_IN;
  assign n11804 = n10364 ^ ~n10363;
  assign n13840 = n10390 ^ ~P1_IR_REG_15__SCAN_IN;
  assign n10390 = ~n10389 | ~P1_IR_REG_31__SCAN_IN;
  assign n11714 = n10189 ^ ~n10188;
  assign n13487 = n10388 ^ n10387;
  assign n12571 = n10266 ^ P1_IR_REG_13__SCAN_IN;
  assign n11519 = n10217 ^ ~n10216;
  assign n12158 = n10058 ^ ~P1_IR_REG_12__SCAN_IN;
  assign n10058 = ~n10265 | ~P1_IR_REG_31__SCAN_IN;
  assign n11262 = n9629 ^ n9628;
  assign n11163 = n9611 ^ n9610;
  assign n11114 = n9587 ^ n9586;
  assign n11282 = n9945 ^ n9944;
  assign n9945 = ~n9968 | ~P1_IR_REG_31__SCAN_IN;
  assign n11054 = ~P2_DATAO_REG_8__SCAN_IN;
  assign n9185 = ~n9512 | ~n9511;
  assign n9540 = n9188 ^ SI_7_;
  assign n11251 = n9916 ^ P1_IR_REG_6__SCAN_IN;
  assign n10991 = n9512 ^ ~n9511;
  assign n9071 = ~n9477 | ~n9478;
  assign n9176 = n9178 ^ SI_5_;
  assign n11044 = n9460 ^ ~n9459;
  assign n9460 = ~n9458 | ~n9457;
  assign n11009 = ~P2_DATAO_REG_2__SCAN_IN;
  assign n12825 = ~n9577 | ~n9553;
  assign n15355 = ~n9364 & ~n11539;
  assign n13596 = n13595 ^ n13594;
  assign n15215 = n15328 ^ ~n15338;
  assign n15222 = ~n15334 | ~n15604;
  assign n13419 = ~n9357 | ~n9379;
  assign n9644 = ~n9643 | ~n9642;
  assign n13418 = ~n13416 | ~n13415;
  assign n12301 = ~P2_REG3_REG_3__SCAN_IN;
  assign n14324 = n14323 ^ ~n14322;
  assign n14322 = n14321 ^ ~n16696;
  assign n14331 = ~n14330 | ~n14329;
  assign n15611 = ~n15610 | ~n15609;
  assign n9604 = ~n9597 | ~n9596;
  assign n12429 = n9428 ^ n16475;
  assign n9427 = ~n10646 | ~n11540;
  assign n14652 = n10598 ^ n10597;
  assign n14625 = n14624 ^ ~n14623;
  assign n14623 = n14622 ^ ~n16721;
  assign n15143 = n15142 ^ ~n15141;
  assign n15150 = ~n15239 | ~n15602;
  assign n13901 = n13900 ^ ~n13899;
  assign n14044 = n14043 ^ ~n14042;
  assign n14042 = n14041 ^ ~n16669;
  assign n15337 = n15336 ^ ~n15335;
  assign n15335 = n15334 ^ ~n15333;
  assign n15347 = ~n16759 | ~n15604;
  assign n9507 = ~n9500 | ~n9499;
  assign n9506 = ~n9505 | ~n9504;
  assign n12981 = ~n9600 | ~n9599;
  assign n12972 = ~n12971 | ~n12970;
  assign n14476 = n14475 ^ ~n14474;
  assign n14483 = ~n14482 | ~n14481;
  assign n14805 = n14804 ^ ~n16734;
  assign n14810 = ~n15602 | ~n14808;
  assign n14165 = n14164 ^ ~n14163;
  assign n14163 = n14162 ^ ~n16676;
  assign n14173 = ~n14172 | ~n14171;
  assign n16550 = ~n13015;
  assign n15596 = ~n9653 & ~n9652;
  assign n9651 = ~n11885 | ~n11537;
  assign n10256 = n10505 ^ ~n10506;
  assign n10257 = ~n16642 | ~n15342;
  assign n10585 = ~n10671 & ~n10584;
  assign n10551 = ~n10548 | ~n10547;
  assign n10170 = ~n10168 | ~n10167;
  assign n16645 = ~n13960;
  assign n10233 = n10232 & n10231;
  assign n10231 = ~n13430 | ~P2_REG0_REG_13__SCAN_IN;
  assign n9374 = n9373 & n9372;
  assign n13325 = ~n13101;
  assign n9581 = n9580 & n9579;
  assign n9535 = n9531 & n9530;
  assign n12402 = ~n16522;
  assign n9441 = ~n13430 | ~P2_REG0_REG_2__SCAN_IN;
  assign n13429 = ~P2_U3893;
  assign n12110 = n9570 ^ P2_IR_REG_8__SCAN_IN;
  assign n9125 = ~n9123 | ~n16958;
  assign n9123 = ~n11322;
  assign n12537 = n12536 ^ n12535;
  assign n13054 = P2_REG2_REG_10__SCAN_IN ^ n13052;
  assign n13277 = n13276 ^ n13275;
  assign n13791 = P2_REG2_REG_12__SCAN_IN ^ ~n13779;
  assign n14600 = P2_REG2_REG_14__SCAN_IN ^ n14598;
  assign n15208 = P2_REG2_REG_16__SCAN_IN ^ n15206;
  assign n15378 = ~n11322 & ~n9344;
  assign n15273 = n15267 & n15266;
  assign n15285 = n15367 ^ ~n15366;
  assign n15255 = n15374 ^ ~n15373;
  assign n15395 = n15393 ^ ~n15392;
  assign n15372 = n15389 ^ n15370;
  assign n15380 = n15385 ^ n15377;
  assign n16359 = ~n16358 | ~n16357;
  assign n15626 = n16353 ^ n15578;
  assign n13744 = ~n16419 | ~n16410;
  assign n15290 = n16910 ^ ~n15451;
  assign n13382 = ~n13381 | ~n15557;
  assign n13381 = n13380 ^ ~n13647;
  assign n13370 = ~n13369 | ~n13368;
  assign n13115 = ~n13233 | ~n16410;
  assign n12938 = ~n12821 | ~n12820;
  assign n12782 = ~n12779 | ~n12778;
  assign n12649 = ~n12646 | ~n12645;
  assign n11531 = ~n9324 & ~n9323;
  assign n9738 = n8999 ^ P2_IR_REG_26__SCAN_IN;
  assign n8999 = ~n9085 & ~n10520;
  assign n10541 = ~n10540 | ~P2_IR_REG_31__SCAN_IN;
  assign n15206 = ~n15192;
  assign n9634 = ~n10204;
  assign n12518 = n9591 ^ P2_IR_REG_9__SCAN_IN;
  assign n12012 = n9544 ^ n9543;
  assign n11585 = ~n11628;
  assign n11570 = n9139 ^ P2_IR_REG_4__SCAN_IN;
  assign n11418 = n9134 ^ ~P2_IR_REG_3__SCAN_IN;
  assign n11002 = ~n9157;
  assign n11356 = n9090 ^ ~P2_IR_REG_1__SCAN_IN;
  assign n10980 = ~n10121 | ~n10135;
  assign n10133 = ~n10121;
  assign n12847 = ~n12375;
  assign n15527 = ~n15517 | ~n15516;
  assign n15524 = ~n15523 | ~n15522;
  assign n10303 = n10302 ^ n10358;
  assign n15090 = n15089 ^ ~n15088;
  assign n13292 = n13291 ^ n13290;
  assign n14438 = n14437 ^ ~n14436;
  assign n14445 = ~n14444 | ~n14443;
  assign n14444 = ~n14442 & ~n14441;
  assign n12877 = ~n12876 | ~n12875;
  assign n12875 = ~n12874 | ~n15511;
  assign n14735 = P1_REG3_REG_21__SCAN_IN ^ n10764;
  assign n14734 = n14733 ^ ~n14732;
  assign n10124 = n10262 ^ n10078;
  assign n14133 = n14132 ^ ~n14131;
  assign n14131 = n14130 ^ ~n14129;
  assign n14058 = P1_REG3_REG_17__SCAN_IN ^ n10452;
  assign n14057 = n14056 ^ n14055;
  assign n15165 = n15164 ^ n15163;
  assign n10009 = ~n10004 | ~n10003;
  assign n10008 = ~n10007 | ~n10006;
  assign n9784 = ~n9783 | ~n9782;
  assign n14609 = n10747 ^ P1_REG3_REG_20__SCAN_IN;
  assign n14608 = n14724 ^ n14725;
  assign n14618 = ~n14617 | ~n14616;
  assign n14617 = ~n15915 | ~n15428;
  assign n13520 = ~n13213;
  assign n14919 = P1_REG3_REG_22__SCAN_IN ^ n10785;
  assign n14911 = n14910 ^ n14909;
  assign n10142 = ~n10144 | ~n10141;
  assign n15427 = n15425 ^ n15424;
  assign n10137 = n10136 & n16328;
  assign n10136 = ~n10134 | ~P1_STATE_REG_SCAN_IN;
  assign n10134 = ~n11644 | ~n10133;
  assign n14111 = n14110 ^ ~n14125;
  assign n10808 = n10803 & n10802;
  assign n10822 = n10817 & n10816;
  assign n10789 = n10784 & n10783;
  assign n10768 = n10763 & n10762;
  assign n10475 = ~n10472 | ~n10471;
  assign n10428 = n10427 & n10426;
  assign n10429 = n10424 & n10423;
  assign n10311 = n10310 & n10309;
  assign n10291 = n10290 & n10289;
  assign n13076 = ~n13283;
  assign n9885 = n9884 & n9883;
  assign n9858 = n9853 & n9852;
  assign n9806 = ~n8923 | ~P1_REG0_REG_2__SCAN_IN;
  assign n15690 = ~n15683;
  assign n9760 = n9754 & n9753;
  assign n11507 = n10021 ^ n10020;
  assign n13497 = ~n13496 | ~n14114;
  assign n14766 = ~n14765 | ~n14764;
  assign n15027 = n16037 ^ ~n14974;
  assign n14981 = n16134 ^ ~n14973;
  assign n15501 = ~n15495 | ~n15654;
  assign n14873 = P1_REG3_REG_24__SCAN_IN ^ ~n10804;
  assign n14670 = n16200 ^ n14818;
  assign n14524 = n16198 ^ ~n14544;
  assign n14335 = n14184 ^ ~n16194;
  assign n14201 = ~n14336 | ~n15659;
  assign n13071 = ~n13070 | ~n13069;
  assign n13069 = ~n13241 | ~n14547;
  assign n11918 = ~n11922;
  assign n16382 = ~n16376 | ~n16375;
  assign n13757 = ~n13756 | ~n13755;
  assign n13627 = ~n13626;
  assign n13624 = ~n13623 | ~n13622;
  assign n12604 = ~n12601 | ~n12600;
  assign n12388 = ~n12694 | ~n12385;
  assign n12272 = ~n12269 | ~n12268;
  assign n12359 = ~n12716 | ~n12356;
  assign n10349 = n10348 ^ SI_31_;
  assign n14155 = ~n14890;
  assign n14005 = ~n9752 | ~n9751;
  assign n9751 = ~n10353;
  assign n13880 = ~n15585;
  assign n13459 = ~n9736 | ~n9735;
  assign n9736 = ~n10323;
  assign n13308 = ~n10114;
  assign n13452 = n10677 ^ n10676;
  assign n16328 = ~n10968 | ~P1_STATE_REG_SCAN_IN;
  assign n13124 = n10642 ^ ~n10641;
  assign n16324 = n9762 ^ P1_IR_REG_20__SCAN_IN;
  assign n12315 = n9692 ^ n9286;
  assign n14754 = ~n15132;
  assign n12564 = ~n13487;
  assign n11600 = ~n12158;
  assign n10055 = ~n10052;
  assign n11609 = n10024 ^ n10023;
  assign n10022 = ~n10021 | ~n10020;
  assign n11299 = n9969 ^ P1_IR_REG_9__SCAN_IN;
  assign n9566 = ~n9565 | ~n9564;
  assign n9567 = ~n9563;
  assign n11492 = n9920 ^ P1_IR_REG_7__SCAN_IN;
  assign n9919 = ~n9918 | ~n9917;
  assign n11039 = n9541 ^ n9540;
  assign n11473 = n9072 ^ ~P1_IR_REG_5__SCAN_IN;
  assign n10996 = n9176 ^ ~n9177;
  assign n11007 = ~n11001;
  assign n10953 = ~n9667 | ~n9666;
  assign n9672 = ~n10967 | ~n10966;
  assign P2_U3893 = ~n9101 & ~P2_U3151;
  assign n10710 = ~n10504 | ~n10503;
  assign n9660 = ~n9659 | ~n9658;
  assign n15363 = ~n15357 | ~n15356;
  assign n13163 = ~P2_U3893 | ~n15589;
  assign n13796 = ~n13788 & ~n13787;
  assign n14039 = ~n14038 | ~n15378;
  assign n14604 = ~n15378 | ~n14603;
  assign n14603 = P2_REG2_REG_15__SCAN_IN ^ ~n14718;
  assign n14721 = n15208 ^ ~n15207;
  assign n15211 = P2_REG2_REG_17__SCAN_IN ^ ~n15252;
  assign n14573 = ~n14572 & ~n14571;
  assign n14432 = ~n14572 & ~n14431;
  assign n14655 = ~n14654 | ~n14653;
  assign n14510 = ~n14509 | ~n14508;
  assign n14384 = ~n14383 | ~n14382;
  assign n13752 = ~n13743 | ~n13742;
  assign n13393 = ~n13392 | ~n13391;
  assign n13450 = ~n16442 | ~n13449;
  assign n13340 = ~n16442 | ~n13339;
  assign n13239 = ~n16442 | ~n13238;
  assign n13447 = ~n16438 | ~n13449;
  assign n13337 = ~n16438 | ~n13339;
  assign n13236 = ~n16438 | ~n13238;
  assign n12654 = ~n12652 | ~n14351;
  assign n10942 = ~n10919 | ~n10918;
  assign n10486 = ~n10485 | ~n10484;
  assign n15139 = ~n15138 | ~n15137;
  assign n15138 = n8924 ^ n15136;
  assign n14253 = ~n14252 | ~n14251;
  assign n14269 = ~n14268 | ~n14267;
  assign n13824 = ~n13823 | ~n13822;
  assign n13933 = ~n13932 | ~n13931;
  assign n13227 = ~n13225 | ~n13224;
  assign n13162 = ~n13156 | ~n13226;
  assign n13208 = ~n16381 | ~n13210;
  assign n13251 = ~n16381 | ~n13250;
  assign n13180 = ~n16381 | ~n13179;
  assign n13211 = ~n16377 | ~n13210;
  assign n13248 = ~n16377 | ~n13250;
  assign n13177 = ~n16377 | ~n13179;
  assign n12913 = ~n16377 | ~n12915;
  assign n13169 = ~n13301 | ~n14154;
  assign n12887 = ~n12882 | ~n14154;
  assign n9332 = ~n10219 & ~P2_IR_REG_13__SCAN_IN;
  assign n16021 = ~n16045;
  assign n13226 = ~n15323;
  assign n8934 = ~n11197 & ~n14900;
  assign n16401 = ~n8932;
  assign n15707 = ~n15717;
  assign n16554 = ~n16553;
  assign n16564 = ~n16563;
  assign n16575 = ~n16574;
  assign n16623 = ~n16621;
  assign n16657 = ~n16658 | ~n16798;
  assign n16699 = ~n16708;
  assign n16048 = ~n16047;
  assign n13646 = ~n13645;
  assign n9471 = ~n12199;
  assign n11582 = ~n11570;
  assign n9386 = ~n11537;
  assign n9940 = ~n9937;
  assign n9559 = ~n9558;
  assign n9542 = ~P1_DATAO_REG_7__SCAN_IN;
  assign n9093 = ~n11344;
  assign n15554 = ~n15555;
  assign n10558 = ~n14426;
  assign n9612 = ~P2_IR_REG_9__SCAN_IN;
  assign n12587 = ~n16077;
  assign n10236 = ~n13466;
  assign n14636 = ~n14773;
  assign n16594 = ~n13362;
  assign n15229 = ~n14997 & ~n16901;
  assign n14638 = ~n14490 & ~n14489;
  assign n9987 = ~n9989;
  assign n10126 = ~n11843;
  assign n15696 = ~n15715;
  assign n9195 = ~n9194;
  assign n10687 = ~n10686;
  assign n10650 = ~P2_REG1_REG_23__SCAN_IN;
  assign n10530 = ~P2_REG1_REG_17__SCAN_IN;
  assign n14787 = ~n14785 | ~n16890;
  assign n16405 = n16404 ^ n16903;
  assign n16730 = ~n10614 & ~n10613;
  assign n13870 = ~n16628;
  assign n9821 = ~n9823;
  assign n10462 = ~n10464;
  assign n10863 = ~n10862;
  assign n14926 = ~n14820 | ~n14819;
  assign n11668 = ~n11910;
  assign n9225 = ~n9222 | ~n9628;
  assign n9944 = ~P1_IR_REG_8__SCAN_IN;
  assign n9457 = ~n9456;
  assign n9003 = ~n9077 | ~n9078;
  assign n12793 = ~n12407;
  assign n16410 = ~n11763 & ~n8926;
  assign n14428 = ~n16412;
  assign n15625 = ~n16386;
  assign n8972 = ~n9012 & ~P1_IR_REG_22__SCAN_IN;
  assign n14129 = ~n10408;
  assign n15835 = ~n15839;
  assign n10141 = ~n10140;
  assign n16130 = ~n16018;
  assign n14402 = ~n14399 & ~n16196;
  assign n14235 = ~n16107;
  assign n11249 = ~P1_REG3_REG_6__SCAN_IN;
  assign n12484 = ~n12479;
  assign n9477 = ~n9066 | ~n9065;
  assign n9004 = ~n9003 | ~P2_IR_REG_31__SCAN_IN;
  assign n9600 = ~n9356;
  assign n11852 = ~P2_REG3_REG_7__SCAN_IN;
  assign n13741 = ~P2_REG2_REG_15__SCAN_IN;
  assign n11989 = ~n11527 & ~n11526;
  assign n14000 = ~P1_DATAO_REG_29__SCAN_IN;
  assign n15776 = ~n15772;
  assign n10353 = ~n9746 & ~P1_IR_REG_29__SCAN_IN;
  assign n13461 = ~P2_DATAO_REG_26__SCAN_IN;
  assign n12733 = ~P2_DATAO_REG_21__SCAN_IN;
  assign n13490 = ~n13840;
  assign n11359 = ~n11203;
  assign n11658 = ~n10121 & ~n10120;
  assign n12882 = ~n12976;
  assign n8936 = ~P1_IR_REG_11__SCAN_IN & ~P1_IR_REG_10__SCAN_IN;
  assign n8935 = ~P1_IR_REG_8__SCAN_IN & ~P1_IR_REG_9__SCAN_IN;
  assign n8940 = ~n8936 | ~n8935;
  assign n8938 = ~P1_IR_REG_6__SCAN_IN & ~P1_IR_REG_5__SCAN_IN;
  assign n8937 = ~P1_IR_REG_7__SCAN_IN & ~P1_IR_REG_4__SCAN_IN;
  assign n8939 = ~n8938 | ~n8937;
  assign n8944 = ~n8940 & ~n8939;
  assign n8941 = ~P1_IR_REG_1__SCAN_IN;
  assign n9811 = ~n11382 | ~n8941;
  assign n9833 = ~P1_IR_REG_2__SCAN_IN;
  assign n8942 = ~P1_IR_REG_3__SCAN_IN;
  assign n9859 = ~n9811 & ~n8943;
  assign n8946 = ~P1_IR_REG_12__SCAN_IN & ~P1_IR_REG_14__SCAN_IN;
  assign n8945 = ~P1_IR_REG_15__SCAN_IN & ~P1_IR_REG_17__SCAN_IN;
  assign n8947 = ~P1_IR_REG_16__SCAN_IN & ~P1_IR_REG_13__SCAN_IN;
  assign n8948 = ~n8947 | ~n10445;
  assign n9005 = ~n9761 & ~P1_IR_REG_20__SCAN_IN;
  assign n8952 = ~n8972 | ~n8954;
  assign n13165 = n8953 ^ P1_IR_REG_24__SCAN_IN;
  assign n9013 = ~P1_IR_REG_22__SCAN_IN;
  assign n8955 = ~n8954 | ~n9013;
  assign n8957 = ~n8955 & ~P1_IR_REG_24__SCAN_IN;
  assign n8956 = ~P1_IR_REG_21__SCAN_IN & ~P1_IR_REG_20__SCAN_IN;
  assign n8966 = ~n8957 | ~n8956;
  assign n8969 = ~n9761 & ~n8966;
  assign n8967 = ~n8966 & ~n8965;
  assign n9017 = ~n9287 | ~n8967;
  assign n13460 = ~n8968 | ~n9017;
  assign n8971 = ~n10116 | ~n10114;
  assign n10121 = ~n13165 & ~n8971;
  assign n8976 = ~P2_IR_REG_11__SCAN_IN & ~P2_IR_REG_12__SCAN_IN;
  assign n8977 = ~n8976 | ~n8975;
  assign n8982 = ~n9493 & ~n8977;
  assign n8978 = ~P2_IR_REG_5__SCAN_IN & ~P2_IR_REG_6__SCAN_IN;
  assign n8980 = ~n9491 | ~n8978;
  assign n9589 = ~n8979 | ~n9543;
  assign n9080 = ~n9332 | ~n8988;
  assign n9077 = ~n9080 & ~P2_IR_REG_21__SCAN_IN;
  assign n8991 = ~n9003 & ~n8990;
  assign n8992 = ~n8991 & ~n10520;
  assign n8998 = ~n8997 | ~n8996;
  assign n9085 = ~n9080 & ~n8998;
  assign n9000 = ~n9003 & ~P2_IR_REG_23__SCAN_IN;
  assign n9007 = ~n9005 & ~n10417;
  assign n9009 = ~n9007 & ~n9006;
  assign n11667 = ~n16236 | ~n16149;
  assign n9744 = ~n9017 & ~P1_IR_REG_27__SCAN_IN;
  assign n9016 = ~n9744 & ~n10417;
  assign n11686 = n9016 ^ P1_IR_REG_28__SCAN_IN;
  assign n9018 = ~n9017 | ~P1_IR_REG_31__SCAN_IN;
  assign n9022 = n13303 ^ ~P2_B_REG_SCAN_IN;
  assign P2_U3241 = n9024 & P2_D_REG_24__SCAN_IN;
  assign P2_U3243 = n9024 & P2_D_REG_22__SCAN_IN;
  assign P2_U3246 = n9024 & P2_D_REG_19__SCAN_IN;
  assign P2_U3240 = n9024 & P2_D_REG_25__SCAN_IN;
  assign P2_U3259 = n9024 & P2_D_REG_6__SCAN_IN;
  assign P2_U3242 = n9024 & P2_D_REG_23__SCAN_IN;
  assign P2_U3261 = n9024 & P2_D_REG_4__SCAN_IN;
  assign P2_U3262 = n9024 & P2_D_REG_3__SCAN_IN;
  assign P2_U3263 = n9024 & P2_D_REG_2__SCAN_IN;
  assign P2_U3244 = n9024 & P2_D_REG_21__SCAN_IN;
  assign P2_U3245 = n9024 & P2_D_REG_20__SCAN_IN;
  assign P2_U3239 = n9024 & P2_D_REG_26__SCAN_IN;
  assign P2_U3251 = n9024 & P2_D_REG_14__SCAN_IN;
  assign P2_U3234 = n9024 & P2_D_REG_31__SCAN_IN;
  assign P2_U3253 = n9024 & P2_D_REG_12__SCAN_IN;
  assign P2_U3254 = n9024 & P2_D_REG_11__SCAN_IN;
  assign P2_U3255 = n9024 & P2_D_REG_10__SCAN_IN;
  assign P2_U3256 = n9024 & P2_D_REG_9__SCAN_IN;
  assign P2_U3257 = n9024 & P2_D_REG_8__SCAN_IN;
  assign P2_U3258 = n9024 & P2_D_REG_7__SCAN_IN;
  assign P2_U3235 = n9024 & P2_D_REG_30__SCAN_IN;
  assign P2_U3260 = n9024 & P2_D_REG_5__SCAN_IN;
  assign P2_U3236 = n9024 & P2_D_REG_29__SCAN_IN;
  assign P2_U3237 = n9024 & P2_D_REG_28__SCAN_IN;
  assign P2_U3238 = n9024 & P2_D_REG_27__SCAN_IN;
  assign P2_U3248 = n9024 & P2_D_REG_17__SCAN_IN;
  assign P2_U3249 = n9024 & P2_D_REG_16__SCAN_IN;
  assign P2_U3250 = n9024 & P2_D_REG_15__SCAN_IN;
  assign P2_U3247 = n9024 & P2_D_REG_18__SCAN_IN;
  assign P2_U3252 = n9024 & P2_D_REG_13__SCAN_IN;
  assign n10345 = ~n9043;
  assign n9032 = ~n8919 | ~SI_0_;
  assign n9418 = n9032 ^ P1_DATAO_REG_0__SCAN_IN;
  assign n9034 = n9418 | P2_STATE_REG_SCAN_IN;
  assign n9033 = ~P2_IR_REG_0__SCAN_IN | ~P2_STATE_REG_SCAN_IN;
  assign P2_U3295 = ~n9034 | ~n9033;
  assign n9036 = ~n9043 | ~SI_0_;
  assign n9035 = ~P2_DATAO_REG_0__SCAN_IN;
  assign n9040 = ~n9036 | ~n9035;
  assign n9048 = ~n9726 & ~n9038;
  assign n9039 = ~n9048;
  assign n9763 = ~n9040 | ~n9039;
  assign n9042 = n9763 | P1_STATE_REG_SCAN_IN;
  assign n9041 = ~P1_IR_REG_0__SCAN_IN | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3355 = ~n9042 | ~n9041;
  assign n9045 = ~n8919 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n9047 = ~n9199 & ~n9046;
  assign n9050 = ~n9037 | ~P1_DATAO_REG_1__SCAN_IN;
  assign n9049 = ~n9199 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n9051 = ~n9050 | ~n9049;
  assign n9436 = ~n9408 | ~SI_1_;
  assign n9434 = ~n9053 & ~n9052;
  assign n9055 = ~n10345 & ~n11009;
  assign n9437 = ~n9055 & ~n9054;
  assign n9456 = ~n9437 & ~n9056;
  assign n9057 = ~n9434 & ~n9456;
  assign n9063 = ~n9436 | ~n9057;
  assign n9059 = ~n8919 | ~P1_DATAO_REG_3__SCAN_IN;
  assign n9064 = ~n9059 | ~n9058;
  assign n9061 = ~n9060 & ~SI_2_;
  assign n9062 = ~n9459 & ~n9061;
  assign n9066 = ~n9063 | ~n9062;
  assign n9177 = ~n9071 | ~n9070;
  assign n9076 = ~n10996 & ~n13123;
  assign n9893 = ~n9859 | ~n9860;
  assign n9072 = ~n9893 | ~P1_IR_REG_31__SCAN_IN;
  assign n9074 = ~n11473 | ~P1_STATE_REG_SCAN_IN;
  assign n13309 = n8919 & P1_U3086;
  assign n9073 = ~n13309 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n9075 = ~n9074 | ~n9073;
  assign P1_U3350 = n9076 | n9075;
  assign n16961 = n9079 ^ n9078;
  assign n9081 = ~n9080 | ~P2_IR_REG_31__SCAN_IN;
  assign n9082 = ~P2_IR_REG_27__SCAN_IN & ~P2_IR_REG_26__SCAN_IN;
  assign n9345 = ~n9085 | ~n9082;
  assign n9083 = ~n9345 | ~P2_IR_REG_31__SCAN_IN;
  assign n9086 = ~n9085 | ~n9084;
  assign n9090 = ~P2_IR_REG_31__SCAN_IN | ~P2_IR_REG_0__SCAN_IN;
  assign n11327 = ~P2_IR_REG_0__SCAN_IN;
  assign n9091 = ~P2_REG1_REG_0__SCAN_IN | ~n11327;
  assign n9092 = ~n11356 | ~n9091;
  assign n9097 = n9131 ^ n9130;
  assign n9105 = ~n15182 & ~n9097;
  assign n9099 = ~n9098;
  assign n9100 = ~n9099 & ~P2_U3151;
  assign n9103 = ~P2_ADDR_REG_2__SCAN_IN | ~n15398;
  assign n9102 = ~P2_REG3_REG_2__SCAN_IN | ~P2_U3151;
  assign n9104 = ~n9103 | ~n9102;
  assign n9111 = ~n9105 & ~n9104;
  assign n11991 = ~P2_REG2_REG_0__SCAN_IN;
  assign n9106 = n11991 | P2_IR_REG_0__SCAN_IN;
  assign n11349 = ~n11356 | ~n9106;
  assign n9108 = ~n11349 | ~P2_REG2_REG_1__SCAN_IN;
  assign n11348 = ~n9107 | ~P2_REG2_REG_0__SCAN_IN;
  assign n9109 = n9145 ^ ~n9144;
  assign n9110 = ~n15378 | ~n9109;
  assign n9129 = ~n9111 | ~n9110;
  assign n9113 = ~n15386 | ~P2_REG2_REG_1__SCAN_IN;
  assign n9112 = ~n15388 | ~P2_REG1_REG_1__SCAN_IN;
  assign n9116 = ~n9113 | ~n9112;
  assign n11342 = n9116 ^ ~n11356;
  assign n9115 = ~n15386 | ~P2_REG2_REG_0__SCAN_IN;
  assign n9114 = ~n15388 | ~P2_REG1_REG_0__SCAN_IN;
  assign n11316 = ~n9115 | ~n9114;
  assign n11341 = ~n11316 & ~n11327;
  assign n9119 = ~n11342 | ~n11341;
  assign n9117 = ~n9116;
  assign n9118 = ~n9117 | ~n11356;
  assign n9121 = ~n15386 | ~P2_REG2_REG_2__SCAN_IN;
  assign n9120 = ~n15388 | ~P2_REG1_REG_2__SCAN_IN;
  assign n9154 = n9156 ^ ~n9157;
  assign n9122 = n9155 ^ ~n9154;
  assign n9127 = ~n9122 | ~n15394;
  assign n9124 = ~P2_U3893 | ~n11319;
  assign n15396 = ~n9125 | ~n9124;
  assign n9126 = ~n15396 | ~n9157;
  assign n9128 = ~n9127 | ~n9126;
  assign P2_U3184 = n9129 | n9128;
  assign n9140 = n11569 ^ ~n11567;
  assign n9143 = ~n15182 & ~n9140;
  assign n12465 = ~P2_REG3_REG_4__SCAN_IN | ~P2_U3151;
  assign n9141 = ~n15398 | ~P2_ADDR_REG_4__SCAN_IN;
  assign n9142 = ~n12465 | ~n9141;
  assign n9153 = ~n9143 & ~n9142;
  assign n9151 = n11581 ^ ~n11580;
  assign n9152 = ~n15378 | ~n9151;
  assign n9175 = ~n9153 | ~n9152;
  assign n9160 = ~n9155 | ~n9154;
  assign n9158 = ~n9156;
  assign n9159 = ~n9158 | ~n9157;
  assign n9163 = n15388 & P2_REG1_REG_3__SCAN_IN;
  assign n9161 = ~P2_REG2_REG_3__SCAN_IN;
  assign n9162 = ~n15388 & ~n9161;
  assign n9164 = ~n9163 & ~n9162;
  assign n9166 = ~n9164 | ~n11418;
  assign n9165 = ~n9164;
  assign n11425 = ~n9166 | ~n9167;
  assign n9168 = ~n9167;
  assign n9170 = ~n15386 | ~P2_REG2_REG_4__SCAN_IN;
  assign n9169 = ~n15388 | ~P2_REG1_REG_4__SCAN_IN;
  assign n9171 = n11553 ^ ~n11552;
  assign n9173 = ~n9171 | ~n15394;
  assign n9172 = ~n15396 | ~n11570;
  assign n9174 = ~n9173 | ~n9172;
  assign P2_U3186 = n9175 | n9174;
  assign n9180 = ~n9177 | ~n9176;
  assign n9541 = ~n9185 | ~n9184;
  assign n9190 = ~n9541 | ~n9540;
  assign n9565 = ~n9190 | ~n9189;
  assign n9611 = ~n9204 | ~n9203;
  assign n10052 = ~n9225 | ~n9224;
  assign n9227 = n8919 & P1_DATAO_REG_12__SCAN_IN;
  assign n10217 = ~n10057 | ~n9233;
  assign n9236 = n8919 & P1_DATAO_REG_13__SCAN_IN;
  assign n9238 = ~n9236 & ~n9235;
  assign n9241 = ~n9239 & ~SI_13_;
  assign n10215 = ~n9240 & ~n9241;
  assign n9243 = ~n10217 | ~n10215;
  assign n10241 = ~n9243 | ~n9242;
  assign n9247 = ~n9245 & ~n9244;
  assign n9250 = ~n9248 & ~SI_14_;
  assign n9252 = ~n10241 | ~n10239;
  assign n10189 = ~n9252 | ~n9251;
  assign n9255 = n8919 & P1_DATAO_REG_15__SCAN_IN;
  assign n9257 = ~n9255 & ~n9254;
  assign n9260 = ~n9258 & ~SI_15_;
  assign n10187 = ~n9259 & ~n9260;
  assign n9262 = ~n10189 | ~n10187;
  assign n9265 = n8919 & P1_DATAO_REG_16__SCAN_IN;
  assign n9267 = ~n9265 & ~n9264;
  assign n9270 = ~n9268 & ~SI_16_;
  assign n10362 = ~n9269 & ~n9270;
  assign n9275 = ~n10415;
  assign n9276 = ~n9274 | ~n9273;
  assign n9277 = ~n9276 | ~SI_17_;
  assign n10439 = ~n9278 | ~n9277;
  assign n9281 = ~n9280 | ~n9279;
  assign n9282 = ~n9281 | ~SI_18_;
  assign n9693 = ~n9285 | ~n9284;
  assign n9292 = ~n12315 & ~n13123;
  assign n9288 = ~n9287 & ~n10417;
  assign n9290 = ~n16322 | ~P1_STATE_REG_SCAN_IN;
  assign n9289 = ~n13309 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n9291 = ~n9290 | ~n9289;
  assign P1_U3336 = n9292 | n9291;
  assign n13037 = ~P2_STATE_REG_SCAN_IN & ~n9365;
  assign n9294 = ~P2_D_REG_4__SCAN_IN & ~P2_D_REG_5__SCAN_IN;
  assign n9293 = ~P2_D_REG_2__SCAN_IN & ~P2_D_REG_3__SCAN_IN;
  assign n9295 = ~n9294 | ~n9293;
  assign n9320 = ~n9295 & ~P2_D_REG_29__SCAN_IN;
  assign n9297 = ~P2_D_REG_12__SCAN_IN & ~P2_D_REG_13__SCAN_IN;
  assign n9296 = ~P2_D_REG_10__SCAN_IN & ~P2_D_REG_11__SCAN_IN;
  assign n9301 = ~n9297 | ~n9296;
  assign n9299 = ~P2_D_REG_8__SCAN_IN & ~P2_D_REG_9__SCAN_IN;
  assign n9298 = ~P2_D_REG_6__SCAN_IN & ~P2_D_REG_7__SCAN_IN;
  assign n9300 = ~n9299 | ~n9298;
  assign n9317 = ~n9301 & ~n9300;
  assign n9303 = ~P2_D_REG_20__SCAN_IN & ~P2_D_REG_21__SCAN_IN;
  assign n9302 = ~P2_D_REG_18__SCAN_IN & ~P2_D_REG_19__SCAN_IN;
  assign n9307 = ~n9303 | ~n9302;
  assign n9305 = ~P2_D_REG_15__SCAN_IN & ~P2_D_REG_17__SCAN_IN;
  assign n9304 = ~P2_D_REG_16__SCAN_IN & ~P2_D_REG_14__SCAN_IN;
  assign n9306 = ~n9305 | ~n9304;
  assign n9315 = ~n9307 & ~n9306;
  assign n9309 = ~P2_D_REG_28__SCAN_IN & ~P2_D_REG_31__SCAN_IN;
  assign n9308 = ~P2_D_REG_26__SCAN_IN & ~P2_D_REG_27__SCAN_IN;
  assign n9313 = ~n9309 | ~n9308;
  assign n9311 = ~P2_D_REG_24__SCAN_IN & ~P2_D_REG_25__SCAN_IN;
  assign n9310 = ~P2_D_REG_22__SCAN_IN & ~P2_D_REG_23__SCAN_IN;
  assign n9312 = ~n9311 | ~n9310;
  assign n9314 = ~n9313 & ~n9312;
  assign n9316 = n9315 & n9314;
  assign n9318 = ~n9317 | ~n9316;
  assign n9319 = ~n9318 & ~P2_D_REG_30__SCAN_IN;
  assign n9321 = n9320 & n9319;
  assign n9330 = ~n9327 | ~n9326;
  assign n11888 = ~n11527 & ~n9331;
  assign n9333 = ~n9332;
  assign n9337 = ~n10247;
  assign n10521 = ~n9337 & ~n9336;
  assign n10540 = ~n10521 | ~n9338;
  assign n9339 = ~n10540 & ~P2_IR_REG_18__SCAN_IN;
  assign n9340 = ~n9343 & ~P2_IR_REG_19__SCAN_IN;
  assign n16798 = ~n16774;
  assign n11539 = ~n14426 | ~n9344;
  assign n9348 = ~n9345 & ~P2_IR_REG_28__SCAN_IN;
  assign n14355 = ~n9348 | ~n9346;
  assign n9359 = n9347 ^ ~P2_IR_REG_30__SCAN_IN;
  assign n9349 = ~n9348 & ~n10520;
  assign n13999 = n9349 ^ ~P2_IR_REG_29__SCAN_IN;
  assign n9358 = ~n13999;
  assign n13434 = ~n14149 & ~n9358;
  assign n9351 = ~n13434 | ~P2_REG2_REG_10__SCAN_IN;
  assign n9350 = ~n13431 | ~P2_REG1_REG_10__SCAN_IN;
  assign n9357 = ~n9600 | ~P2_REG3_REG_10__SCAN_IN;
  assign n10631 = n9359 | n9358;
  assign n9377 = ~n15355 | ~n13325;
  assign n9369 = ~n9380 | ~P2_REG3_REG_12__SCAN_IN;
  assign n9375 = n9371 & n9370;
  assign n9373 = ~n13434 | ~P2_REG2_REG_12__SCAN_IN;
  assign n9372 = ~n13430 | ~P2_REG0_REG_12__SCAN_IN;
  assign n9376 = ~n15604 | ~n16466;
  assign n9378 = ~n9377 | ~n9376;
  assign n9402 = ~n13037 & ~n9378;
  assign n9381 = ~n9379 | ~P2_REG3_REG_11__SCAN_IN;
  assign n11767 = ~n8922 & ~n8925;
  assign n9403 = ~n11767 | ~n16939;
  assign n9650 = ~n16847 & ~n11528;
  assign n11885 = ~n11527 & ~n9389;
  assign n9390 = ~n11888;
  assign n9400 = n9394 | P2_U3151;
  assign n12653 = ~n8922 | ~P2_STATE_REG_SCAN_IN;
  assign n12316 = ~n8926 | ~P2_STATE_REG_SCAN_IN;
  assign n9396 = ~n12653 | ~n12316;
  assign n9397 = n9396 & n16774;
  assign n9401 = ~n13395 | ~n15602;
  assign n9661 = ~n9402 | ~n9401;
  assign n16947 = ~n8922 | ~n16917;
  assign n9404 = ~n9403 | ~n16947;
  assign n9407 = ~n16401 | ~P1_DATAO_REG_1__SCAN_IN;
  assign n9406 = ~n10558 | ~n11356;
  assign n11026 = n9408 ^ SI_1_;
  assign n9409 = ~n11026;
  assign n9410 = ~n10218 & ~n9409;
  assign n9412 = ~n13431 | ~P2_REG1_REG_1__SCAN_IN;
  assign n9415 = ~n8930 | ~P2_REG3_REG_1__SCAN_IN;
  assign n9414 = ~n13434 | ~P2_REG2_REG_1__SCAN_IN;
  assign n9416 = ~n9415 | ~n9414;
  assign n9420 = ~n10558 & ~n9418;
  assign n9419 = ~n14426 & ~n11327;
  assign n11540 = ~n9420 & ~n9419;
  assign n9422 = ~n13430 | ~P2_REG0_REG_0__SCAN_IN;
  assign n9421 = ~n13431 | ~P2_REG1_REG_0__SCAN_IN;
  assign n9426 = ~n9422 | ~n9421;
  assign n9424 = ~n8930 | ~P2_REG3_REG_0__SCAN_IN;
  assign n9423 = ~n13434 | ~P2_REG2_REG_0__SCAN_IN;
  assign n16471 = ~n9426 & ~n9425;
  assign n16470 = ~n11540;
  assign n16472 = ~n16471 | ~n16470;
  assign n12430 = ~n9427 | ~n16472;
  assign n9429 = ~n9428 | ~n16475;
  assign n11971 = ~n9430 | ~n9429;
  assign n9433 = ~n8933 & ~n9431;
  assign n9432 = ~n14426 & ~n11002;
  assign n9435 = ~n9434;
  assign n9455 = ~n9436 | ~n9435;
  assign n9453 = n9437 ^ SI_2_;
  assign n11001 = n9455 ^ n9453;
  assign n12255 = ~n9439 | ~n9438;
  assign n9445 = n9441 & n9440;
  assign n9443 = ~n8930 | ~P2_REG3_REG_2__SCAN_IN;
  assign n9442 = ~n13434 | ~P2_REG2_REG_2__SCAN_IN;
  assign n9444 = n9443 & n9442;
  assign n12421 = ~n9445 | ~n9444;
  assign n11969 = ~n9446 & ~n12421;
  assign n9448 = ~n11971 & ~n11969;
  assign n9447 = ~n9446;
  assign n16495 = ~n12421;
  assign n11970 = ~n9447 & ~n16495;
  assign n12201 = ~n9448 & ~n11970;
  assign n9449 = ~P1_DATAO_REG_3__SCAN_IN;
  assign n9452 = ~n8933 & ~n9449;
  assign n9451 = ~n14426 & ~n9450;
  assign n9462 = ~n9452 & ~n9451;
  assign n9454 = ~n9453;
  assign n9458 = ~n9455 | ~n9454;
  assign n9461 = ~n11044 | ~n8921;
  assign n9465 = ~n8930 | ~n12301;
  assign n9469 = n9465 & n9464;
  assign n9467 = ~n13434 | ~P2_REG2_REG_3__SCAN_IN;
  assign n9466 = ~n13431 | ~P2_REG1_REG_3__SCAN_IN;
  assign n9468 = n9467 & n9466;
  assign n16506 = ~n9469 | ~n9468;
  assign n9470 = ~n12199 | ~n16506;
  assign n9473 = ~n12201 | ~n9470;
  assign n16517 = ~n16506;
  assign n9472 = ~n9471 | ~n16517;
  assign n12458 = ~n9473 | ~n9472;
  assign n9475 = ~n10558 | ~n11570;
  assign n11049 = n9478 ^ n9477;
  assign n9479 = n11049 & n8921;
  assign n16523 = ~n9480 & ~n9479;
  assign n9482 = ~n13430 | ~P2_REG0_REG_4__SCAN_IN;
  assign n9481 = ~n13431 | ~P2_REG1_REG_4__SCAN_IN;
  assign n9487 = ~n9482 | ~n9481;
  assign n9483 = ~P2_REG3_REG_4__SCAN_IN | ~P2_REG3_REG_3__SCAN_IN;
  assign n12659 = ~n9502 | ~n9483;
  assign n9484 = ~n13434 | ~P2_REG2_REG_4__SCAN_IN;
  assign n16522 = ~n9487 & ~n9486;
  assign n9490 = ~n12458 | ~n12459;
  assign n9489 = ~n9488 | ~n16522;
  assign n12186 = ~n9490 | ~n9489;
  assign n9498 = ~n10996 & ~n15584;
  assign n9496 = ~n16401 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n9495 = ~n10558 | ~n11628;
  assign n9500 = ~n13434 | ~P2_REG2_REG_5__SCAN_IN;
  assign n9499 = ~n13431 | ~P2_REG1_REG_5__SCAN_IN;
  assign n9528 = ~n9501;
  assign n9503 = ~n9502 | ~P2_REG3_REG_5__SCAN_IN;
  assign n12790 = ~n9528 | ~n9503;
  assign n9505 = ~n8930 | ~n12790;
  assign n9504 = ~n13430 | ~P2_REG0_REG_5__SCAN_IN;
  assign n12467 = ~n9507 & ~n9506;
  assign n9510 = ~n12186 | ~n12187;
  assign n12673 = ~n9510 | ~n9509;
  assign n9513 = ~n10991;
  assign n9514 = ~P1_DATAO_REG_6__SCAN_IN;
  assign n9525 = ~n8933 & ~n9514;
  assign n9524 = ~n14426 & ~n11872;
  assign n9526 = ~n9525 & ~n9524;
  assign n9529 = ~n9528 | ~P2_REG3_REG_6__SCAN_IN;
  assign n12684 = ~n9529 | ~n9552;
  assign n9531 = ~n8930 | ~n12684;
  assign n9530 = ~n13430 | ~P2_REG0_REG_6__SCAN_IN;
  assign n9533 = ~n13434 | ~P2_REG2_REG_6__SCAN_IN;
  assign n9532 = ~n13431 | ~P2_REG1_REG_6__SCAN_IN;
  assign n9534 = n9533 & n9532;
  assign n9539 = ~n12673 | ~n9536;
  assign n9537 = ~n12671;
  assign n12761 = ~n12769;
  assign n9538 = ~n9537 | ~n12761;
  assign n12548 = ~n9539 | ~n9538;
  assign n9546 = ~n8933 & ~n9542;
  assign n9545 = ~n14426 & ~n12020;
  assign n9547 = ~n9546 & ~n9545;
  assign n9558 = n16551 ^ n15591;
  assign n9550 = ~n13434 | ~P2_REG2_REG_7__SCAN_IN;
  assign n9549 = ~n13430 | ~P2_REG0_REG_7__SCAN_IN;
  assign n9557 = n9550 & n9549;
  assign n9577 = ~n9551;
  assign n9553 = ~n9552 | ~P2_REG3_REG_7__SCAN_IN;
  assign n9555 = ~n8930 | ~n12825;
  assign n9554 = ~n13431 | ~P2_REG1_REG_7__SCAN_IN;
  assign n9556 = n9555 & n9554;
  assign n9560 = ~n9559 | ~n16550;
  assign n9562 = ~n9561;
  assign n9574 = ~n11070 | ~n8921;
  assign n9572 = ~n8933 & ~n9568;
  assign n9571 = ~n14426 & ~n12121;
  assign n9573 = ~n9572 & ~n9571;
  assign n13016 = ~n9574 | ~n9573;
  assign n9576 = ~n13430 | ~P2_REG0_REG_8__SCAN_IN;
  assign n9575 = ~n13431 | ~P2_REG1_REG_8__SCAN_IN;
  assign n9582 = n9576 & n9575;
  assign n9578 = ~n9577 | ~P2_REG3_REG_8__SCAN_IN;
  assign n9580 = ~n8930 | ~n13026;
  assign n9579 = ~n13434 | ~P2_REG2_REG_8__SCAN_IN;
  assign n9585 = ~n13013 & ~n13010;
  assign n9584 = ~n9583;
  assign n12966 = ~n9585 & ~n13011;
  assign n9595 = ~n11114 | ~n8921;
  assign n9588 = ~P1_DATAO_REG_9__SCAN_IN;
  assign n9593 = ~n8933 & ~n9588;
  assign n9613 = ~n9590 & ~n9589;
  assign n9592 = ~n14426 & ~n12536;
  assign n9594 = ~n9593 & ~n9592;
  assign n13315 = ~n9595 | ~n9594;
  assign n9597 = ~n13434 | ~P2_REG2_REG_9__SCAN_IN;
  assign n9596 = ~n13431 | ~P2_REG1_REG_9__SCAN_IN;
  assign n9599 = ~n9598 | ~P2_REG3_REG_9__SCAN_IN;
  assign n9602 = ~n8930 | ~n12981;
  assign n9606 = ~n9605;
  assign n9607 = ~n9606 | ~n13023;
  assign n13406 = ~n12968 & ~n9609;
  assign n9615 = ~n9618 | ~P2_IR_REG_31__SCAN_IN;
  assign n13052 = ~n9620 | ~n9630;
  assign n13041 = ~n13052;
  assign n13230 = ~n9624 & ~n9623;
  assign n9627 = ~n13406 | ~n13407;
  assign n10201 = ~n9627 | ~n9626;
  assign n9637 = ~n13276 & ~n14426;
  assign n9636 = ~n8933 & ~n9635;
  assign n16610 = ~n9639 | ~n9638;
  assign n9643 = ~n13430 | ~P2_REG0_REG_11__SCAN_IN;
  assign n9642 = ~n13434 | ~P2_REG2_REG_11__SCAN_IN;
  assign n9648 = ~n10202 & ~n10200;
  assign n9652 = n9651 & n11883;
  assign n9655 = ~n10958 & ~n16433;
  assign n9658 = ~n16610 | ~n15342;
  assign P2_U3176 = n9661 | n9660;
  assign n9690 = P2_ADDR_REG_19__SCAN_IN ^ n9662;
  assign n13182 = ~P2_ADDR_REG_18__SCAN_IN | ~P1_ADDR_REG_18__SCAN_IN;
  assign n13006 = P2_ADDR_REG_17__SCAN_IN & P1_ADDR_REG_17__SCAN_IN;
  assign n12687 = P2_ADDR_REG_16__SCAN_IN & P1_ADDR_REG_16__SCAN_IN;
  assign n12416 = P2_ADDR_REG_15__SCAN_IN & P1_ADDR_REG_15__SCAN_IN;
  assign n12078 = P2_ADDR_REG_14__SCAN_IN & P1_ADDR_REG_14__SCAN_IN;
  assign n11902 = P2_ADDR_REG_13__SCAN_IN & P1_ADDR_REG_13__SCAN_IN;
  assign n11706 = P2_ADDR_REG_12__SCAN_IN & P1_ADDR_REG_12__SCAN_IN;
  assign n11548 = P2_ADDR_REG_11__SCAN_IN & P1_ADDR_REG_11__SCAN_IN;
  assign n11389 = P2_ADDR_REG_10__SCAN_IN & P1_ADDR_REG_10__SCAN_IN;
  assign n9679 = ~P2_ADDR_REG_9__SCAN_IN & ~P1_ADDR_REG_9__SCAN_IN;
  assign n9677 = ~P2_ADDR_REG_8__SCAN_IN & ~P1_ADDR_REG_8__SCAN_IN;
  assign n9675 = ~P2_ADDR_REG_7__SCAN_IN & ~P1_ADDR_REG_7__SCAN_IN;
  assign n9673 = ~P2_ADDR_REG_6__SCAN_IN | ~P1_ADDR_REG_6__SCAN_IN;
  assign n10967 = P2_ADDR_REG_6__SCAN_IN ^ P1_ADDR_REG_6__SCAN_IN;
  assign n9671 = ~P2_ADDR_REG_5__SCAN_IN & ~P1_ADDR_REG_5__SCAN_IN;
  assign n9669 = ~P2_ADDR_REG_4__SCAN_IN & ~P1_ADDR_REG_4__SCAN_IN;
  assign n9667 = ~P1_ADDR_REG_3__SCAN_IN | ~P2_ADDR_REG_3__SCAN_IN;
  assign n10951 = P1_ADDR_REG_3__SCAN_IN ^ P2_ADDR_REG_3__SCAN_IN;
  assign n9665 = ~P1_ADDR_REG_2__SCAN_IN | ~P2_ADDR_REG_2__SCAN_IN;
  assign n10943 = P1_ADDR_REG_0__SCAN_IN & P2_ADDR_REG_0__SCAN_IN;
  assign n10946 = ~P1_ADDR_REG_1__SCAN_IN & ~n10943;
  assign n10945 = P1_ADDR_REG_1__SCAN_IN & n10943;
  assign n9663 = ~P2_ADDR_REG_1__SCAN_IN & ~n10945;
  assign n10949 = ~n10946 & ~n9663;
  assign n10948 = P1_ADDR_REG_2__SCAN_IN ^ P2_ADDR_REG_2__SCAN_IN;
  assign n9664 = ~n10949 | ~n10948;
  assign n10950 = ~n9665 | ~n9664;
  assign n9666 = ~n10951 | ~n10950;
  assign n10952 = P2_ADDR_REG_4__SCAN_IN ^ ~P1_ADDR_REG_4__SCAN_IN;
  assign n9668 = ~n10953 & ~n10952;
  assign n10954 = P2_ADDR_REG_5__SCAN_IN ^ ~P1_ADDR_REG_5__SCAN_IN;
  assign n9670 = ~n10955 & ~n10954;
  assign n11024 = P2_ADDR_REG_7__SCAN_IN ^ ~P1_ADDR_REG_7__SCAN_IN;
  assign n11076 = P2_ADDR_REG_8__SCAN_IN ^ ~P1_ADDR_REG_8__SCAN_IN;
  assign n11171 = P2_ADDR_REG_9__SCAN_IN ^ ~P1_ADDR_REG_9__SCAN_IN;
  assign n11390 = ~P2_ADDR_REG_10__SCAN_IN & ~P1_ADDR_REG_10__SCAN_IN;
  assign n11549 = ~P2_ADDR_REG_11__SCAN_IN & ~P1_ADDR_REG_11__SCAN_IN;
  assign n11707 = ~P2_ADDR_REG_12__SCAN_IN & ~P1_ADDR_REG_12__SCAN_IN;
  assign n11903 = ~P2_ADDR_REG_13__SCAN_IN & ~P1_ADDR_REG_13__SCAN_IN;
  assign n12079 = ~P2_ADDR_REG_14__SCAN_IN & ~P1_ADDR_REG_14__SCAN_IN;
  assign n12417 = ~P2_ADDR_REG_15__SCAN_IN & ~P1_ADDR_REG_15__SCAN_IN;
  assign n12688 = ~P2_ADDR_REG_16__SCAN_IN & ~P1_ADDR_REG_16__SCAN_IN;
  assign n13007 = ~P2_ADDR_REG_17__SCAN_IN & ~P1_ADDR_REG_17__SCAN_IN;
  assign n13183 = P2_ADDR_REG_18__SCAN_IN | P1_ADDR_REG_18__SCAN_IN;
  assign n9688 = ~n13184 | ~n13183;
  assign n9689 = ~n13182 | ~n9688;
  assign ADD_1068_U4 = n9690 ^ ~n9689;
  assign n9695 = ~n9692 | ~n9691;
  assign n9698 = ~n9697 | ~n9696;
  assign n9701 = ~n8919 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n9703 = ~n9702 | ~n9701;
  assign n9704 = ~n9703 | ~SI_21_;
  assign n9708 = ~n9707 | ~n9706;
  assign n9713 = ~n9712 | ~n9711;
  assign n9714 = ~n9713 | ~SI_23_;
  assign n9716 = ~n8919 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n9718 = ~n9717 | ~n9716;
  assign n9723 = ~n9722 | ~n9721;
  assign n9725 = ~n10677 | ~n10676;
  assign n9730 = ~n9728 & ~n9727;
  assign n10321 = ~n9730 | ~n9729;
  assign n10323 = ~n9734 & ~n9733;
  assign n9740 = ~n9738 | ~P2_STATE_REG_SCAN_IN;
  assign n14356 = ~n10344 | ~P2_U3151;
  assign n9739 = ~n13683 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n9741 = ~n9740 | ~n9739;
  assign P2_U3269 = n9742 | n9741;
  assign n9746 = ~n9744 | ~n9743;
  assign n9745 = ~n10353 & ~n10417;
  assign n9781 = ~n14156 & ~n14005;
  assign n9753 = ~n8923 | ~P1_REG0_REG_0__SCAN_IN;
  assign n9758 = ~n11100 | ~P1_REG2_REG_0__SCAN_IN;
  assign n9757 = ~n8928 | ~P1_REG1_REG_0__SCAN_IN;
  assign n9759 = n9758 & n9757;
  assign n11719 = ~n9760 | ~n9759;
  assign n9762 = ~n9761 | ~P1_IR_REG_31__SCAN_IN;
  assign n11843 = ~n16236 | ~n16324;
  assign n15534 = ~n11910 | ~n16324;
  assign n11840 = ~n15534 & ~n16322;
  assign n9769 = ~n11719 | ~n10906;
  assign n9765 = n10730 & P1_IR_REG_0__SCAN_IN;
  assign n9764 = ~n10730 & ~n9763;
  assign n11922 = ~n9765 & ~n9764;
  assign n9767 = ~n10826 & ~n11922;
  assign n9766 = ~n10133 & ~n11382;
  assign n9768 = ~n9767 & ~n9766;
  assign n11377 = ~n9769 | ~n9768;
  assign n9775 = ~n11377;
  assign n9774 = ~n11719 | ~n9957;
  assign n10901 = ~n9770;
  assign n9772 = ~n10901 | ~n11918;
  assign n9771 = ~n10121 | ~P1_REG1_REG_0__SCAN_IN;
  assign n9773 = n9772 & n9771;
  assign n11378 = ~n9774 | ~n9773;
  assign n9778 = ~n9775 | ~n11378;
  assign n9776 = ~n16149 | ~n8924;
  assign n9777 = ~n9798 | ~n10904;
  assign n9794 = ~n9778 | ~n9777;
  assign n9780 = ~n8923 | ~P1_REG0_REG_1__SCAN_IN;
  assign n9779 = ~n8928 | ~P1_REG1_REG_1__SCAN_IN;
  assign n9785 = ~n9780 | ~n9779;
  assign n9783 = ~n8920 | ~P1_REG3_REG_1__SCAN_IN;
  assign n9782 = ~n11100 | ~P1_REG2_REG_1__SCAN_IN;
  assign n15683 = ~n9785 & ~n9784;
  assign n9792 = ~n15683 & ~n10826;
  assign n9788 = ~n9810 | ~n11026;
  assign n9786 = ~P1_IR_REG_31__SCAN_IN | ~P1_IR_REG_0__SCAN_IN;
  assign n11198 = n9786 ^ ~P1_IR_REG_1__SCAN_IN;
  assign n9787 = ~n10730 | ~n11198;
  assign n9790 = ~n9788 | ~n9787;
  assign n11014 = ~P2_DATAO_REG_1__SCAN_IN;
  assign n9789 = ~n14970 & ~n11014;
  assign n9793 = ~n9792 & ~n9791;
  assign n9797 = n9793 ^ n11662;
  assign n11723 = ~n9794 | ~n9797;
  assign n9796 = ~n15690 | ~n10906;
  assign n15701 = ~n15684;
  assign n9795 = ~n15701 | ~n9957;
  assign n9802 = ~n9797;
  assign n9800 = ~n9798 | ~n11662;
  assign n9799 = ~n11377 | ~n11378;
  assign n11747 = ~n9803 | ~n11722;
  assign n9805 = ~n11100 | ~P1_REG2_REG_2__SCAN_IN;
  assign n9804 = ~n8928 | ~P1_REG1_REG_2__SCAN_IN;
  assign n9809 = n9805 & n9804;
  assign n9808 = n9807 & n9806;
  assign n12496 = ~n9809 | ~n9808;
  assign n9817 = ~n12496 | ~n9957;
  assign n9815 = ~n14967 & ~n11001;
  assign n9834 = ~n9811 | ~P1_IR_REG_31__SCAN_IN;
  assign n11407 = n9834 ^ n9833;
  assign n9812 = ~n10730 | ~n11407;
  assign n12480 = ~n9815 & ~n9814;
  assign n9816 = ~n11812 | ~n10901;
  assign n9818 = ~n9817 | ~n9816;
  assign n9822 = n9818 ^ n10904;
  assign n9820 = ~n12496 | ~n10906;
  assign n9819 = ~n11812 | ~n9957;
  assign n9823 = ~n9820 | ~n9819;
  assign n9825 = ~n11747 | ~n11744;
  assign n9824 = ~n9822;
  assign n12509 = ~n9825 | ~n11745;
  assign n9827 = ~n11100 | ~P1_REG2_REG_3__SCAN_IN;
  assign n9826 = ~n8928 | ~P1_REG1_REG_3__SCAN_IN;
  assign n9828 = ~P1_REG3_REG_3__SCAN_IN;
  assign n9830 = ~n8920 | ~n9828;
  assign n9829 = ~n8923 | ~P1_REG0_REG_3__SCAN_IN;
  assign n9831 = n9830 & n9829;
  assign n15715 = ~n9832 | ~n9831;
  assign n9843 = ~n15715 | ~n9957;
  assign n10842 = ~n14967;
  assign n9835 = ~n9834 | ~n9833;
  assign n9836 = ~n9835 | ~P1_IR_REG_31__SCAN_IN;
  assign n11226 = n9836 ^ P1_IR_REG_3__SCAN_IN;
  assign n9839 = ~n10969 & ~n11226;
  assign n9837 = ~P2_DATAO_REG_3__SCAN_IN;
  assign n9838 = ~n14970 & ~n9837;
  assign n9840 = ~n9839 & ~n9838;
  assign n15714 = ~n9841 | ~n9840;
  assign n9842 = ~n15714 | ~n10901;
  assign n9844 = ~n9843 | ~n9842;
  assign n9848 = n9844 ^ n10904;
  assign n9846 = ~n15715 | ~n10906;
  assign n9845 = ~n15714 | ~n9957;
  assign n9849 = ~n9846 | ~n9845;
  assign n9847 = ~n9849;
  assign n12506 = ~n9848 & ~n9847;
  assign n9851 = ~n12509 & ~n12506;
  assign n9850 = ~n9848;
  assign n12507 = ~n9850 & ~n9849;
  assign n12085 = ~n9851 & ~n12507;
  assign n9853 = ~n11100 | ~P1_REG2_REG_4__SCAN_IN;
  assign n9854 = ~P1_REG3_REG_4__SCAN_IN & ~P1_REG3_REG_3__SCAN_IN;
  assign n12084 = ~n9898 & ~n9854;
  assign n9856 = ~n8920 | ~n12084;
  assign n9855 = ~n8923 | ~P1_REG0_REG_4__SCAN_IN;
  assign n9857 = n9856 & n9855;
  assign n15722 = ~n9858 | ~n9857;
  assign n9868 = ~n15722 | ~n9957;
  assign n9866 = ~n11049 | ~n10842;
  assign n9861 = ~n9859 & ~n10417;
  assign n11203 = n9861 ^ n9860;
  assign n9864 = ~n10969 & ~n11203;
  assign n9862 = ~P2_DATAO_REG_4__SCAN_IN;
  assign n9863 = ~n14970 & ~n9862;
  assign n9865 = ~n9864 & ~n9863;
  assign n15723 = ~n9866 | ~n9865;
  assign n9867 = ~n15723 | ~n10901;
  assign n9869 = ~n9868 | ~n9867;
  assign n9873 = n9869 ^ n11662;
  assign n9871 = ~n15722 | ~n10906;
  assign n9870 = ~n15723 | ~n9957;
  assign n9875 = ~n12085 | ~n12086;
  assign n12324 = ~n9875 | ~n9874;
  assign n9879 = ~n10996 & ~n14967;
  assign n9877 = ~n10864 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n9876 = ~n10730 | ~n11473;
  assign n9878 = ~n9877 | ~n9876;
  assign n12349 = ~n9879 & ~n9878;
  assign n9888 = ~n15738 | ~n10901;
  assign n9881 = ~n11100 | ~P1_REG2_REG_5__SCAN_IN;
  assign n9880 = ~n8923 | ~P1_REG0_REG_5__SCAN_IN;
  assign n9886 = n9881 & n9880;
  assign n12707 = n9882 ^ ~P1_REG3_REG_5__SCAN_IN;
  assign n9884 = ~n8920 | ~n12707;
  assign n9883 = ~n8928 | ~P1_REG1_REG_5__SCAN_IN;
  assign n15739 = ~n9886 | ~n9885;
  assign n9887 = ~n15739 | ~n9957;
  assign n9891 = ~n12217 & ~n10827;
  assign n9890 = ~n12349 & ~n10826;
  assign n9892 = ~n12322 & ~n12435;
  assign n9912 = ~n12324 & ~n9892;
  assign n9897 = ~n10991 & ~n14967;
  assign n9895 = ~n10864 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n9894 = ~n10730 | ~n11251;
  assign n12371 = ~n9897 & ~n9896;
  assign n9906 = ~n12371 & ~n9770;
  assign n12449 = n9925 ^ ~P1_REG3_REG_6__SCAN_IN;
  assign n9900 = ~n8920 | ~n12449;
  assign n9899 = ~n11100 | ~P1_REG2_REG_6__SCAN_IN;
  assign n9904 = n9900 & n9899;
  assign n9902 = ~n8923 | ~P1_REG0_REG_6__SCAN_IN;
  assign n9901 = ~n8928 | ~P1_REG1_REG_6__SCAN_IN;
  assign n9903 = n9902 & n9901;
  assign n9905 = ~n12847 & ~n10826;
  assign n9907 = ~n9906 & ~n9905;
  assign n9909 = ~n12371 & ~n10826;
  assign n9908 = ~n12847 & ~n10827;
  assign n9910 = ~n12322 | ~n12435;
  assign n9918 = ~n9916;
  assign n9917 = ~P1_IR_REG_6__SCAN_IN;
  assign n9922 = ~n10969 & ~n11492;
  assign n11019 = ~P2_DATAO_REG_7__SCAN_IN;
  assign n9921 = ~n14970 & ~n11019;
  assign n15750 = ~n9924 | ~n9923;
  assign n12850 = n9950 ^ P1_REG3_REG_7__SCAN_IN;
  assign n9927 = ~n8920 | ~n12850;
  assign n9926 = ~n8923 | ~P1_REG0_REG_7__SCAN_IN;
  assign n9931 = n9927 & n9926;
  assign n9929 = ~n11100 | ~P1_REG2_REG_7__SCAN_IN;
  assign n9928 = ~n8928 | ~P1_REG1_REG_7__SCAN_IN;
  assign n9930 = n9929 & n9928;
  assign n9936 = ~n15750 | ~n9957;
  assign n9935 = ~n15751 | ~n10906;
  assign n9941 = ~n12839 | ~n12836;
  assign n9963 = ~n9941 | ~n12837;
  assign n9942 = ~P1_IR_REG_6__SCAN_IN & ~P1_IR_REG_7__SCAN_IN;
  assign n11055 = ~n11282;
  assign n9947 = ~n10969 & ~n11055;
  assign n9946 = ~n14970 & ~n11054;
  assign n9948 = ~n9947 & ~n9946;
  assign n12879 = n9975 ^ ~P1_REG3_REG_8__SCAN_IN;
  assign n9952 = ~n8920 | ~n12879;
  assign n9951 = ~n8928 | ~P1_REG1_REG_8__SCAN_IN;
  assign n9956 = n9952 & n9951;
  assign n9954 = ~n11100 | ~P1_REG2_REG_8__SCAN_IN;
  assign n9953 = ~n8923 | ~P1_REG0_REG_8__SCAN_IN;
  assign n9955 = n9954 & n9953;
  assign n9958 = ~n15773 | ~n9957;
  assign n12870 = ~n9963 | ~n9964;
  assign n9962 = ~n15772 | ~n10907;
  assign n9961 = ~n15773 | ~n10906;
  assign n9967 = ~n12870 | ~n12872;
  assign n12871 = ~n9966 | ~n9965;
  assign n12857 = ~n9967 | ~n12871;
  assign n9974 = ~n11114 | ~n10842;
  assign n9972 = ~n10969 & ~n11211;
  assign n9970 = ~P2_DATAO_REG_9__SCAN_IN;
  assign n9971 = ~n14970 & ~n9970;
  assign n15788 = ~n9974 | ~n9973;
  assign n9983 = ~n15788 | ~n10901;
  assign n12920 = n10002 ^ P1_REG3_REG_9__SCAN_IN;
  assign n9977 = ~n8920 | ~n12920;
  assign n9976 = ~n8928 | ~P1_REG1_REG_9__SCAN_IN;
  assign n9981 = n9977 & n9976;
  assign n9979 = ~n11100 | ~P1_REG2_REG_9__SCAN_IN;
  assign n9978 = ~n8923 | ~P1_REG0_REG_9__SCAN_IN;
  assign n9980 = n9979 & n9978;
  assign n9985 = ~n15789 | ~n10906;
  assign n9994 = ~n12857 & ~n12858;
  assign n15802 = ~n10001 & ~n10000;
  assign n13298 = n10032 ^ ~P1_REG3_REG_10__SCAN_IN;
  assign n10004 = ~n8920 | ~n13298;
  assign n10003 = ~n8923 | ~P1_REG0_REG_10__SCAN_IN;
  assign n10007 = ~n11100 | ~P1_REG2_REG_10__SCAN_IN;
  assign n10006 = ~n8928 | ~P1_REG1_REG_10__SCAN_IN;
  assign n10010 = ~n15803 & ~n10826;
  assign n13288 = ~n10015 | ~n10016;
  assign n10014 = ~n15802 & ~n10826;
  assign n10013 = ~n15803 & ~n10827;
  assign n10019 = ~n13288 | ~n13290;
  assign n10018 = ~n10015;
  assign n13289 = ~n10018 | ~n10017;
  assign n10023 = ~P1_IR_REG_11__SCAN_IN;
  assign n11497 = ~n11609;
  assign n10027 = ~n11497 & ~n10969;
  assign n10026 = ~n14970 & ~n10025;
  assign n13517 = ~n10029 | ~n10028;
  assign n10031 = ~n11100 | ~P1_REG2_REG_11__SCAN_IN;
  assign n10030 = ~n8928 | ~P1_REG1_REG_11__SCAN_IN;
  assign n10034 = ~n10035;
  assign n10033 = ~P1_REG3_REG_11__SCAN_IN;
  assign n10036 = ~n10034 | ~n10033;
  assign n13501 = ~n10036 | ~n10150;
  assign n10037 = ~n13501;
  assign n10039 = ~n8920 | ~n10037;
  assign n10038 = ~n8923 | ~P1_REG0_REG_11__SCAN_IN;
  assign n10051 = ~n13511 & ~n10047;
  assign n10262 = ~n10051 & ~n10050;
  assign n10054 = ~n10053;
  assign n11435 = ~n10057 | ~n10056;
  assign n10060 = ~n10969 & ~n11600;
  assign n10059 = ~n14970 & ~n11267;
  assign n15819 = ~n10062 | ~n10061;
  assign n10070 = ~n15819 | ~n10901;
  assign n13060 = n10150 ^ ~P1_REG3_REG_12__SCAN_IN;
  assign n10064 = ~n8920 | ~n13060;
  assign n10063 = ~n8928 | ~P1_REG1_REG_12__SCAN_IN;
  assign n10068 = n10064 & n10063;
  assign n10066 = ~n11100 | ~P1_REG2_REG_12__SCAN_IN;
  assign n10065 = ~n8923 | ~P1_REG0_REG_12__SCAN_IN;
  assign n10067 = n10066 & n10065;
  assign n10073 = ~n15819 | ~n10907;
  assign n10072 = ~n15820 | ~n10906;
  assign n10078 = ~n10263 | ~n10261;
  assign n10080 = ~P1_D_REG_4__SCAN_IN & ~P1_D_REG_5__SCAN_IN;
  assign n10079 = ~P1_D_REG_2__SCAN_IN & ~P1_D_REG_3__SCAN_IN;
  assign n10081 = ~n10080 | ~n10079;
  assign n10106 = ~n10081 & ~P1_D_REG_29__SCAN_IN;
  assign n10083 = ~P1_D_REG_12__SCAN_IN & ~P1_D_REG_13__SCAN_IN;
  assign n10082 = ~P1_D_REG_10__SCAN_IN & ~P1_D_REG_11__SCAN_IN;
  assign n10087 = ~n10083 | ~n10082;
  assign n10085 = ~P1_D_REG_8__SCAN_IN & ~P1_D_REG_9__SCAN_IN;
  assign n10084 = ~P1_D_REG_6__SCAN_IN & ~P1_D_REG_7__SCAN_IN;
  assign n10086 = ~n10085 | ~n10084;
  assign n10103 = ~n10087 & ~n10086;
  assign n10089 = ~P1_D_REG_20__SCAN_IN & ~P1_D_REG_21__SCAN_IN;
  assign n10088 = ~P1_D_REG_18__SCAN_IN & ~P1_D_REG_19__SCAN_IN;
  assign n10093 = ~n10089 | ~n10088;
  assign n10091 = ~P1_D_REG_15__SCAN_IN & ~P1_D_REG_17__SCAN_IN;
  assign n10090 = ~P1_D_REG_16__SCAN_IN & ~P1_D_REG_14__SCAN_IN;
  assign n10092 = ~n10091 | ~n10090;
  assign n10101 = ~n10093 & ~n10092;
  assign n10095 = ~P1_D_REG_28__SCAN_IN & ~P1_D_REG_31__SCAN_IN;
  assign n10094 = ~P1_D_REG_26__SCAN_IN & ~P1_D_REG_27__SCAN_IN;
  assign n10099 = ~n10095 | ~n10094;
  assign n10097 = ~P1_D_REG_24__SCAN_IN & ~P1_D_REG_25__SCAN_IN;
  assign n10096 = ~P1_D_REG_22__SCAN_IN & ~P1_D_REG_23__SCAN_IN;
  assign n10098 = ~n10097 | ~n10096;
  assign n10100 = ~n10099 & ~n10098;
  assign n10102 = n10101 & n10100;
  assign n10104 = ~n10103 | ~n10102;
  assign n10105 = ~n10104 & ~P1_D_REG_30__SCAN_IN;
  assign n10113 = ~n10106 | ~n10105;
  assign n10108 = ~P1_B_REG_SCAN_IN;
  assign n10109 = ~n13165 | ~n10108;
  assign n10117 = ~n13165;
  assign n13221 = ~n11910 | ~n16224;
  assign n10122 = ~n11910 | ~n16322;
  assign n16369 = ~n13221 | ~n10122;
  assign n10129 = ~n10144;
  assign n10125 = ~n13221;
  assign n10140 = ~n11658 | ~n10125;
  assign n10127 = ~n10126 | ~n8924;
  assign n16332 = ~n16149;
  assign n11911 = ~n10127 & ~n16332;
  assign n10128 = ~n10140 | ~n16331;
  assign n10130 = ~n16324 | ~n8924;
  assign n10132 = ~n10144 & ~n10131;
  assign n10968 = ~n10135;
  assign n10138 = ~n13060 | ~n15516;
  assign n11654 = ~n15534 & ~n8924;
  assign n10162 = ~n15819 | ~n15428;
  assign n10143 = ~n16331;
  assign n10145 = ~n15094 & ~n13283;
  assign n11603 = ~P1_STATE_REG_SCAN_IN & ~n10149;
  assign n10160 = n10145 | n11603;
  assign n13881 = ~n11686;
  assign n15515 = ~n10146 | ~n13881;
  assign n10153 = ~n10151;
  assign n10152 = ~P1_REG3_REG_13__SCAN_IN;
  assign n10154 = ~n10153 | ~n10152;
  assign n10159 = ~n15515 & ~n15840;
  assign n10161 = ~n10160 & ~n10159;
  assign n10163 = ~n10162 | ~n10161;
  assign P1_U3224 = n10164 | n10163;
  assign n14583 = ~P2_STATE_REG_SCAN_IN & ~n10166;
  assign n10184 = ~n10228 & ~P2_REG3_REG_14__SCAN_IN;
  assign n10168 = ~n13430 | ~P2_REG0_REG_16__SCAN_IN;
  assign n10167 = ~n13431 | ~P2_REG1_REG_16__SCAN_IN;
  assign n13973 = ~P2_REG2_REG_16__SCAN_IN;
  assign n10182 = ~n14079 | ~n15604;
  assign n10176 = ~n10184;
  assign n10175 = ~n10228 | ~P2_REG3_REG_14__SCAN_IN;
  assign n13869 = ~n10176 | ~n10175;
  assign n10178 = ~n8930 | ~n13869;
  assign n10181 = ~n15355 | ~n16631;
  assign n10183 = ~n10182 | ~n10181;
  assign n10186 = ~n14583 & ~n10183;
  assign n10185 = ~n13746 | ~n15602;
  assign n10260 = ~n10186 | ~n10185;
  assign n10510 = ~n10247 & ~n10520;
  assign n16637 = ~n10193 & ~n10192;
  assign n10507 = n16637 ^ n15591;
  assign n10195 = ~n13746 | ~n8930;
  assign n10203 = ~n10201 & ~n10200;
  assign n13635 = ~n10210 | ~n10209;
  assign n10221 = ~n10219 | ~P2_IR_REG_31__SCAN_IN;
  assign n10220 = ~P2_IR_REG_13__SCAN_IN;
  assign n16461 = ~n10225 & ~n10224;
  assign n10227 = ~n10226 | ~P2_REG3_REG_13__SCAN_IN;
  assign n13653 = ~n10228 | ~n10227;
  assign n10230 = ~n8930 | ~n13653;
  assign n10234 = n10230 & n10229;
  assign n10232 = ~n13434 | ~P2_REG2_REG_13__SCAN_IN;
  assign n10235 = ~n13466 | ~n13859;
  assign n10238 = ~n13468 | ~n10235;
  assign n13594 = ~n10238 | ~n10237;
  assign n10242 = ~P1_DATAO_REG_14__SCAN_IN;
  assign n10250 = ~n8933 & ~n10242;
  assign n10244 = ~n9332 & ~n10520;
  assign n10243 = ~P2_IR_REG_14__SCAN_IN;
  assign n10246 = ~n10244 & ~n10243;
  assign n10245 = ~n10520 & ~P2_IR_REG_14__SCAN_IN;
  assign n10248 = ~n10246 & ~n10245;
  assign n14587 = ~n10248 & ~n10247;
  assign n10249 = ~n14426 & ~n14598;
  assign n16628 = ~n10252 | ~n10251;
  assign n10255 = ~n13594 | ~n13595;
  assign n10506 = ~n10255 | ~n10254;
  assign P2_U3181 = n10260 | n10259;
  assign n10264 = ~n10262 | ~n10261;
  assign n13524 = ~n10264 | ~n10263;
  assign n10368 = ~n10265 & ~P1_IR_REG_12__SCAN_IN;
  assign n10266 = ~n10368 & ~n10417;
  assign n15839 = ~n10270 & ~n10269;
  assign n10271 = ~n15840 & ~n10826;
  assign n10365 = ~P1_IR_REG_13__SCAN_IN;
  assign n10281 = ~n10368 | ~n10365;
  assign n10284 = ~n10969 & ~n12564;
  assign n10283 = ~n14970 & ~n10282;
  assign n15849 = ~n10286 | ~n10285;
  assign n13536 = n10375 ^ ~P1_REG3_REG_14__SCAN_IN;
  assign n10288 = ~n8920 | ~n13536;
  assign n10287 = ~n8923 | ~P1_REG0_REG_14__SCAN_IN;
  assign n10292 = n10288 & n10287;
  assign n10290 = ~n11100 | ~P1_REG2_REG_14__SCAN_IN;
  assign n10289 = ~n8928 | ~P1_REG1_REG_14__SCAN_IN;
  assign n10360 = ~n10297 | ~n10296;
  assign n10359 = ~n10299 | ~n10298;
  assign n10302 = ~n10360 | ~n10359;
  assign n10300 = ~n15850 | ~n10906;
  assign n10318 = ~n15516 | ~n13536;
  assign n10316 = ~n13604 & ~n15518;
  assign n10304 = ~n15094 & ~n15840;
  assign n10305 = ~P1_REG3_REG_14__SCAN_IN;
  assign n12565 = ~P1_STATE_REG_SCAN_IN & ~n10305;
  assign n10314 = ~n10304 & ~n12565;
  assign n10306 = ~n10375 & ~n10305;
  assign n14112 = n10306 ^ P1_REG3_REG_15__SCAN_IN;
  assign n10308 = ~n14112 | ~n8920;
  assign n10307 = ~n8923 | ~P1_REG0_REG_15__SCAN_IN;
  assign n10312 = n10308 & n10307;
  assign n10310 = ~n11100 | ~P1_REG2_REG_15__SCAN_IN;
  assign n10309 = ~n8928 | ~P1_REG1_REG_15__SCAN_IN;
  assign n10313 = ~n15439 | ~n14136;
  assign n10315 = ~n10314 | ~n10313;
  assign n10317 = ~n10316 & ~n10315;
  assign n10319 = ~n10318 | ~n10317;
  assign P1_U3215 = n10320 | n10319;
  assign n10326 = ~n10325 | ~n10324;
  assign n10328 = ~n10692 | ~n10690;
  assign n10331 = ~n10330 | ~n10329;
  assign n10333 = ~n10898 | ~n10897;
  assign n10335 = ~n10344 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n10334 = ~n8919 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n10338 = ~n13998 | ~n13997;
  assign n10340 = ~n10344 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n10339 = ~n10345 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n10343 = ~n14148 | ~n14147;
  assign n10347 = ~n10344 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n10346 = ~n10345 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n10348 = ~n10347 | ~n10346;
  assign n10351 = ~P1_IR_REG_31__SCAN_IN | ~P1_STATE_REG_SCAN_IN;
  assign n10352 = ~n10351 & ~P1_IR_REG_30__SCAN_IN;
  assign n10355 = ~n10353 | ~n10352;
  assign n10354 = ~n13309 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n10356 = ~n10355 | ~n10354;
  assign P1_U3324 = n10357 | n10356;
  assign n10361 = ~n10359 | ~n10358;
  assign n14109 = ~n10361 | ~n10360;
  assign n10366 = ~n10365 | ~n10387;
  assign n10367 = ~n10366 & ~P1_IR_REG_15__SCAN_IN;
  assign n10369 = ~n10416 | ~P1_IR_REG_31__SCAN_IN;
  assign n10370 = ~n10730 | ~n14457;
  assign n13797 = ~n10373 & ~n10372;
  assign n14134 = n10425 ^ P1_REG3_REG_16__SCAN_IN;
  assign n10377 = ~n14134 | ~n8920;
  assign n10376 = ~n8923 | ~P1_REG0_REG_16__SCAN_IN;
  assign n10381 = n10377 & n10376;
  assign n10379 = ~n11100 | ~P1_REG2_REG_16__SCAN_IN;
  assign n10378 = ~n8928 | ~P1_REG1_REG_16__SCAN_IN;
  assign n10380 = n10379 & n10378;
  assign n10382 = ~n14116 & ~n10826;
  assign n10385 = ~n14060 | ~n10906;
  assign n10389 = ~n10388 | ~n10387;
  assign n10391 = ~n10730 | ~n13840;
  assign n13619 = ~n10394 & ~n10393;
  assign n10395 = ~n13694 & ~n10826;
  assign n10398 = ~n14136 | ~n10906;
  assign n10413 = ~n14109 | ~n10402;
  assign n14055 = ~n10413 | ~n10412;
  assign n10443 = ~n10416 & ~P1_IR_REG_16__SCAN_IN;
  assign n10418 = ~n10443 & ~n10417;
  assign n15888 = ~n10422 & ~n10421;
  assign n10424 = ~n11100 | ~P1_REG2_REG_17__SCAN_IN;
  assign n10423 = ~n8928 | ~P1_REG1_REG_17__SCAN_IN;
  assign n10426 = ~n8923 | ~P1_REG0_REG_17__SCAN_IN;
  assign n10430 = ~n15885 & ~n10826;
  assign n10438 = ~n14055 | ~n14056;
  assign n10465 = ~n10438 | ~n10437;
  assign n10463 = ~n10465;
  assign n10442 = ~P1_IR_REG_17__SCAN_IN;
  assign n10444 = ~n10443 | ~n10442;
  assign n10446 = ~n10444 | ~P1_IR_REG_31__SCAN_IN;
  assign n10449 = ~n10969 & ~n14754;
  assign n10447 = ~P2_DATAO_REG_18__SCAN_IN;
  assign n10448 = ~n14970 & ~n10447;
  assign n15880 = ~n10451 | ~n10450;
  assign n10456 = ~n11100 | ~P1_REG2_REG_18__SCAN_IN;
  assign n10455 = ~n8923 | ~P1_REG0_REG_18__SCAN_IN;
  assign n10728 = ~n10463 | ~n10462;
  assign n10468 = ~n10728 | ~n10727;
  assign n10466 = ~n15883 | ~n10906;
  assign n10485 = ~n15516 | ~n13819;
  assign n10483 = ~n14178 & ~n15518;
  assign n10477 = ~n14439 | ~n8920;
  assign n10472 = ~n11100 | ~P1_REG2_REG_19__SCAN_IN;
  assign n10471 = ~n8923 | ~P1_REG0_REG_19__SCAN_IN;
  assign n10473 = ~P1_REG1_REG_19__SCAN_IN;
  assign n10474 = ~n8927 & ~n10473;
  assign n10481 = ~n15901 | ~n15439;
  assign n10479 = ~n15094 & ~n15885;
  assign n14762 = ~P1_STATE_REG_SCAN_IN & ~n10478;
  assign n10480 = ~n10479 & ~n14762;
  assign n10482 = ~n10481 | ~n10480;
  assign P1_U3238 = n10487 | n10486;
  assign n10563 = ~P2_REG3_REG_18__SCAN_IN & ~n10546;
  assign n10581 = ~n10563 | ~n10489;
  assign n10491 = ~n8930 | ~n15460;
  assign n10493 = ~n13434 | ~P2_REG2_REG_26__SCAN_IN;
  assign n10492 = ~n13430 | ~P2_REG0_REG_26__SCAN_IN;
  assign n10494 = n10493 & n10492;
  assign n10504 = ~n15355 | ~n15572;
  assign n10497 = ~n13430 | ~P2_REG0_REG_28__SCAN_IN;
  assign n10496 = ~n13431 | ~P2_REG1_REG_28__SCAN_IN;
  assign n10502 = n10497 & n10496;
  assign n10697 = P2_REG3_REG_26__SCAN_IN | n10498;
  assign n13400 = n10697 | P2_REG3_REG_27__SCAN_IN;
  assign n10500 = ~n8930 | ~n16357;
  assign n10499 = ~n13434 | ~P2_REG2_REG_28__SCAN_IN;
  assign n15589 = ~n10502 | ~n10501;
  assign n10509 = ~n10506 | ~n10505;
  assign n10516 = ~n11804 & ~n15584;
  assign n10511 = ~n10510 & ~P2_IR_REG_15__SCAN_IN;
  assign n10512 = ~n10511 & ~n10520;
  assign n14075 = ~n10516 & ~n10515;
  assign n10519 = ~n13900 & ~n13898;
  assign n14043 = ~n10519 & ~n13897;
  assign n10522 = ~n10521 & ~n10520;
  assign n16658 = ~n10526 & ~n10525;
  assign n10529 = ~n13434 | ~P2_REG2_REG_17__SCAN_IN;
  assign n10528 = ~n13430 | ~P2_REG0_REG_17__SCAN_IN;
  assign n10531 = ~n10671 & ~n10530;
  assign n10539 = ~P1_DATAO_REG_18__SCAN_IN;
  assign n10543 = ~n8933 & ~n10539;
  assign n10542 = ~n14426 & ~n15381;
  assign n16679 = ~n10545 | ~n10544;
  assign n10548 = ~n13430 | ~P2_REG0_REG_18__SCAN_IN;
  assign n10547 = ~n13431 | ~P2_REG1_REG_18__SCAN_IN;
  assign n14296 = ~P2_REG2_REG_18__SCAN_IN;
  assign n16680 = ~n10553 | ~n10552;
  assign n10557 = ~n14164 | ~n10554;
  assign n14323 = ~n10557 | ~n10556;
  assign n16695 = ~n10562 & ~n10561;
  assign n10570 = ~n14381 | ~n8930;
  assign n10565 = ~n13434 | ~P2_REG2_REG_19__SCAN_IN;
  assign n10564 = ~n13431 | ~P2_REG1_REG_19__SCAN_IN;
  assign n10566 = ~P2_REG0_REG_19__SCAN_IN;
  assign n10567 = ~n10631 & ~n10566;
  assign n14492 = ~n10570 | ~n10569;
  assign n10574 = ~n14323 | ~n10571;
  assign n14475 = ~n10574 | ~n10573;
  assign n12490 = n10577 ^ n10576;
  assign n10578 = ~P1_DATAO_REG_20__SCAN_IN;
  assign n10588 = ~n14507 | ~n8930;
  assign n10583 = ~n13434 | ~P2_REG2_REG_20__SCAN_IN;
  assign n10582 = ~n13430 | ~P2_REG0_REG_20__SCAN_IN;
  assign n10584 = ~P2_REG1_REG_20__SCAN_IN;
  assign n10591 = ~n14475 & ~n14473;
  assign n10594 = ~P1_DATAO_REG_21__SCAN_IN;
  assign n10597 = ~P2_REG3_REG_21__SCAN_IN;
  assign n10605 = ~n14652 | ~n8930;
  assign n10600 = ~n13431 | ~P2_REG1_REG_21__SCAN_IN;
  assign n10599 = ~n13434 | ~P2_REG2_REG_21__SCAN_IN;
  assign n10601 = ~P2_REG0_REG_21__SCAN_IN;
  assign n10602 = ~n10631 & ~n10601;
  assign n16724 = ~n10605 | ~n10604;
  assign n10609 = ~n14624 | ~n10606;
  assign n10612 = ~P1_DATAO_REG_22__SCAN_IN;
  assign n10616 = ~n13434 | ~P2_REG2_REG_22__SCAN_IN;
  assign n10615 = ~n13430 | ~P2_REG0_REG_22__SCAN_IN;
  assign n10621 = n10616 & n10615;
  assign n10619 = ~n8930 | ~n14808;
  assign n10626 = ~n14804 & ~n16734;
  assign n10625 = ~n10624 & ~n10623;
  assign n15330 = ~n10626 & ~n10625;
  assign n10635 = ~n15341 | ~n8930;
  assign n10629 = ~n13431 | ~P2_REG1_REG_24__SCAN_IN;
  assign n10628 = ~n13434 | ~P2_REG2_REG_24__SCAN_IN;
  assign n10630 = ~P2_REG0_REG_24__SCAN_IN;
  assign n10632 = ~n10631 & ~n10630;
  assign n15343 = ~n10640 | ~n10639;
  assign n10643 = ~P1_DATAO_REG_23__SCAN_IN;
  assign n10654 = ~n15218 | ~n8930;
  assign n10649 = ~n13434 | ~P2_REG2_REG_23__SCAN_IN;
  assign n10648 = ~n13430 | ~P2_REG0_REG_23__SCAN_IN;
  assign n10651 = ~n10671 & ~n10650;
  assign n10665 = ~n15330 & ~n10657;
  assign n10666 = ~P2_REG3_REG_25__SCAN_IN;
  assign n10675 = ~n15239 | ~n8930;
  assign n10669 = ~n13430 | ~P2_REG0_REG_25__SCAN_IN;
  assign n10668 = ~n13434 | ~P2_REG2_REG_25__SCAN_IN;
  assign n10670 = ~P2_REG1_REG_25__SCAN_IN;
  assign n10672 = ~n10671 & ~n10670;
  assign n10683 = ~n15142 & ~n15141;
  assign n15353 = ~n10683 & ~n10682;
  assign n10685 = ~n13459 | ~n8921;
  assign n10689 = ~n15353 & ~n15352;
  assign n10694 = ~n13672 | ~n8921;
  assign n16778 = ~n10694 | ~n10693;
  assign n10696 = ~n13430 | ~P2_REG0_REG_27__SCAN_IN;
  assign n10695 = ~n13431 | ~P2_REG1_REG_27__SCAN_IN;
  assign n10701 = n10696 & n10695;
  assign n10699 = ~n8930 | ~n15565;
  assign n10702 = n15583 ^ ~n15582;
  assign n10708 = ~n10702 | ~n15596;
  assign n10704 = ~n15602 | ~n15565;
  assign n10703 = ~P2_U3151 | ~P2_REG3_REG_27__SCAN_IN;
  assign n10709 = ~n10708 | ~n10707;
  assign P2_U3154 = n10710 | n10709;
  assign n10886 = ~P1_REG3_REG_27__SCAN_IN;
  assign n10713 = ~n8923 | ~P1_REG0_REG_27__SCAN_IN;
  assign n10712 = ~n8928 | ~P1_REG1_REG_27__SCAN_IN;
  assign n15322 = ~P1_REG2_REG_27__SCAN_IN;
  assign n10715 = ~n10714 & ~n15322;
  assign n10717 = ~n10716 & ~n10715;
  assign n10720 = ~n13680 & ~n14967;
  assign n13674 = ~P2_DATAO_REG_27__SCAN_IN;
  assign n14437 = ~n10729 | ~n10728;
  assign n10731 = ~n10730 | ~n16322;
  assign n15902 = ~n10734 & ~n10733;
  assign n10735 = ~n14610 & ~n10826;
  assign n12491 = ~P2_DATAO_REG_20__SCAN_IN;
  assign n10754 = ~n14609 | ~n8920;
  assign n10749 = ~n11100 | ~P1_REG2_REG_20__SCAN_IN;
  assign n10748 = ~n8928 | ~P1_REG1_REG_20__SCAN_IN;
  assign n10750 = ~P1_REG0_REG_20__SCAN_IN;
  assign n10751 = ~n10926 & ~n10750;
  assign n10753 = ~n10752 & ~n10751;
  assign n10755 = ~n14737 & ~n10826;
  assign n10760 = ~n14970 & ~n12733;
  assign n14400 = ~n10761 & ~n10760;
  assign n10763 = ~n11100 | ~P1_REG2_REG_21__SCAN_IN;
  assign n10766 = ~n8920 | ~n14735;
  assign n10769 = ~n14914 & ~n10826;
  assign n10780 = ~n10777 & ~n10776;
  assign n12883 = ~P2_DATAO_REG_22__SCAN_IN;
  assign n10784 = ~n11100 | ~P1_REG2_REG_22__SCAN_IN;
  assign n10787 = ~n8920 | ~n14919;
  assign n10790 = ~n15937 & ~n10826;
  assign n14908 = ~n10795 | ~n10796;
  assign n10794 = ~n15936 & ~n10826;
  assign n10793 = ~n15937 & ~n10827;
  assign n10799 = ~n14908 | ~n14909;
  assign n10798 = ~n10795;
  assign n14907 = ~n10798 | ~n10797;
  assign n10803 = ~n11100 | ~P1_REG2_REG_24__SCAN_IN;
  assign n10802 = ~n8928 | ~P1_REG1_REG_24__SCAN_IN;
  assign n13125 = ~P2_DATAO_REG_23__SCAN_IN;
  assign n10817 = ~n11100 | ~P1_REG2_REG_23__SCAN_IN;
  assign n10816 = ~n8928 | ~P1_REG1_REG_23__SCAN_IN;
  assign n10820 = ~n8920 | ~n15091;
  assign n15949 = ~n10822 | ~n10821;
  assign n10823 = ~n15953 & ~n10826;
  assign n10829 = ~n15952 & ~n10826;
  assign n15038 = ~n10841 | ~n10840;
  assign n10846 = ~n11100 | ~P1_REG2_REG_25__SCAN_IN;
  assign n15983 = ~n10851 & ~n10850;
  assign n15039 = ~n15038 | ~n15037;
  assign n15425 = ~n15039 | ~n10863;
  assign n10868 = ~n11100 | ~P1_REG2_REG_26__SCAN_IN;
  assign n10867 = ~n8928 | ~P1_REG1_REG_26__SCAN_IN;
  assign n10873 = n10868 & n10867;
  assign n10870 = ~n8923 | ~P1_REG0_REG_26__SCAN_IN;
  assign n10884 = ~n15425 | ~n15424;
  assign n10885 = ~n15513;
  assign n10891 = ~n11100 | ~P1_REG2_REG_28__SCAN_IN;
  assign n10890 = ~n8928 | ~P1_REG1_REG_28__SCAN_IN;
  assign n10892 = ~P1_REG0_REG_28__SCAN_IN;
  assign n10893 = ~n10926 & ~n10892;
  assign n10895 = ~n10894 & ~n10893;
  assign n15673 = ~n10896 | ~n10895;
  assign n10900 = ~n15585 & ~n14967;
  assign n13882 = ~P2_DATAO_REG_28__SCAN_IN;
  assign n10919 = ~n10912 | ~n10922;
  assign n10916 = ~n15513 & ~n10915;
  assign n10918 = ~n10917 | ~n10916;
  assign n10924 = ~n11100 | ~P1_REG2_REG_29__SCAN_IN;
  assign n10923 = ~n8928 | ~P1_REG1_REG_29__SCAN_IN;
  assign n10928 = ~n10924 | ~n10923;
  assign n10925 = ~P1_REG0_REG_29__SCAN_IN;
  assign n10927 = ~n10926 & ~n10925;
  assign n10929 = ~n10928 & ~n10927;
  assign n10938 = ~n16130 & ~n15515;
  assign n10934 = ~n15998 & ~n15094;
  assign n10931 = ~P1_REG3_REG_28__SCAN_IN | ~P1_U3086;
  assign P1_U3220 = n10942 | n10941;
  assign U123 = P1_WR_REG_SCAN_IN ^ ~P2_WR_REG_SCAN_IN;
  assign U126 = P1_RD_REG_SCAN_IN ^ ~P2_RD_REG_SCAN_IN;
  assign n10944 = ~P1_ADDR_REG_0__SCAN_IN & ~P2_ADDR_REG_0__SCAN_IN;
  assign ADD_1068_U46 = ~n10944 & ~n10943;
  assign n10947 = ~n10946 & ~n10945;
  assign ADD_1068_U5 = n10947 ^ P2_ADDR_REG_1__SCAN_IN;
  assign ADD_1068_U54 = n10949 ^ n10948;
  assign ADD_1068_U53 = n10951 ^ n10950;
  assign ADD_1068_U52 = n10953 ^ ~n10952;
  assign ADD_1068_U51 = n10955 ^ ~n10954;
  assign n10957 = ~P2_D_REG_1__SCAN_IN | ~n10958;
  assign n10956 = ~n11891 | ~n11531;
  assign P2_U3377 = ~n10957 | ~n10956;
  assign n10960 = ~n11524 | ~n11891;
  assign n10959 = ~n10958 | ~P2_D_REG_0__SCAN_IN;
  assign P2_U3376 = ~n10960 | ~n10959;
  assign P1_U3311 = P1_D_REG_14__SCAN_IN & n10963;
  assign P1_U3318 = P1_D_REG_7__SCAN_IN & n10963;
  assign P1_U3312 = P1_D_REG_13__SCAN_IN & n10963;
  assign P1_U3309 = P1_D_REG_16__SCAN_IN & n10963;
  assign P1_U3317 = P1_D_REG_8__SCAN_IN & n10963;
  assign P1_U3310 = P1_D_REG_15__SCAN_IN & n10963;
  assign P1_U3319 = P1_D_REG_6__SCAN_IN & n10963;
  assign P1_U3295 = P1_D_REG_30__SCAN_IN & n10963;
  assign P1_U3294 = P1_D_REG_31__SCAN_IN & n10963;
  assign P1_U3316 = P1_D_REG_9__SCAN_IN & n10963;
  assign P1_U3315 = P1_D_REG_10__SCAN_IN & n10963;
  assign P1_U3298 = P1_D_REG_27__SCAN_IN & n10963;
  assign P1_U3314 = P1_D_REG_11__SCAN_IN & n10963;
  assign P1_U3296 = P1_D_REG_29__SCAN_IN & n10963;
  assign P1_U3320 = P1_D_REG_5__SCAN_IN & n10963;
  assign P1_U3323 = P1_D_REG_2__SCAN_IN & n10963;
  assign P1_U3306 = P1_D_REG_19__SCAN_IN & n10963;
  assign P1_U3305 = P1_D_REG_20__SCAN_IN & n10963;
  assign P1_U3304 = P1_D_REG_21__SCAN_IN & n10963;
  assign P1_U3313 = P1_D_REG_12__SCAN_IN & n10963;
  assign P1_U3321 = P1_D_REG_4__SCAN_IN & n10963;
  assign P1_U3301 = P1_D_REG_24__SCAN_IN & n10963;
  assign P1_U3300 = P1_D_REG_25__SCAN_IN & n10963;
  assign P1_U3299 = P1_D_REG_26__SCAN_IN & n10963;
  assign P1_U3307 = P1_D_REG_18__SCAN_IN & n10963;
  assign P1_U3297 = P1_D_REG_28__SCAN_IN & n10963;
  assign P1_U3303 = P1_D_REG_22__SCAN_IN & n10963;
  assign P1_U3302 = P1_D_REG_23__SCAN_IN & n10963;
  assign P1_U3322 = P1_D_REG_3__SCAN_IN & n10963;
  assign P1_U3308 = P1_D_REG_17__SCAN_IN & n10963;
  assign n10965 = ~P1_D_REG_1__SCAN_IN | ~n10963;
  assign n10964 = n10963 | n10962;
  assign P1_U3440 = ~n10965 | ~n10964;
  assign ADD_1068_U50 = n10967 ^ n10966;
  assign n10979 = P1_U3086 & P1_REG3_REG_0__SCAN_IN;
  assign n10971 = ~n10968 & ~n11667;
  assign n10970 = ~n10969 | ~P1_STATE_REG_SCAN_IN;
  assign n10972 = ~n10971 & ~n10970;
  assign n13673 = ~n14900;
  assign n11185 = ~P1_REG1_REG_0__SCAN_IN;
  assign n10975 = n13673 & n11185;
  assign n10973 = ~P1_REG2_REG_0__SCAN_IN;
  assign n10974 = ~n14900 | ~n10973;
  assign n11381 = ~n11686 | ~n10974;
  assign n10976 = ~n10975 & ~n11381;
  assign n10977 = n10976 ^ ~P1_IR_REG_0__SCAN_IN;
  assign n10978 = ~n11197 & ~n10977;
  assign n10983 = ~n10979 & ~n10978;
  assign n10981 = ~n10980;
  assign n15122 = ~P1_U3085 & ~n10981;
  assign n10982 = ~P1_ADDR_REG_0__SCAN_IN | ~n15122;
  assign P1_U3243 = ~n10983 | ~n10982;
  assign n10985 = ~n11658 & ~P1_D_REG_0__SCAN_IN;
  assign P1_U3439 = ~n10985 & ~n11832;
  assign n10988 = ~n10991 & ~n13123;
  assign n10986 = ~n11251;
  assign n10987 = ~n10986 & ~P1_U3086;
  assign n10990 = ~n10988 & ~n10987;
  assign n10989 = ~n13309 | ~P2_DATAO_REG_6__SCAN_IN;
  assign P1_U3349 = ~n10990 | ~n10989;
  assign n10993 = ~n10991 & ~n13679;
  assign n10992 = ~n11872 & ~P2_U3151;
  assign n10995 = ~n10993 & ~n10992;
  assign n10994 = ~n13683 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P2_U3289 = ~n10995 | ~n10994;
  assign n10998 = ~n10996 & ~n13679;
  assign n10997 = ~n11585 & ~P2_U3151;
  assign n11000 = ~n10998 & ~n10997;
  assign n10999 = ~n13683 | ~P1_DATAO_REG_5__SCAN_IN;
  assign P2_U3290 = ~n11000 | ~n10999;
  assign n11004 = ~n11001 & ~n13679;
  assign n11003 = ~n11002 & ~P2_U3151;
  assign n11006 = ~n11004 & ~n11003;
  assign n11005 = ~n13683 | ~P1_DATAO_REG_2__SCAN_IN;
  assign P2_U3293 = ~n11006 | ~n11005;
  assign n11013 = ~n11007 | ~n14154;
  assign n11008 = ~n11407;
  assign n11011 = ~n11008 & ~P1_U3086;
  assign n11010 = ~n14157 & ~n11009;
  assign n11012 = ~n11011 & ~n11010;
  assign P1_U3353 = ~n11013 | ~n11012;
  assign n11018 = ~n11026 | ~n14154;
  assign n11016 = ~n14157 & ~n11014;
  assign n11455 = ~n11198;
  assign n11015 = ~n11455 & ~P1_U3086;
  assign n11017 = ~n11016 & ~n11015;
  assign P1_U3354 = ~n11018 | ~n11017;
  assign n11023 = ~n11039 | ~n14154;
  assign n11021 = ~n11492 & ~P1_U3086;
  assign n11020 = ~n14157 & ~n11019;
  assign n11022 = ~n11021 & ~n11020;
  assign P1_U3348 = ~n11023 | ~n11022;
  assign ADD_1068_U49 = n11025 ^ ~n11024;
  assign n11028 = ~n11026 | ~n14351;
  assign n11027 = ~n11356 | ~P2_STATE_REG_SCAN_IN;
  assign n11030 = n11028 & n11027;
  assign n11029 = ~n13683 | ~P1_DATAO_REG_1__SCAN_IN;
  assign P2_U3294 = ~n11030 | ~n11029;
  assign n11032 = ~n11044 | ~n14351;
  assign n11031 = ~n11418 | ~P2_STATE_REG_SCAN_IN;
  assign n11034 = n11032 & n11031;
  assign n11033 = ~n13683 | ~P1_DATAO_REG_3__SCAN_IN;
  assign P2_U3292 = ~n11034 | ~n11033;
  assign n11036 = ~n11049 | ~n14351;
  assign n11035 = ~n11570 | ~P2_STATE_REG_SCAN_IN;
  assign n11038 = n11036 & n11035;
  assign n11037 = ~n13683 | ~P1_DATAO_REG_4__SCAN_IN;
  assign P2_U3291 = ~n11038 | ~n11037;
  assign n11041 = ~n11039 | ~n14351;
  assign n11040 = ~n12012 | ~P2_STATE_REG_SCAN_IN;
  assign n11043 = n11041 & n11040;
  assign n11042 = ~n13683 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P2_U3288 = ~n11043 | ~n11042;
  assign n11046 = ~n11044 | ~n14154;
  assign n11201 = ~n11226;
  assign n11045 = ~n11201 | ~P1_STATE_REG_SCAN_IN;
  assign n11048 = n11046 & n11045;
  assign n11047 = ~n13309 | ~P2_DATAO_REG_3__SCAN_IN;
  assign P1_U3352 = ~n11048 | ~n11047;
  assign n11051 = ~n11049 | ~n14154;
  assign n11050 = ~n11359 | ~P1_STATE_REG_SCAN_IN;
  assign n11053 = n11051 & n11050;
  assign n11052 = ~n13309 | ~P2_DATAO_REG_4__SCAN_IN;
  assign P1_U3351 = ~n11053 | ~n11052;
  assign n11059 = ~n11070 | ~n14154;
  assign n11057 = ~n14157 & ~n11054;
  assign n11056 = ~P1_U3086 & ~n11055;
  assign n11058 = ~n11057 & ~n11056;
  assign P1_U3347 = ~n11059 | ~n11058;
  assign n12312 = ~P1_U3973;
  assign n11061 = ~P1_DATAO_REG_19__SCAN_IN | ~n12312;
  assign n11060 = ~P1_U3973 | ~n15901;
  assign P1_U3573 = ~n11061 | ~n11060;
  assign n11063 = ~n12421 | ~P2_U3893;
  assign n11062 = ~n13429 | ~P2_DATAO_REG_2__SCAN_IN;
  assign P2_U3493 = ~n11063 | ~n11062;
  assign n11065 = ~n12420 | ~P2_U3893;
  assign n11064 = ~n13429 | ~P2_DATAO_REG_0__SCAN_IN;
  assign P2_U3491 = ~n11065 | ~n11064;
  assign n11067 = ~n16506 | ~P2_U3893;
  assign n11066 = ~n13429 | ~P2_DATAO_REG_3__SCAN_IN;
  assign P2_U3494 = ~n11067 | ~n11066;
  assign n11069 = ~n16482 | ~P2_U3893;
  assign n11068 = ~n13429 | ~P2_DATAO_REG_1__SCAN_IN;
  assign P2_U3492 = ~n11069 | ~n11068;
  assign n11071 = ~n11070;
  assign n11073 = ~n11071 & ~n13679;
  assign n11072 = ~n12121 & ~P2_U3151;
  assign n11075 = ~n11073 & ~n11072;
  assign n11074 = ~n13683 | ~P1_DATAO_REG_8__SCAN_IN;
  assign P2_U3287 = ~n11075 | ~n11074;
  assign ADD_1068_U48 = n11077 ^ ~n11076;
  assign P2_U3150 = ~P2_U3893 & ~n15398;
  assign n11083 = ~P1_DATAO_REG_31__SCAN_IN | ~n12312;
  assign n11079 = ~n11100 | ~P1_REG2_REG_31__SCAN_IN;
  assign n11078 = ~n8923 | ~P1_REG0_REG_31__SCAN_IN;
  assign n11081 = n11079 & n11078;
  assign n11080 = ~n8928 | ~P1_REG1_REG_31__SCAN_IN;
  assign n11082 = ~P1_U3973 | ~n16133;
  assign P1_U3585 = ~n11083 | ~n11082;
  assign n11085 = ~P2_DATAO_REG_17__SCAN_IN | ~n13429;
  assign n11084 = ~P2_U3893 | ~n16665;
  assign P2_U3508 = ~n11085 | ~n11084;
  assign n11087 = ~n12312 | ~P1_DATAO_REG_9__SCAN_IN;
  assign n11086 = ~n15789 | ~P1_U3973;
  assign P1_U3563 = ~n11087 | ~n11086;
  assign n11089 = ~n12312 | ~P1_DATAO_REG_2__SCAN_IN;
  assign n11088 = ~n12496 | ~P1_U3973;
  assign P1_U3556 = ~n11089 | ~n11088;
  assign n11091 = ~n13076 | ~P1_U3973;
  assign n11090 = ~n12312 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P1_U3565 = ~n11091 | ~n11090;
  assign n11093 = ~P2_DATAO_REG_16__SCAN_IN | ~n13429;
  assign n11092 = ~P2_U3893 | ~n14079;
  assign P2_U3507 = ~n11093 | ~n11092;
  assign n11095 = ~n12312 | ~P1_DATAO_REG_0__SCAN_IN;
  assign n11094 = ~n11719 | ~P1_U3973;
  assign P1_U3554 = ~n11095 | ~n11094;
  assign n11097 = ~n15690 | ~P1_U3973;
  assign n11096 = ~n12312 | ~P1_DATAO_REG_1__SCAN_IN;
  assign P1_U3555 = ~n11097 | ~n11096;
  assign n11099 = ~n16466 | ~P2_U3893;
  assign n11098 = ~n13429 | ~P2_DATAO_REG_12__SCAN_IN;
  assign P2_U3503 = ~n11099 | ~n11098;
  assign n11107 = ~P1_DATAO_REG_30__SCAN_IN | ~n12312;
  assign n11103 = ~n11100 | ~P1_REG2_REG_30__SCAN_IN;
  assign n11102 = ~n8923 | ~P1_REG0_REG_30__SCAN_IN;
  assign n11105 = ~n11103 | ~n11102;
  assign n11104 = n8928 & P1_REG1_REG_30__SCAN_IN;
  assign n11106 = n12312 | n16313;
  assign P1_U3584 = ~n11107 | ~n11106;
  assign n11109 = ~n13859 | ~P2_U3893;
  assign n11108 = ~n13429 | ~P2_DATAO_REG_13__SCAN_IN;
  assign P2_U3504 = ~n11109 | ~n11108;
  assign n11111 = ~n11114 | ~n14351;
  assign n11110 = ~n12518 | ~P2_STATE_REG_SCAN_IN;
  assign n11113 = n11111 & n11110;
  assign n11112 = ~n13683 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P2_U3286 = ~n11113 | ~n11112;
  assign n11116 = ~n11114 | ~n14154;
  assign n11115 = ~n11299 | ~P1_STATE_REG_SCAN_IN;
  assign n11118 = n11116 & n11115;
  assign n11117 = ~n13309 | ~P2_DATAO_REG_9__SCAN_IN;
  assign P1_U3346 = ~n11118 | ~n11117;
  assign n11120 = ~n16631 | ~P2_U3893;
  assign n11119 = ~n13429 | ~P2_DATAO_REG_14__SCAN_IN;
  assign P2_U3505 = ~n11120 | ~n11119;
  assign n11122 = ~n16605 | ~P2_U3893;
  assign n11121 = ~n13429 | ~P2_DATAO_REG_11__SCAN_IN;
  assign P2_U3502 = ~n11122 | ~n11121;
  assign n11124 = ~n13410 | ~P2_U3893;
  assign n11123 = ~n13429 | ~P2_DATAO_REG_9__SCAN_IN;
  assign P2_U3500 = ~n11124 | ~n11123;
  assign n11126 = ~n13503 | ~P1_U3973;
  assign n11125 = ~n12312 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P1_U3564 = ~n11126 | ~n11125;
  assign n11128 = ~n13015 | ~P2_U3893;
  assign n11127 = ~n13429 | ~P2_DATAO_REG_7__SCAN_IN;
  assign P2_U3498 = ~n11128 | ~n11127;
  assign n11130 = ~n12769 | ~P2_U3893;
  assign n11129 = ~n13429 | ~P2_DATAO_REG_6__SCAN_IN;
  assign P2_U3497 = ~n11130 | ~n11129;
  assign n11132 = ~n12997 | ~P2_U3893;
  assign n11131 = ~n13429 | ~P2_DATAO_REG_8__SCAN_IN;
  assign P2_U3499 = ~n11132 | ~n11131;
  assign n11134 = ~P2_DATAO_REG_19__SCAN_IN | ~n13429;
  assign n11133 = ~P2_U3893 | ~n14492;
  assign P2_U3510 = ~n11134 | ~n11133;
  assign n11136 = ~n16645 | ~P2_U3893;
  assign n11135 = ~n13429 | ~P2_DATAO_REG_15__SCAN_IN;
  assign P2_U3506 = ~n11136 | ~n11135;
  assign n11138 = ~n13325 | ~P2_U3893;
  assign n11137 = ~n13429 | ~P2_DATAO_REG_10__SCAN_IN;
  assign P2_U3501 = ~n11138 | ~n11137;
  assign n11140 = ~P1_DATAO_REG_20__SCAN_IN | ~n12312;
  assign n11139 = ~P1_U3973 | ~n15916;
  assign P1_U3574 = ~n11140 | ~n11139;
  assign n11142 = ~n15883 | ~P1_U3973;
  assign n11141 = ~n12312 | ~P1_DATAO_REG_18__SCAN_IN;
  assign P1_U3572 = ~n11142 | ~n11141;
  assign n11144 = ~P2_DATAO_REG_18__SCAN_IN | ~n13429;
  assign n11143 = ~P2_U3893 | ~n16680;
  assign P2_U3509 = ~n11144 | ~n11143;
  assign n11146 = ~n12402 | ~P2_U3893;
  assign n11145 = ~n13429 | ~P2_DATAO_REG_4__SCAN_IN;
  assign P2_U3495 = ~n11146 | ~n11145;
  assign n11148 = ~n12675 | ~P2_U3893;
  assign n11147 = ~n13429 | ~P2_DATAO_REG_5__SCAN_IN;
  assign P2_U3496 = ~n11148 | ~n11147;
  assign n11150 = ~n12312 | ~P1_DATAO_REG_8__SCAN_IN;
  assign n11149 = ~n15773 | ~P1_U3973;
  assign P1_U3562 = ~n11150 | ~n11149;
  assign n11152 = ~n12312 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n11151 = ~n15751 | ~P1_U3973;
  assign P1_U3561 = ~n11152 | ~n11151;
  assign n11154 = ~n12312 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n11153 = ~n12375 | ~P1_U3973;
  assign P1_U3560 = ~n11154 | ~n11153;
  assign n11156 = ~n12312 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n11155 = ~n15850 | ~P1_U3973;
  assign P1_U3568 = ~n11156 | ~n11155;
  assign n11158 = ~P1_DATAO_REG_21__SCAN_IN | ~n12312;
  assign n11157 = ~P1_U3973 | ~n14611;
  assign P1_U3575 = ~n11158 | ~n11157;
  assign n11160 = ~n11163 & ~n13679;
  assign n11159 = ~n13052 & ~P2_U3151;
  assign n11162 = ~n11160 & ~n11159;
  assign n11161 = ~n13683 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P2_U3285 = ~n11162 | ~n11161;
  assign n11166 = ~n11163 & ~n13123;
  assign n11164 = ~n11507;
  assign n11165 = ~n11164 & ~P1_U3086;
  assign n11168 = ~n11166 & ~n11165;
  assign n11167 = ~n13309 | ~P2_DATAO_REG_10__SCAN_IN;
  assign P1_U3345 = ~n11168 | ~n11167;
  assign n11170 = ~n12312 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n11169 = ~n15739 | ~P1_U3973;
  assign P1_U3559 = ~n11170 | ~n11169;
  assign ADD_1068_U47 = n11172 ^ ~n11171;
  assign n11174 = ~n12312 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n11173 = ~n15722 | ~P1_U3973;
  assign P1_U3558 = ~n11174 | ~n11173;
  assign n11176 = ~n12312 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n11175 = ~n14136 | ~P1_U3973;
  assign P1_U3569 = ~n11176 | ~n11175;
  assign n11178 = ~n12312 | ~P1_DATAO_REG_12__SCAN_IN;
  assign n11177 = ~n15820 | ~P1_U3973;
  assign P1_U3566 = ~n11178 | ~n11177;
  assign n11180 = ~n12312 | ~P1_DATAO_REG_3__SCAN_IN;
  assign n11179 = ~n15715 | ~P1_U3973;
  assign P1_U3557 = ~n11180 | ~n11179;
  assign n11182 = ~n12312 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n11181 = ~n13808 | ~P1_U3973;
  assign P1_U3571 = ~n11182 | ~n11181;
  assign n11184 = ~n12312 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n11183 = ~n14060 | ~P1_U3973;
  assign P1_U3570 = ~n11184 | ~n11183;
  assign n12853 = ~P1_REG3_REG_9__SCAN_IN | ~P1_U3086;
  assign n11193 = ~P1_REG1_REG_8__SCAN_IN | ~n11282;
  assign n11447 = n11198 ^ P1_REG1_REG_1__SCAN_IN;
  assign n11446 = ~n11382 & ~n11185;
  assign n11448 = ~n11447 | ~n11446;
  assign n11186 = ~n11198 | ~P1_REG1_REG_1__SCAN_IN;
  assign n11394 = ~n11448 | ~n11186;
  assign n11393 = n11407 ^ P1_REG1_REG_2__SCAN_IN;
  assign n11395 = ~n11394 | ~n11393;
  assign n11187 = ~n11407 | ~P1_REG1_REG_2__SCAN_IN;
  assign n11222 = ~n11395 | ~n11187;
  assign n11221 = n11226 ^ ~P1_REG1_REG_3__SCAN_IN;
  assign n11223 = ~n11222 | ~n11221;
  assign n11188 = ~n11201 | ~P1_REG1_REG_3__SCAN_IN;
  assign n11371 = ~n11223 | ~n11188;
  assign n11370 = n11203 ^ ~P1_REG1_REG_4__SCAN_IN;
  assign n11372 = ~n11371 | ~n11370;
  assign n11189 = ~n11359 | ~P1_REG1_REG_4__SCAN_IN;
  assign n11466 = ~n11372 | ~n11189;
  assign n11465 = n11473 ^ P1_REG1_REG_5__SCAN_IN;
  assign n11467 = ~n11466 | ~n11465;
  assign n11190 = ~n11473 | ~P1_REG1_REG_5__SCAN_IN;
  assign n11240 = ~n11467 | ~n11190;
  assign n11239 = n11251 ^ P1_REG1_REG_6__SCAN_IN;
  assign n11191 = ~n11251 | ~P1_REG1_REG_6__SCAN_IN;
  assign n11484 = n11492 ^ ~P1_REG1_REG_7__SCAN_IN;
  assign n11207 = ~n11492;
  assign n11192 = ~n11207 | ~P1_REG1_REG_7__SCAN_IN;
  assign n11276 = P1_REG1_REG_8__SCAN_IN ^ n11282;
  assign n11194 = n11301 ^ ~n11300;
  assign n11195 = ~n11194 | ~n8934;
  assign n11216 = ~n12853 | ~n11195;
  assign n11196 = ~n11197;
  assign n15119 = ~n14450;
  assign n11214 = ~n15119 | ~n11299;
  assign n16330 = ~n11686 | ~n14900;
  assign n15137 = ~n11197 & ~n16330;
  assign n11210 = ~P1_REG2_REG_8__SCAN_IN & ~n11282;
  assign n11273 = P1_REG2_REG_8__SCAN_IN ^ ~n11282;
  assign n11442 = n11198 ^ P1_REG2_REG_1__SCAN_IN;
  assign n11441 = P1_IR_REG_0__SCAN_IN & P1_REG2_REG_0__SCAN_IN;
  assign n11443 = ~n11442 | ~n11441;
  assign n11199 = ~n11198 | ~P1_REG2_REG_1__SCAN_IN;
  assign n11399 = ~n11443 | ~n11199;
  assign n11398 = n11407 ^ P1_REG2_REG_2__SCAN_IN;
  assign n11400 = ~n11399 | ~n11398;
  assign n11200 = ~n11407 | ~P1_REG2_REG_2__SCAN_IN;
  assign n11228 = ~n11400 | ~n11200;
  assign n11227 = n11226 ^ ~P1_REG2_REG_3__SCAN_IN;
  assign n11229 = ~n11228 | ~n11227;
  assign n11202 = ~n11201 | ~P1_REG2_REG_3__SCAN_IN;
  assign n11363 = ~n11229 | ~n11202;
  assign n11362 = n11203 ^ ~P1_REG2_REG_4__SCAN_IN;
  assign n11364 = ~n11363 | ~n11362;
  assign n11204 = ~n11359 | ~P1_REG2_REG_4__SCAN_IN;
  assign n11461 = ~n11364 | ~n11204;
  assign n11460 = n11473 ^ P1_REG2_REG_5__SCAN_IN;
  assign n11462 = ~n11461 | ~n11460;
  assign n11205 = ~n11473 | ~P1_REG2_REG_5__SCAN_IN;
  assign n11245 = ~n11462 | ~n11205;
  assign n11244 = n11251 ^ P1_REG2_REG_6__SCAN_IN;
  assign n11246 = ~n11245 | ~n11244;
  assign n11206 = ~n11251 | ~P1_REG2_REG_6__SCAN_IN;
  assign n11479 = n11492 ^ ~P1_REG2_REG_7__SCAN_IN;
  assign n11208 = ~n11207 | ~P1_REG2_REG_7__SCAN_IN;
  assign n11291 = n11211 ^ P1_REG2_REG_9__SCAN_IN;
  assign n11212 = n11292 ^ ~n11291;
  assign n11213 = ~n15137 | ~n11212;
  assign n11215 = ~n11214 | ~n11213;
  assign n11218 = ~n11216 & ~n11215;
  assign n11217 = ~n15122 | ~P1_ADDR_REG_9__SCAN_IN;
  assign P1_U3252 = ~n11218 | ~n11217;
  assign n11220 = ~n15836 | ~P1_U3973;
  assign n11219 = ~n12312 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P1_U3567 = ~n11220 | ~n11219;
  assign n11225 = ~n11222 & ~n11221;
  assign n11224 = ~n8934 | ~n11223;
  assign n11236 = ~n11225 & ~n11224;
  assign n11233 = ~n14450 & ~n11226;
  assign n11231 = ~n11228 & ~n11227;
  assign n11230 = ~n15137 | ~n11229;
  assign n11232 = ~n11231 & ~n11230;
  assign n11234 = ~n11233 & ~n11232;
  assign n12499 = ~P1_REG3_REG_3__SCAN_IN | ~P1_U3086;
  assign n11235 = ~n11234 | ~n12499;
  assign n11238 = ~n11236 & ~n11235;
  assign n11237 = ~n15122 | ~P1_ADDR_REG_3__SCAN_IN;
  assign P1_U3246 = ~n11238 | ~n11237;
  assign n11243 = ~n11240 & ~n11239;
  assign n11242 = ~n8934 | ~n11241;
  assign n11255 = ~n11243 & ~n11242;
  assign n11248 = ~n11245 & ~n11244;
  assign n11247 = ~n15137 | ~n11246;
  assign n11250 = ~n11248 & ~n11247;
  assign n12448 = ~P1_STATE_REG_SCAN_IN & ~n11249;
  assign n11253 = ~n11250 & ~n12448;
  assign n11252 = ~n15119 | ~n11251;
  assign n11254 = ~n11253 | ~n11252;
  assign n11257 = ~n11255 & ~n11254;
  assign n11256 = ~P1_ADDR_REG_6__SCAN_IN | ~n15122;
  assign P1_U3249 = ~n11257 | ~n11256;
  assign n11259 = ~n11262 | ~n14154;
  assign n11258 = ~n11609 | ~P1_STATE_REG_SCAN_IN;
  assign n11261 = n11259 & n11258;
  assign n11260 = ~n13309 | ~P2_DATAO_REG_11__SCAN_IN;
  assign P1_U3344 = ~n11261 | ~n11260;
  assign n11264 = ~n11262 | ~n14351;
  assign n11263 = ~n13258 | ~P2_STATE_REG_SCAN_IN;
  assign n11266 = n11264 & n11263;
  assign n11265 = ~n13683 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P2_U3284 = ~n11266 | ~n11265;
  assign n11271 = ~n11435 | ~n14154;
  assign n11269 = ~n14157 & ~n11267;
  assign n11268 = ~P1_U3086 & ~n11600;
  assign n11270 = ~n11269 & ~n11268;
  assign P1_U3343 = ~n11271 | ~n11270;
  assign n11274 = n11273 ^ n11272;
  assign n11601 = ~n15137;
  assign n11286 = ~n11274 & ~n11601;
  assign n11279 = ~n11276 & ~n11275;
  assign n11278 = ~n11277 | ~n8934;
  assign n11281 = ~n11279 & ~n11278;
  assign n12868 = ~P1_STATE_REG_SCAN_IN & ~n11280;
  assign n11284 = ~n11281 & ~n12868;
  assign n11283 = ~n15119 | ~n11282;
  assign n11285 = ~n11284 | ~n11283;
  assign n11288 = ~n11286 & ~n11285;
  assign n11287 = ~P1_ADDR_REG_8__SCAN_IN | ~n15122;
  assign P1_U3251 = ~n11288 | ~n11287;
  assign n11290 = ~P2_DATAO_REG_21__SCAN_IN | ~n13429;
  assign n11289 = ~P2_U3893 | ~n16724;
  assign P2_U3512 = ~n11290 | ~n11289;
  assign n11295 = n11507 ^ P1_REG2_REG_10__SCAN_IN;
  assign n11294 = ~n11299 & ~P1_REG2_REG_9__SCAN_IN;
  assign n11298 = ~n11295 & ~n11296;
  assign n11297 = ~n15137 | ~n11508;
  assign n11313 = ~n11298 & ~n11297;
  assign n11303 = ~n11299 & ~P1_REG1_REG_9__SCAN_IN;
  assign n11307 = ~n11304 & ~n11305;
  assign n11306 = ~n11501 | ~n8934;
  assign n11309 = ~n11307 & ~n11306;
  assign n13284 = ~P1_STATE_REG_SCAN_IN & ~n11308;
  assign n11311 = ~n11309 & ~n13284;
  assign n11310 = ~n15122 | ~P1_ADDR_REG_10__SCAN_IN;
  assign n11312 = ~n11311 | ~n11310;
  assign n11315 = ~n11313 & ~n11312;
  assign n11314 = ~n15119 | ~n11507;
  assign P1_U3253 = ~n11315 | ~n11314;
  assign n11317 = ~n11316;
  assign n11320 = ~n11317 & ~P2_IR_REG_0__SCAN_IN;
  assign n11318 = ~n11320 & ~n11341;
  assign n11334 = ~n15268 & ~n11318;
  assign n11321 = ~n11320 | ~n11319;
  assign n11330 = ~n11322 & ~n11321;
  assign n11325 = ~n15378 | ~n11991;
  assign n11323 = ~P2_REG1_REG_0__SCAN_IN;
  assign n11324 = ~n15371 | ~n11323;
  assign n11326 = ~n11325 | ~n11324;
  assign n11328 = ~n15396 & ~n11326;
  assign n11329 = ~n11328 & ~n11327;
  assign n11332 = ~n11330 & ~n11329;
  assign n11331 = ~P2_REG3_REG_0__SCAN_IN | ~P2_U3151;
  assign n11333 = ~n11332 | ~n11331;
  assign n11336 = ~n11334 & ~n11333;
  assign n11335 = ~P2_ADDR_REG_0__SCAN_IN | ~n15398;
  assign P2_U3182 = ~n11336 | ~n11335;
  assign n11338 = ~P1_DATAO_REG_22__SCAN_IN | ~n12312;
  assign n11337 = ~P1_U3973 | ~n15933;
  assign P1_U3576 = ~n11338 | ~n11337;
  assign n11340 = ~P2_ADDR_REG_1__SCAN_IN | ~n15398;
  assign n11339 = ~P2_REG3_REG_1__SCAN_IN | ~P2_U3151;
  assign n11355 = ~n11340 | ~n11339;
  assign n11343 = n11342 ^ n11341;
  assign n11347 = ~n11343 & ~n15268;
  assign n11345 = n11344 ^ ~P2_REG1_REG_1__SCAN_IN;
  assign n11346 = ~n15182 & ~n11345;
  assign n11353 = ~n11347 & ~n11346;
  assign n11350 = n11349 & n11348;
  assign n11351 = P2_REG2_REG_1__SCAN_IN ^ ~n11350;
  assign n11352 = ~n15378 | ~n11351;
  assign n11354 = ~n11353 | ~n11352;
  assign n11358 = ~n11355 & ~n11354;
  assign n11357 = ~n15396 | ~n11356;
  assign P2_U3183 = ~n11358 | ~n11357;
  assign n11361 = ~n15122 | ~P1_ADDR_REG_4__SCAN_IN;
  assign n11360 = ~n15119 | ~n11359;
  assign n11368 = ~n11361 | ~n11360;
  assign n11366 = ~n11363 & ~n11362;
  assign n11365 = ~n15137 | ~n11364;
  assign n11367 = ~n11366 & ~n11365;
  assign n11369 = ~n11368 & ~n11367;
  assign n12090 = ~P1_REG3_REG_4__SCAN_IN | ~P1_U3086;
  assign n11376 = ~n11369 | ~n12090;
  assign n11374 = ~n11371 & ~n11370;
  assign n11373 = ~n8934 | ~n11372;
  assign n11375 = ~n11374 & ~n11373;
  assign n11388 = ~n11376 & ~n11375;
  assign n11646 = n11378 ^ n11377;
  assign n11379 = ~n11686 | ~n13673;
  assign n11387 = n11646 | n11379;
  assign n11380 = ~n16330;
  assign n11384 = ~n11380 | ~n11441;
  assign n11383 = ~n11382 | ~n11381;
  assign n11385 = ~n11384 | ~n11383;
  assign n11386 = ~n12312 & ~n11385;
  assign n11412 = ~n11387 | ~n11386;
  assign P1_U3247 = ~n11388 | ~n11412;
  assign n11392 = ~n11390 & ~n11389;
  assign ADD_1068_U63 = n11392 ^ n11391;
  assign n11397 = ~n11394 & ~n11393;
  assign n11396 = ~n8934 | ~n11395;
  assign n11411 = ~n11397 & ~n11396;
  assign n11402 = ~n11399 & ~n11398;
  assign n11401 = ~n15137 | ~n11400;
  assign n11406 = ~n11402 & ~n11401;
  assign n11404 = ~P1_ADDR_REG_2__SCAN_IN | ~n15122;
  assign n11403 = ~P1_REG3_REG_2__SCAN_IN | ~P1_U3086;
  assign n11405 = ~n11404 | ~n11403;
  assign n11409 = ~n11406 & ~n11405;
  assign n11408 = ~n15119 | ~n11407;
  assign n11410 = ~n11409 | ~n11408;
  assign n11413 = ~n11411 & ~n11410;
  assign P1_U3245 = ~n11413 | ~n11412;
  assign n11415 = ~P2_DATAO_REG_20__SCAN_IN | ~n13429;
  assign n11414 = ~P2_U3893 | ~n14641;
  assign P2_U3511 = ~n11415 | ~n11414;
  assign n12205 = ~P2_STATE_REG_SCAN_IN & ~n12301;
  assign n11417 = n11416 ^ P2_REG1_REG_3__SCAN_IN;
  assign n11424 = ~n15182 & ~n11417;
  assign n11422 = ~n15396 | ~n11418;
  assign n11420 = n11419 ^ ~P2_REG2_REG_3__SCAN_IN;
  assign n11421 = ~n15378 | ~n11420;
  assign n11423 = ~n11422 | ~n11421;
  assign n11431 = ~n11424 & ~n11423;
  assign n11427 = ~n11426 | ~n11425;
  assign n11429 = ~n11427 | ~n15394;
  assign n11430 = n11429 | n11428;
  assign n11432 = ~n11431 | ~n11430;
  assign n11434 = ~n12205 & ~n11432;
  assign n11433 = ~P2_ADDR_REG_3__SCAN_IN | ~n15398;
  assign P2_U3185 = ~n11434 | ~n11433;
  assign n11436 = ~n11435;
  assign n11438 = ~n11436 & ~n13679;
  assign n11437 = ~n13789 & ~P2_U3151;
  assign n11440 = ~n11438 & ~n11437;
  assign n11439 = ~n13683 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P2_U3283 = ~n11440 | ~n11439;
  assign n11445 = ~n11442 & ~n11441;
  assign n11444 = ~n15137 | ~n11443;
  assign n11452 = ~n11445 & ~n11444;
  assign n11450 = ~n11447 & ~n11446;
  assign n11449 = ~n8934 | ~n11448;
  assign n11451 = ~n11450 & ~n11449;
  assign n11454 = ~n11452 & ~n11451;
  assign n11453 = ~P1_REG3_REG_1__SCAN_IN | ~P1_U3086;
  assign n11457 = ~n11454 | ~n11453;
  assign n11456 = ~n14450 & ~n11455;
  assign n11459 = ~n11457 & ~n11456;
  assign n11458 = ~P1_ADDR_REG_1__SCAN_IN | ~n15122;
  assign P1_U3244 = ~n11459 | ~n11458;
  assign n11464 = ~n11461 & ~n11460;
  assign n11463 = ~n15137 | ~n11462;
  assign n11471 = ~n11464 & ~n11463;
  assign n11469 = ~n11466 & ~n11465;
  assign n11468 = ~n8934 | ~n11467;
  assign n11470 = ~n11469 & ~n11468;
  assign n11472 = ~n11471 & ~n11470;
  assign n12329 = ~P1_REG3_REG_5__SCAN_IN | ~P1_U3086;
  assign n11476 = ~n11472 | ~n12329;
  assign n11474 = ~n11473;
  assign n11475 = ~n14450 & ~n11474;
  assign n11478 = ~n11476 & ~n11475;
  assign n11477 = ~n15122 | ~P1_ADDR_REG_5__SCAN_IN;
  assign P1_U3248 = ~n11478 | ~n11477;
  assign n11483 = ~n11480 & ~n11479;
  assign n11482 = ~n15137 | ~n11481;
  assign n11490 = ~n11483 & ~n11482;
  assign n11488 = ~n11485 & ~n11484;
  assign n11487 = ~n8934 | ~n11486;
  assign n11489 = ~n11488 & ~n11487;
  assign n11491 = ~n11490 & ~n11489;
  assign n12845 = ~P1_REG3_REG_7__SCAN_IN | ~P1_U3086;
  assign n11494 = ~n11491 | ~n12845;
  assign n11493 = ~n14450 & ~n11492;
  assign n11496 = ~n11494 & ~n11493;
  assign n11495 = ~n15122 | ~P1_ADDR_REG_7__SCAN_IN;
  assign P1_U3250 = ~n11496 | ~n11495;
  assign n11500 = ~n14450 & ~n11497;
  assign n11498 = ~n15122 | ~P1_ADDR_REG_11__SCAN_IN;
  assign n13504 = ~P1_REG3_REG_11__SCAN_IN | ~P1_U3086;
  assign n11499 = ~n11498 | ~n13504;
  assign n11514 = ~n11500 & ~n11499;
  assign n11502 = ~n11507 | ~P1_REG1_REG_10__SCAN_IN;
  assign n11506 = ~n11504 & ~n11503;
  assign n11505 = ~n11610 | ~n8934;
  assign n11512 = ~n11506 & ~n11505;
  assign n11509 = ~n11507 | ~P1_REG2_REG_10__SCAN_IN;
  assign n11510 = n11597 ^ n11596;
  assign n11511 = ~n11510 & ~n11601;
  assign n11513 = ~n11512 & ~n11511;
  assign P1_U3254 = ~n11514 | ~n11513;
  assign n11516 = ~n11519 & ~n13679;
  assign n11515 = ~n14034 & ~P2_U3151;
  assign n11518 = ~n11516 & ~n11515;
  assign n11517 = ~n13683 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P2_U3282 = ~n11518 | ~n11517;
  assign n11521 = ~n11519 & ~n13123;
  assign n12149 = ~n12571;
  assign n11520 = ~n12149 & ~P1_U3086;
  assign n11523 = ~n11521 & ~n11520;
  assign n11522 = ~n13309 | ~P2_DATAO_REG_13__SCAN_IN;
  assign P1_U3342 = ~n11523 | ~n11522;
  assign n11985 = ~n11532 & ~n11530;
  assign n11545 = ~P2_REG1_REG_0__SCAN_IN | ~n16444;
  assign n11774 = ~n12420 | ~n16470;
  assign n11536 = ~n16471 | ~n11540;
  assign n16854 = ~n11774 | ~n11536;
  assign n11538 = ~n16854;
  assign n11543 = ~n11538 | ~n11537;
  assign n15559 = ~n11539 | ~n16591;
  assign n11999 = ~n16475 & ~n15559;
  assign n11541 = ~n11540 & ~n16433;
  assign n11542 = ~n11999 & ~n11541;
  assign n11896 = ~n11543 | ~n11542;
  assign n11544 = ~n16442 | ~n11896;
  assign P2_U3459 = ~n11545 | ~n11544;
  assign n11547 = ~P1_DATAO_REG_23__SCAN_IN | ~n12312;
  assign n11546 = ~P1_U3973 | ~n15949;
  assign P1_U3577 = ~n11547 | ~n11546;
  assign n11551 = ~n11549 & ~n11548;
  assign ADD_1068_U62 = n11551 ^ n11550;
  assign n11555 = ~n11554;
  assign n11559 = ~n15386 | ~P2_REG2_REG_5__SCAN_IN;
  assign n11558 = ~n15388 | ~P2_REG1_REG_5__SCAN_IN;
  assign n11561 = ~n11560;
  assign n11565 = ~n15386 | ~P2_REG2_REG_6__SCAN_IN;
  assign n11564 = ~n15388 | ~P2_REG1_REG_6__SCAN_IN;
  assign n11566 = n11859 ^ n11858;
  assign n11593 = ~n11566 & ~n15268;
  assign n11576 = n11853 ^ n11854;
  assign n11579 = ~n11576 & ~n15182;
  assign n12680 = ~P2_REG3_REG_6__SCAN_IN | ~P2_U3151;
  assign n11577 = ~n15398 | ~P2_ADDR_REG_6__SCAN_IN;
  assign n11578 = ~n12680 | ~n11577;
  assign n11591 = ~n11579 & ~n11578;
  assign n11589 = n11874 ^ ~n11873;
  assign n11590 = ~n15378 | ~n11589;
  assign n11592 = ~n11591 | ~n11590;
  assign n11595 = ~n11593 & ~n11592;
  assign n11861 = ~n11872;
  assign n11594 = ~n11861 | ~n15396;
  assign P2_U3188 = ~n11595 | ~n11594;
  assign n11608 = ~n14450 & ~n11600;
  assign n11599 = ~n11609 & ~P1_REG2_REG_11__SCAN_IN;
  assign n12150 = P1_REG2_REG_12__SCAN_IN ^ n11600;
  assign n11602 = n12151 ^ n12150;
  assign n11604 = ~n11602 & ~n11601;
  assign n11606 = ~n11604 & ~n11603;
  assign n11605 = ~n15122 | ~P1_ADDR_REG_12__SCAN_IN;
  assign n11607 = ~n11606 | ~n11605;
  assign n11614 = ~n11608 & ~n11607;
  assign n11611 = ~n11609 | ~P1_REG1_REG_11__SCAN_IN;
  assign n12159 = P1_REG1_REG_12__SCAN_IN ^ ~n12158;
  assign n11612 = n12160 ^ ~n12159;
  assign n11613 = ~n11612 | ~n8934;
  assign P1_U3255 = ~n11614 | ~n11613;
  assign n11620 = ~n11615;
  assign n11617 = ~n11620 & ~n13679;
  assign n11616 = ~n14598 & ~P2_U3151;
  assign n11619 = ~n11617 & ~n11616;
  assign n11618 = ~n13683 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P2_U3281 = ~n11619 | ~n11618;
  assign n11622 = ~n11620 & ~n13123;
  assign n11621 = ~n12564 & ~P1_U3086;
  assign n11624 = ~n11622 & ~n11621;
  assign n11623 = ~n13309 | ~P2_DATAO_REG_14__SCAN_IN;
  assign P1_U3341 = ~n11624 | ~n11623;
  assign n11625 = ~P2_REG3_REG_5__SCAN_IN;
  assign n12191 = ~P2_STATE_REG_SCAN_IN & ~n11625;
  assign n11627 = P2_REG1_REG_5__SCAN_IN ^ n11626;
  assign n11635 = ~n11627 & ~n15182;
  assign n11633 = ~n11628 | ~n15396;
  assign n11631 = n11630 ^ ~n11629;
  assign n11632 = ~n11631 | ~n15394;
  assign n11634 = ~n11633 | ~n11632;
  assign n11639 = ~n11635 & ~n11634;
  assign n11637 = P2_REG2_REG_5__SCAN_IN ^ ~n11636;
  assign n11638 = ~n15378 | ~n11637;
  assign n11640 = ~n11639 | ~n11638;
  assign n11642 = ~n12191 & ~n11640;
  assign n11641 = ~n15398 | ~P2_ADDR_REG_5__SCAN_IN;
  assign P2_U3187 = ~n11642 | ~n11641;
  assign n11645 = n11644 & n11643;
  assign n11739 = ~n11658 | ~n11645;
  assign n11652 = ~P1_REG3_REG_0__SCAN_IN | ~n11739;
  assign n11650 = ~n15515 & ~n15683;
  assign n11648 = ~n15428 | ~n11918;
  assign n11647 = ~n15511 | ~n11646;
  assign n11649 = ~n11648 | ~n11647;
  assign n11651 = ~n11650 & ~n11649;
  assign P1_U3232 = ~n11652 | ~n11651;
  assign n11656 = ~n11654 & ~n11653;
  assign n11657 = n11656 & n11655;
  assign n11673 = ~P1_REG0_REG_0__SCAN_IN | ~n16378;
  assign n15691 = ~n11719 & ~n11922;
  assign n11931 = ~n11719;
  assign n16238 = ~n11931 & ~n11918;
  assign n16158 = ~n15691 & ~n16238;
  assign n15816 = ~n16045;
  assign n15103 = n15816 & n16324;
  assign n14669 = ~n11663 | ~n16365;
  assign n11665 = ~n16236 | ~n16224;
  assign n11664 = ~n16149 | ~n16322;
  assign n15637 = ~n11665 | ~n11664;
  assign n11666 = ~n14669 & ~n15637;
  assign n11671 = n16158 | n11666;
  assign n15533 = ~n11667 & ~n11686;
  assign n11913 = ~n15683 & ~n14935;
  assign n11669 = ~n11922 & ~n11668;
  assign n11670 = ~n11913 & ~n11669;
  assign n11676 = ~n11671 | ~n11670;
  assign n11672 = ~n16377 | ~n11676;
  assign P1_U3453 = ~n11673 | ~n11672;
  assign n11678 = ~P1_REG1_REG_0__SCAN_IN | ~n16383;
  assign n11677 = ~n16381 | ~n11676;
  assign P1_U3522 = ~n11678 | ~n11677;
  assign n11702 = ~P1_REG0_REG_2__SCAN_IN | ~n16378;
  assign n15703 = ~n15691;
  assign n11925 = ~n15683 | ~n15701;
  assign n16237 = ~n15690 | ~n15684;
  assign n11930 = ~n12496;
  assign n16242 = ~n11930 & ~n11812;
  assign n11680 = ~n16242;
  assign n15680 = ~n12496 & ~n12480;
  assign n16245 = ~n15680;
  assign n11815 = ~n11680 | ~n16245;
  assign n11681 = n16235 ^ n11815;
  assign n11690 = ~n11681 & ~n15479;
  assign n11928 = ~n11719 | ~n11918;
  assign n11682 = ~n15683 | ~n15684;
  assign n11685 = ~n11683 | ~n11682;
  assign n15687 = ~n15683 & ~n15684;
  assign n12478 = n11811 ^ ~n11815;
  assign n11688 = n12478 | n11663;
  assign n11687 = ~n15690 | ~n15484;
  assign n11689 = ~n11688 | ~n11687;
  assign n12479 = ~n11690 & ~n11689;
  assign n11699 = ~n12478 & ~n16365;
  assign n11691 = ~n12480 | ~n11922;
  assign n12041 = ~n11691 & ~n15701;
  assign n11694 = ~n12041;
  assign n11692 = ~n15684 | ~n11922;
  assign n11693 = ~n11812 | ~n11692;
  assign n12472 = ~n11694 | ~n11693;
  assign n11697 = n12472 | n15534;
  assign n12482 = ~n15696 & ~n14935;
  assign n11695 = ~n12480 & ~n15536;
  assign n11696 = ~n12482 & ~n11695;
  assign n11698 = ~n11697 | ~n11696;
  assign n11700 = ~n11699 & ~n11698;
  assign n11703 = ~n12479 | ~n11700;
  assign n11701 = ~n16377 | ~n11703;
  assign P1_U3459 = ~n11702 | ~n11701;
  assign n11705 = ~P1_REG1_REG_2__SCAN_IN | ~n16383;
  assign n11704 = ~n16381 | ~n11703;
  assign P1_U3524 = ~n11705 | ~n11704;
  assign n11709 = ~n11707 & ~n11706;
  assign ADD_1068_U61 = n11709 ^ n11708;
  assign n11711 = ~n11714 & ~n13679;
  assign n11710 = ~n14717 & ~P2_U3151;
  assign n11713 = ~n11711 & ~n11710;
  assign n11712 = ~n13683 | ~P1_DATAO_REG_15__SCAN_IN;
  assign P2_U3280 = ~n11713 | ~n11712;
  assign n11716 = ~n11714 & ~n13123;
  assign n11715 = ~n13490 & ~P1_U3086;
  assign n11718 = ~n11716 & ~n11715;
  assign n11717 = ~n13309 | ~P2_DATAO_REG_15__SCAN_IN;
  assign P1_U3340 = ~n11718 | ~n11717;
  assign n11721 = ~n15439 | ~n12496;
  assign n11720 = ~n15521 | ~n11719;
  assign n11730 = ~n11721 | ~n11720;
  assign n11728 = ~n15428 | ~n15701;
  assign n11725 = ~n11723 | ~n11722;
  assign n11726 = n11725 ^ ~n11724;
  assign n11727 = ~n15511 | ~n11726;
  assign n11729 = ~n11728 | ~n11727;
  assign n11732 = ~n11730 & ~n11729;
  assign n11731 = ~P1_REG3_REG_1__SCAN_IN | ~n11739;
  assign P1_U3222 = ~n11732 | ~n11731;
  assign n11734 = ~P2_DATAO_REG_22__SCAN_IN | ~n13429;
  assign n11733 = ~P2_U3893 | ~n16734;
  assign P2_U3513 = ~n11734 | ~n11733;
  assign n11736 = ~P1_DATAO_REG_24__SCAN_IN | ~n12312;
  assign n11735 = ~P1_U3973 | ~n15964;
  assign P1_U3578 = ~n11736 | ~n11735;
  assign n11738 = ~n15439 | ~n15715;
  assign n11737 = ~n15521 | ~n15690;
  assign n11743 = ~n11738 | ~n11737;
  assign n11741 = ~P1_REG3_REG_2__SCAN_IN | ~n11739;
  assign n11740 = ~n15428 | ~n11812;
  assign n11742 = ~n11741 | ~n11740;
  assign n11750 = ~n11743 & ~n11742;
  assign n11746 = ~n11745 | ~n11744;
  assign n11748 = n11747 ^ ~n11746;
  assign n11749 = ~n11748 | ~n15511;
  assign P1_U3237 = ~n11750 | ~n11749;
  assign n11771 = ~P2_REG1_REG_1__SCAN_IN | ~n16444;
  assign n16479 = ~n16476;
  assign n16489 = ~n16482 | ~n16479;
  assign n11772 = ~n16475 | ~n16476;
  assign n16853 = ~n16489 | ~n11772;
  assign n11753 = n16853 ^ ~n11774;
  assign n11752 = n16947 & n11751;
  assign n11758 = ~n11753 & ~n11752;
  assign n16411 = ~n11754 | ~n16591;
  assign n11756 = ~n12420 | ~n16345;
  assign n11755 = ~n12421 | ~n16346;
  assign n11757 = ~n11756 | ~n11755;
  assign n11765 = ~n11758 & ~n11757;
  assign n12724 = n16853 ^ n16472;
  assign n11762 = ~n11759 & ~n16961;
  assign n11764 = ~n12724 | ~n16410;
  assign n12729 = ~n11765 | ~n11764;
  assign n11766 = ~n16476 & ~n16433;
  assign n11769 = ~n12729 & ~n11766;
  assign n16431 = ~n11767 | ~n16961;
  assign n11768 = ~n12724 | ~n13731;
  assign n11899 = ~n11769 | ~n11768;
  assign n11770 = ~n16442 | ~n11899;
  assign P2_U3460 = ~n11771 | ~n11770;
  assign n11799 = ~P2_REG1_REG_2__SCAN_IN | ~n16444;
  assign n11776 = ~n11774 & ~n11773;
  assign n11775 = ~n16489;
  assign n11778 = ~n11776 & ~n11775;
  assign n11777 = ~n16495 & ~n12255;
  assign n12135 = ~n12421 & ~n16496;
  assign n16850 = ~n11777 & ~n12135;
  assign n11790 = ~n16850;
  assign n12131 = ~n11778 | ~n11790;
  assign n11780 = ~n12131;
  assign n11779 = ~n11778 & ~n11790;
  assign n11781 = ~n11780 & ~n11779;
  assign n11785 = ~n11781 & ~n11752;
  assign n11783 = ~n16482 | ~n16345;
  assign n11782 = ~n16506 | ~n16346;
  assign n11784 = ~n11783 | ~n11782;
  assign n11794 = ~n11785 & ~n11784;
  assign n11788 = ~n16482 | ~n16476;
  assign n11787 = ~n16472 | ~n11786;
  assign n11789 = ~n11788 | ~n11787;
  assign n12136 = ~n11790 & ~n11789;
  assign n11792 = ~n12136;
  assign n11791 = ~n11790 | ~n11789;
  assign n12251 = ~n11792 | ~n11791;
  assign n11793 = ~n12251 | ~n16410;
  assign n12253 = ~n11794 | ~n11793;
  assign n11795 = ~n16496 & ~n16433;
  assign n11797 = ~n12253 & ~n11795;
  assign n11796 = ~n12251 | ~n13731;
  assign n11893 = ~n11797 | ~n11796;
  assign n11798 = ~n16442 | ~n11893;
  assign P2_U3461 = ~n11799 | ~n11798;
  assign n11801 = ~n11804 & ~n13679;
  assign n11800 = ~n15206 & ~P2_U3151;
  assign n11803 = ~n11801 & ~n11800;
  assign n11802 = ~n13683 | ~P1_DATAO_REG_16__SCAN_IN;
  assign P2_U3279 = ~n11803 | ~n11802;
  assign n11806 = ~n11804 & ~n13123;
  assign n13828 = ~n14457;
  assign n11805 = ~n13828 & ~P1_U3086;
  assign n11808 = ~n11806 & ~n11805;
  assign n11807 = ~n13309 | ~P2_DATAO_REG_16__SCAN_IN;
  assign P1_U3339 = ~n11808 | ~n11807;
  assign n11828 = ~P1_REG1_REG_3__SCAN_IN | ~n16383;
  assign n11842 = n12041 ^ n15714;
  assign n11810 = ~n11842 & ~n15534;
  assign n11809 = ~n12038 & ~n15536;
  assign n11826 = ~n11810 & ~n11809;
  assign n16063 = ~n15696 & ~n15714;
  assign n16160 = ~n16065 & ~n16063;
  assign n16159 = ~n11815;
  assign n11813 = ~n12496 & ~n11812;
  assign n12043 = ~n11814 & ~n11813;
  assign n11844 = n16160 ^ ~n12043;
  assign n11824 = n11844 & n15103;
  assign n11816 = ~n16235 & ~n11815;
  assign n16064 = ~n11816 & ~n15680;
  assign n11817 = n16160 ^ ~n16064;
  assign n11821 = ~n11817 & ~n15479;
  assign n11819 = ~n12496 | ~n15484;
  assign n11818 = ~n15722 | ~n15533;
  assign n11820 = ~n11819 | ~n11818;
  assign n11823 = ~n11821 & ~n11820;
  assign n11822 = ~n11844 | ~n15057;
  assign n11846 = ~n11823 | ~n11822;
  assign n11825 = ~n11824 & ~n11846;
  assign n11829 = ~n11826 | ~n11825;
  assign n11827 = ~n16381 | ~n11829;
  assign P1_U3525 = ~n11828 | ~n11827;
  assign n11831 = ~P1_REG0_REG_3__SCAN_IN | ~n16378;
  assign n11830 = ~n16377 | ~n11829;
  assign P1_U3462 = ~n11831 | ~n11830;
  assign n11839 = ~n14874 & ~P1_REG3_REG_3__SCAN_IN;
  assign n15660 = ~n15323 & ~n13221;
  assign n11837 = ~n15660 | ~n15714;
  assign n11836 = ~n15323 | ~P1_REG2_REG_3__SCAN_IN;
  assign n11838 = ~n11837 | ~n11836;
  assign n11851 = ~n11839 & ~n11838;
  assign n15074 = ~n11841 | ~n11840;
  assign n11849 = ~n15074 & ~n11842;
  assign n12477 = ~n11843 & ~n8924;
  assign n11845 = n11844 & n12477;
  assign n11847 = ~n11846 & ~n11845;
  assign n11848 = ~n15323 & ~n11847;
  assign n11850 = ~n11849 & ~n11848;
  assign P1_U3290 = ~n11851 | ~n11850;
  assign n12545 = ~P2_STATE_REG_SCAN_IN & ~n11852;
  assign n11857 = P2_REG1_REG_7__SCAN_IN ^ n12005;
  assign n11871 = ~n11857 & ~n15182;
  assign n11869 = ~n12012 | ~n15396;
  assign n11862 = ~n11860;
  assign n11866 = ~n15386 | ~P2_REG2_REG_7__SCAN_IN;
  assign n11865 = ~n15388 | ~P2_REG1_REG_7__SCAN_IN;
  assign n11867 = n12010 ^ ~n12009;
  assign n11868 = ~n11867 | ~n15394;
  assign n11870 = ~n11869 | ~n11868;
  assign n11879 = ~n11871 & ~n11870;
  assign n11877 = P2_REG2_REG_7__SCAN_IN ^ ~n12021;
  assign n11878 = ~n15378 | ~n11877;
  assign n11880 = ~n11879 | ~n11878;
  assign n11882 = ~n12545 & ~n11880;
  assign n11881 = ~n15398 | ~P2_ADDR_REG_7__SCAN_IN;
  assign P2_U3189 = ~n11882 | ~n11881;
  assign n11895 = ~P2_REG0_REG_2__SCAN_IN | ~n16439;
  assign n11894 = ~n16438 | ~n11893;
  assign P2_U3396 = ~n11895 | ~n11894;
  assign n11898 = ~P2_REG0_REG_0__SCAN_IN | ~n16439;
  assign n11897 = ~n16438 | ~n11896;
  assign P2_U3390 = ~n11898 | ~n11897;
  assign n11901 = ~P2_REG0_REG_1__SCAN_IN | ~n16439;
  assign n11900 = ~n16438 | ~n11899;
  assign P2_U3393 = ~n11901 | ~n11900;
  assign n11905 = ~n11903 & ~n11902;
  assign ADD_1068_U60 = n11905 ^ n11904;
  assign n11907 = ~P1_DATAO_REG_25__SCAN_IN | ~n12312;
  assign n11906 = ~P1_U3973 | ~n15969;
  assign P1_U3579 = ~n11907 | ~n11906;
  assign n11909 = ~n15323 | ~P1_REG2_REG_0__SCAN_IN;
  assign n11908 = ~P1_REG3_REG_0__SCAN_IN | ~n15654;
  assign n11917 = ~n11909 | ~n11908;
  assign n11912 = n11911 | n11910;
  assign n11914 = ~n16158 & ~n11912;
  assign n11915 = ~n11914 & ~n11913;
  assign n11916 = ~n15323 & ~n11915;
  assign n11921 = ~n11917 & ~n11916;
  assign n11919 = ~n15497 | ~n15074;
  assign n11920 = ~n11919 | ~n11918;
  assign P1_U3293 = ~n11921 | ~n11920;
  assign n11940 = ~P1_REG0_REG_1__SCAN_IN | ~n16378;
  assign n11948 = n15684 ^ ~n11922;
  assign n11924 = ~n11948 & ~n15534;
  assign n11923 = ~n15684 & ~n15536;
  assign n11938 = ~n11924 & ~n11923;
  assign n11927 = ~n11925;
  assign n11926 = ~n16237;
  assign n16161 = ~n11927 & ~n11926;
  assign n11950 = n16161 ^ ~n11928;
  assign n11936 = ~n11950 & ~n12892;
  assign n11929 = n16161 ^ ~n15691;
  assign n11935 = ~n11929 | ~n15637;
  assign n11933 = ~n11930 & ~n14935;
  assign n11932 = ~n11931 & ~n15639;
  assign n11934 = ~n11933 & ~n11932;
  assign n11952 = ~n11935 | ~n11934;
  assign n11937 = ~n11936 & ~n11952;
  assign n11941 = ~n11938 | ~n11937;
  assign n11939 = ~n16377 | ~n11941;
  assign P1_U3456 = ~n11940 | ~n11939;
  assign n11943 = ~P1_REG1_REG_1__SCAN_IN | ~n16383;
  assign n11942 = ~n16381 | ~n11941;
  assign P1_U3523 = ~n11943 | ~n11942;
  assign n11945 = ~n15323 | ~P1_REG2_REG_1__SCAN_IN;
  assign n11944 = ~P1_REG3_REG_1__SCAN_IN | ~n15654;
  assign n11947 = ~n11945 | ~n11944;
  assign n11946 = ~n15497 & ~n15684;
  assign n11957 = ~n11947 & ~n11946;
  assign n11955 = ~n15074 & ~n11948;
  assign n12952 = ~n11949;
  assign n11951 = ~n11950 & ~n12952;
  assign n11953 = ~n11952 & ~n11951;
  assign n11954 = ~n15323 & ~n11953;
  assign n11956 = ~n11955 & ~n11954;
  assign P1_U3292 = ~n11957 | ~n11956;
  assign n11959 = ~n11962 & ~n13679;
  assign n11958 = ~n15281 & ~P2_U3151;
  assign n11961 = ~n11959 & ~n11958;
  assign n11960 = ~n13683 | ~P1_DATAO_REG_17__SCAN_IN;
  assign P2_U3278 = ~n11961 | ~n11960;
  assign n11964 = ~n11962 & ~n13123;
  assign n14449 = ~n14755;
  assign n11963 = ~n14449 & ~P1_U3086;
  assign n11966 = ~n11964 & ~n11963;
  assign n11965 = ~n13309 | ~P2_DATAO_REG_17__SCAN_IN;
  assign P1_U3338 = ~n11966 | ~n11965;
  assign n11968 = ~n15604 | ~n16506;
  assign n11967 = ~n15342 | ~n12255;
  assign n11977 = ~n11968 | ~n11967;
  assign n11972 = ~n11970 & ~n11969;
  assign n11973 = n11972 ^ ~n11971;
  assign n11975 = ~n11973 | ~n15596;
  assign n11974 = ~n15355 | ~n16482;
  assign n11976 = ~n11975 | ~n11974;
  assign n11979 = ~n11977 & ~n11976;
  assign n14167 = ~n15602;
  assign n11978 = ~P2_REG3_REG_2__SCAN_IN | ~n12424;
  assign P2_U3177 = ~n11979 | ~n11978;
  assign n11981 = ~P2_DATAO_REG_23__SCAN_IN | ~n13429;
  assign n11980 = ~P2_U3893 | ~n15338;
  assign P2_U3514 = ~n11981 | ~n11980;
  assign n11983 = ~n11985;
  assign n11992 = ~n11989 | ~n11988;
  assign n11996 = ~n11991 & ~n16419;
  assign n12307 = n11992 | n15564;
  assign n11994 = ~n16424 | ~n16470;
  assign n11993 = ~n16358 | ~P2_REG3_REG_0__SCAN_IN;
  assign n11995 = ~n11994 | ~n11993;
  assign n12003 = ~n11996 & ~n11995;
  assign n11998 = ~n11997 | ~n16433;
  assign n12000 = ~n16854 & ~n11998;
  assign n12001 = n12000 | n11999;
  assign n12002 = ~n12001 | ~n16419;
  assign P2_U3233 = ~n12003 | ~n12002;
  assign n12008 = n12098 ^ n12099;
  assign n12031 = ~n12008 & ~n15182;
  assign n12013 = ~n12011;
  assign n12017 = ~n15386 | ~P2_REG2_REG_8__SCAN_IN;
  assign n12016 = ~n15388 | ~P2_REG1_REG_8__SCAN_IN;
  assign n12018 = n12108 ^ n12107;
  assign n12027 = ~n12018 & ~n15268;
  assign n13021 = ~P2_REG3_REG_8__SCAN_IN | ~P2_U3151;
  assign n12024 = n12123 ^ ~n12122;
  assign n12025 = ~n12024 | ~n15378;
  assign n12026 = ~n13021 | ~n12025;
  assign n12029 = ~n12027 & ~n12026;
  assign n12028 = ~n15398 | ~P2_ADDR_REG_8__SCAN_IN;
  assign n12030 = ~n12029 | ~n12028;
  assign n12033 = ~n12031 & ~n12030;
  assign n12032 = ~n12110 | ~n15396;
  assign P2_U3190 = ~n12033 | ~n12032;
  assign n12063 = ~n15723;
  assign n12037 = ~n15497 & ~n12063;
  assign n12035 = ~n15323 | ~P1_REG2_REG_4__SCAN_IN;
  assign n12034 = ~n15654 | ~n12084;
  assign n12036 = ~n12035 | ~n12034;
  assign n12059 = ~n12037 & ~n12036;
  assign n12039 = ~n12041 | ~n12038;
  assign n12042 = ~n12039 | ~n15723;
  assign n12040 = ~n15723 & ~n15714;
  assign n12062 = ~n12042 | ~n12348;
  assign n12057 = ~n15074 & ~n12062;
  assign n12343 = ~n15722;
  assign n16067 = ~n12343 & ~n15723;
  assign n12366 = ~n12343 | ~n15723;
  assign n12215 = ~n12235;
  assign n12044 = ~n15715 & ~n15714;
  assign n12236 = ~n12045 & ~n12044;
  assign n12066 = n12215 ^ n12236;
  assign n12049 = ~n12066 & ~n11663;
  assign n12047 = ~n15715 | ~n15484;
  assign n12046 = ~n15739 | ~n15533;
  assign n12048 = ~n12047 | ~n12046;
  assign n12053 = ~n12049 & ~n12048;
  assign n16244 = ~n16065;
  assign n12051 = n12235 ^ ~n12367;
  assign n12052 = ~n12051 | ~n15637;
  assign n12067 = ~n12053 | ~n12052;
  assign n13560 = ~n12477;
  assign n12054 = ~n12066 & ~n13560;
  assign n12055 = ~n12067 & ~n12054;
  assign n12056 = ~n15323 & ~n12055;
  assign n12058 = ~n12057 & ~n12056;
  assign P1_U3289 = ~n12059 | ~n12058;
  assign n12061 = ~P2_DATAO_REG_25__SCAN_IN | ~n13429;
  assign n12060 = ~P2_U3893 | ~n16759;
  assign P2_U3516 = ~n12061 | ~n12060;
  assign n12072 = ~P1_REG0_REG_4__SCAN_IN | ~n16378;
  assign n12065 = ~n12062 & ~n15534;
  assign n12064 = ~n12063 & ~n15536;
  assign n12070 = ~n12065 & ~n12064;
  assign n12068 = ~n12066 & ~n16365;
  assign n12069 = ~n12068 & ~n12067;
  assign n12073 = ~n12070 | ~n12069;
  assign n12071 = ~n16377 | ~n12073;
  assign P1_U3465 = ~n12072 | ~n12071;
  assign n12075 = ~P1_REG1_REG_4__SCAN_IN | ~n16383;
  assign n12074 = ~n16381 | ~n12073;
  assign P1_U3526 = ~n12075 | ~n12074;
  assign n12077 = ~P1_DATAO_REG_26__SCAN_IN | ~n12312;
  assign n12076 = ~P1_U3973 | ~n15520;
  assign P1_U3580 = ~n12077 | ~n12076;
  assign n12081 = ~n12079 & ~n12078;
  assign ADD_1068_U59 = n12081 ^ n12080;
  assign n12083 = ~P2_DATAO_REG_24__SCAN_IN | ~n13429;
  assign n12082 = ~P2_U3893 | ~n15334;
  assign P2_U3515 = ~n12083 | ~n12082;
  assign n12097 = ~n15516 | ~n12084;
  assign n12087 = n12086 ^ ~n12085;
  assign n12095 = ~n12087 & ~n15426;
  assign n12089 = ~n15439 | ~n15739;
  assign n12088 = ~n15521 | ~n15715;
  assign n12093 = ~n12089 | ~n12088;
  assign n12091 = ~n15428 | ~n15723;
  assign n12092 = ~n12091 | ~n12090;
  assign n12094 = n12093 | n12092;
  assign n12096 = ~n12095 & ~n12094;
  assign P1_U3230 = ~n12097 | ~n12096;
  assign n12102 = P2_REG1_REG_9__SCAN_IN ^ n12529;
  assign n12120 = ~n12102 & ~n15182;
  assign n12103 = ~P2_REG3_REG_9__SCAN_IN;
  assign n12963 = ~P2_STATE_REG_SCAN_IN & ~n12103;
  assign n12105 = ~n15398 | ~P2_ADDR_REG_9__SCAN_IN;
  assign n12104 = ~n12518 | ~n15396;
  assign n12106 = ~n12105 | ~n12104;
  assign n12118 = ~n12963 & ~n12106;
  assign n12111 = ~n12109;
  assign n12112 = ~n12111 | ~n12110;
  assign n12115 = ~n15386 | ~P2_REG2_REG_9__SCAN_IN;
  assign n12114 = ~n15388 | ~P2_REG1_REG_9__SCAN_IN;
  assign n12116 = n12516 ^ ~n12515;
  assign n12117 = ~n12116 | ~n15394;
  assign n12119 = ~n12118 | ~n12117;
  assign n12128 = ~n12120 & ~n12119;
  assign n12126 = P2_REG2_REG_9__SCAN_IN ^ ~n12537;
  assign n12127 = ~n15378 | ~n12126;
  assign P2_U3191 = ~n12128 | ~n12127;
  assign n12145 = ~P2_REG1_REG_3__SCAN_IN | ~n16444;
  assign n12129 = ~n16517 & ~n16507;
  assign n12287 = ~n16506 & ~n16516;
  assign n16849 = ~n12129 & ~n12287;
  assign n12285 = ~n16849;
  assign n12130 = ~n16495 | ~n16496;
  assign n12275 = ~n12131 | ~n12130;
  assign n12132 = n12285 ^ ~n12275;
  assign n12134 = ~n12132 | ~n15557;
  assign n12133 = ~n12421 | ~n16345;
  assign n12140 = ~n12134 | ~n12133;
  assign n12286 = ~n12136 & ~n12135;
  assign n12300 = n12285 ^ n12286;
  assign n12138 = n12300 | n15455;
  assign n12137 = ~n12402 | ~n16346;
  assign n12139 = ~n12138 | ~n12137;
  assign n12303 = ~n12140 & ~n12139;
  assign n12142 = ~n12300 & ~n16431;
  assign n12141 = ~n16516 & ~n16433;
  assign n12143 = ~n12142 & ~n12141;
  assign n12146 = ~n12303 | ~n12143;
  assign n12144 = ~n16442 | ~n12146;
  assign P2_U3462 = ~n12145 | ~n12144;
  assign n12148 = ~P2_REG0_REG_3__SCAN_IN | ~n16439;
  assign n12147 = ~n16438 | ~n12146;
  assign P2_U3399 = ~n12148 | ~n12147;
  assign n12171 = ~n14450 & ~n12149;
  assign n12154 = P1_REG2_REG_13__SCAN_IN ^ n12571;
  assign n12153 = ~P1_REG2_REG_12__SCAN_IN & ~n12158;
  assign n12157 = ~n12154 & ~n12155;
  assign n12156 = ~n15137 | ~n12572;
  assign n12168 = ~n12157 & ~n12156;
  assign n12163 = P1_REG1_REG_13__SCAN_IN ^ n12571;
  assign n12162 = ~P1_REG1_REG_12__SCAN_IN & ~n12158;
  assign n12166 = ~n12163 & ~n12164;
  assign n12165 = ~n12558 | ~n8934;
  assign n12167 = ~n12166 & ~n12165;
  assign n12169 = ~n12168 & ~n12167;
  assign n13526 = ~P1_REG3_REG_13__SCAN_IN | ~P1_U3086;
  assign n12170 = ~n12169 | ~n13526;
  assign n12173 = ~n12171 & ~n12170;
  assign n12172 = ~n15122 | ~P1_ADDR_REG_13__SCAN_IN;
  assign P1_U3256 = ~n12173 | ~n12172;
  assign n12175 = ~P1_DATAO_REG_29__SCAN_IN | ~n12312;
  assign n12174 = ~P1_U3973 | ~n16018;
  assign P1_U3583 = ~n12175 | ~n12174;
  assign n12178 = ~n12181 & ~n13679;
  assign n12177 = ~n15381 & ~P2_U3151;
  assign n12180 = ~n12178 & ~n12177;
  assign n12179 = ~n13683 | ~P1_DATAO_REG_18__SCAN_IN;
  assign P2_U3277 = ~n12180 | ~n12179;
  assign n12183 = ~n12181 & ~n13123;
  assign n12182 = ~n14754 & ~P1_U3086;
  assign n12185 = ~n12183 & ~n12182;
  assign n12184 = ~n13309 | ~P2_DATAO_REG_18__SCAN_IN;
  assign P1_U3337 = ~n12185 | ~n12184;
  assign n12188 = n12187 ^ n12186;
  assign n12196 = ~n12188 & ~n15617;
  assign n12190 = ~n15603 & ~n16522;
  assign n12189 = ~n15146 & ~n12761;
  assign n12194 = ~n12190 & ~n12189;
  assign n12192 = ~n15601 & ~n12407;
  assign n12193 = ~n12192 & ~n12191;
  assign n12195 = ~n12194 | ~n12193;
  assign n12198 = ~n12196 & ~n12195;
  assign n12197 = ~n12790 | ~n15602;
  assign P2_U3167 = ~n12198 | ~n12197;
  assign n12200 = n12199 ^ ~n16506;
  assign n12202 = n12201 ^ ~n12200;
  assign n12210 = ~n12202 & ~n15617;
  assign n12204 = ~n15603 & ~n16495;
  assign n12203 = ~n15146 & ~n16522;
  assign n12208 = ~n12204 & ~n12203;
  assign n12206 = ~n15601 & ~n16516;
  assign n12207 = ~n12206 & ~n12205;
  assign n12209 = ~n12208 | ~n12207;
  assign n12212 = ~n12210 & ~n12209;
  assign n12211 = ~n15602 | ~n12301;
  assign P2_U3158 = ~n12212 | ~n12211;
  assign n12214 = ~P1_DATAO_REG_27__SCAN_IN | ~n12312;
  assign n12213 = ~P1_U3973 | ~n15999;
  assign P1_U3581 = ~n12214 | ~n12213;
  assign n12216 = ~n12367 | ~n12215;
  assign n12338 = n12216 & n16249;
  assign n15730 = ~n12349 | ~n15739;
  assign n12341 = ~n15730 | ~n15731;
  assign n12337 = ~n12338 & ~n12341;
  assign n16254 = ~n15730;
  assign n12218 = ~n12337 & ~n16254;
  assign n12447 = ~n12371;
  assign n12362 = ~n12371 & ~n12847;
  assign n12242 = ~n12364 & ~n12362;
  assign n12219 = n12218 ^ ~n12242;
  assign n12223 = ~n12219 & ~n15479;
  assign n12221 = ~n15751 | ~n15533;
  assign n12220 = ~n15739 | ~n15484;
  assign n12222 = ~n12221 | ~n12220;
  assign n12269 = ~n12223 & ~n12222;
  assign n12234 = ~n15323 & ~n12269;
  assign n12224 = ~n12348 & ~n15738;
  assign n12226 = ~n12596;
  assign n12225 = ~n12224 & ~n12371;
  assign n12263 = ~n12226 & ~n12225;
  assign n12230 = n15659 & n12263;
  assign n12228 = ~n15660 | ~n12447;
  assign n12227 = ~n15323 | ~P1_REG2_REG_6__SCAN_IN;
  assign n12229 = ~n12228 | ~n12227;
  assign n12232 = ~n12230 & ~n12229;
  assign n12231 = ~n12449 | ~n15654;
  assign n12233 = ~n12232 | ~n12231;
  assign n12244 = ~n12234 & ~n12233;
  assign n12237 = ~n15722 | ~n15723;
  assign n12342 = ~n12238 | ~n12237;
  assign n15742 = ~n15738 & ~n15739;
  assign n12239 = ~n15742;
  assign n12241 = ~n12342 | ~n12239;
  assign n12240 = ~n15738 | ~n15739;
  assign n12363 = ~n12241 | ~n12240;
  assign n12262 = n12363 ^ ~n12242;
  assign n12918 = ~n14547;
  assign n12243 = n12262 | n12918;
  assign P1_U3287 = ~n12244 | ~n12243;
  assign n12250 = ~P2_REG3_REG_0__SCAN_IN | ~n12424;
  assign n12248 = ~n15617 & ~n16854;
  assign n12246 = ~n15604 | ~n16482;
  assign n12245 = ~n15342 | ~n16470;
  assign n12247 = ~n12246 | ~n12245;
  assign n12249 = ~n12248 & ~n12247;
  assign P2_U3172 = ~n12250 | ~n12249;
  assign n12609 = ~n13871 & ~n16939;
  assign n12252 = n12251 & n12609;
  assign n12254 = ~n12253 & ~n12252;
  assign n12259 = ~n15240 & ~n12254;
  assign n12257 = ~n16424 | ~n12255;
  assign n12256 = ~n15240 | ~P2_REG2_REG_2__SCAN_IN;
  assign n12258 = ~n12257 | ~n12256;
  assign n12261 = ~n12259 & ~n12258;
  assign n12260 = ~n16358 | ~P2_REG3_REG_2__SCAN_IN;
  assign P2_U3231 = ~n12261 | ~n12260;
  assign n12271 = ~P1_REG1_REG_6__SCAN_IN | ~n16383;
  assign n12267 = ~n12262 & ~n12892;
  assign n12265 = ~n12263 | ~n16367;
  assign n12264 = ~n12447 | ~n16369;
  assign n12266 = ~n12265 | ~n12264;
  assign n12268 = ~n12267 & ~n12266;
  assign n12270 = ~n16381 | ~n12272;
  assign P1_U3528 = ~n12271 | ~n12270;
  assign n12274 = ~P1_REG0_REG_6__SCAN_IN | ~n16378;
  assign n12273 = ~n16377 | ~n12272;
  assign P1_U3471 = ~n12274 | ~n12273;
  assign n12295 = ~P2_REG1_REG_4__SCAN_IN | ~n16444;
  assign n12277 = ~n12275 | ~n12285;
  assign n16510 = ~n16506 & ~n16507;
  assign n12276 = ~n16510;
  assign n12278 = n12277 & n12276;
  assign n16855 = n16522 ^ n16523;
  assign n12394 = ~n12278 | ~n16855;
  assign n12279 = ~n12278 & ~n16855;
  assign n12280 = ~n12279 & ~n11752;
  assign n12284 = ~n12394 | ~n12280;
  assign n12282 = ~n16517 & ~n16411;
  assign n12281 = ~n12467 & ~n15559;
  assign n12283 = ~n12282 & ~n12281;
  assign n12290 = ~n12284 | ~n12283;
  assign n12288 = ~n12286 & ~n12285;
  assign n12401 = ~n12288 & ~n12287;
  assign n12663 = n16855 ^ n12401;
  assign n12289 = ~n12663 & ~n15455;
  assign n12668 = n12290 | n12289;
  assign n12291 = ~n16523 & ~n16433;
  assign n12293 = ~n12668 & ~n12291;
  assign n12292 = n12663 | n16431;
  assign n12296 = ~n12293 | ~n12292;
  assign n12294 = ~n16442 | ~n12296;
  assign P2_U3463 = ~n12295 | ~n12294;
  assign n12298 = ~P2_REG0_REG_4__SCAN_IN | ~n16439;
  assign n12297 = ~n16438 | ~n12296;
  assign P2_U3402 = ~n12298 | ~n12297;
  assign n12299 = ~n12609;
  assign n12305 = ~n12300 & ~n12299;
  assign n12302 = ~n16358 | ~n12301;
  assign n12304 = ~n12303 | ~n12302;
  assign n12306 = ~n12305 & ~n12304;
  assign n12309 = ~n15240 & ~n12306;
  assign n12308 = ~n12307 & ~n16516;
  assign n12311 = ~n12309 & ~n12308;
  assign n12310 = ~P2_REG2_REG_3__SCAN_IN | ~n15240;
  assign P2_U3230 = ~n12311 | ~n12310;
  assign n12314 = ~P1_DATAO_REG_28__SCAN_IN | ~n12312;
  assign n12313 = ~P1_U3973 | ~n15673;
  assign P1_U3582 = ~n12314 | ~n12313;
  assign n12318 = ~n12315 & ~n13679;
  assign n12317 = ~n12316;
  assign n12320 = ~n12318 & ~n12317;
  assign n12319 = ~n13683 | ~P1_DATAO_REG_19__SCAN_IN;
  assign P2_U3276 = ~n12320 | ~n12319;
  assign n12336 = ~n15516 | ~n12707;
  assign n12321 = ~n12324;
  assign n12437 = ~n12321 | ~n12322;
  assign n12323 = ~n12322;
  assign n12325 = ~n12324 | ~n12323;
  assign n12326 = n12434 ^ ~n12435;
  assign n12334 = ~n12326 & ~n15426;
  assign n12328 = ~n15439 | ~n12375;
  assign n12327 = ~n15521 | ~n15722;
  assign n12332 = ~n12328 | ~n12327;
  assign n12330 = ~n15428 | ~n15738;
  assign n12331 = ~n12330 | ~n12329;
  assign n12333 = n12332 | n12331;
  assign n12335 = ~n12334 & ~n12333;
  assign P1_U3227 = ~n12336 | ~n12335;
  assign n12358 = ~P1_REG1_REG_5__SCAN_IN | ~n16383;
  assign n12340 = ~n15479 & ~n12337;
  assign n12339 = ~n12338 | ~n12341;
  assign n12347 = ~n12340 | ~n12339;
  assign n12706 = n12342 ^ ~n12341;
  assign n12345 = ~n12706 & ~n11663;
  assign n12344 = ~n12343 & ~n15639;
  assign n12346 = ~n12345 & ~n12344;
  assign n12716 = n12347 & n12346;
  assign n12355 = ~n12706 & ~n16365;
  assign n12717 = n12348 ^ ~n12349;
  assign n12353 = ~n12717 | ~n16367;
  assign n12351 = ~n12847 & ~n14935;
  assign n12350 = ~n12349 & ~n15536;
  assign n12352 = ~n12351 & ~n12350;
  assign n12354 = ~n12353 | ~n12352;
  assign n12356 = ~n12355 & ~n12354;
  assign n12357 = ~n16381 | ~n12359;
  assign P1_U3527 = ~n12358 | ~n12357;
  assign n12361 = ~P1_REG0_REG_5__SCAN_IN | ~n16378;
  assign n12360 = ~n16377 | ~n12359;
  assign P1_U3468 = ~n12361 | ~n12360;
  assign n12387 = ~P1_REG0_REG_7__SCAN_IN | ~n16378;
  assign n15759 = ~n15751;
  assign n16077 = ~n15750 & ~n15759;
  assign n12580 = ~n12365 & ~n12364;
  assign n12379 = ~n12696 & ~n11663;
  assign n12368 = ~n15731 | ~n16067;
  assign n12369 = ~n12368 | ~n15730;
  assign n16166 = ~n12371 & ~n12375;
  assign n12585 = ~n12373 & ~n16170;
  assign n12588 = ~n12585 & ~n15479;
  assign n12374 = ~n12373 | ~n16170;
  assign n12377 = ~n12588 | ~n12374;
  assign n12376 = ~n12375 | ~n15484;
  assign n12378 = ~n12377 | ~n12376;
  assign n12384 = ~n12696 & ~n16365;
  assign n12697 = n12596 ^ ~n15750;
  assign n12382 = ~n12697 & ~n15534;
  assign n12380 = ~n15750 | ~n16369;
  assign n12693 = ~n15773 | ~n15533;
  assign n12381 = ~n12380 | ~n12693;
  assign n12383 = n12382 | n12381;
  assign n12385 = ~n12384 & ~n12383;
  assign n12386 = ~n16377 | ~n12388;
  assign P1_U3474 = ~n12387 | ~n12386;
  assign n12390 = ~P1_REG1_REG_7__SCAN_IN | ~n16383;
  assign n12389 = ~n16381 | ~n12388;
  assign P1_U3529 = ~n12390 | ~n12389;
  assign n12412 = ~P2_REG1_REG_5__SCAN_IN | ~n16444;
  assign n12393 = ~n12402 | ~n12662;
  assign n12617 = ~n12394 | ~n12393;
  assign n12395 = n16851 ^ ~n12617;
  assign n12399 = ~n12395 & ~n11752;
  assign n12397 = ~n12402 | ~n16345;
  assign n12396 = ~n12769 | ~n16346;
  assign n12398 = ~n12397 | ~n12396;
  assign n12406 = ~n12399 & ~n12398;
  assign n12616 = ~n16851;
  assign n12404 = ~n12401 | ~n12400;
  assign n12403 = ~n12402 | ~n16523;
  assign n12607 = ~n12404 | ~n12403;
  assign n12794 = n12616 ^ n12607;
  assign n12405 = ~n12794 | ~n16410;
  assign n12799 = ~n12406 | ~n12405;
  assign n12408 = ~n12407 & ~n16433;
  assign n12410 = ~n12799 & ~n12408;
  assign n12409 = ~n12794 | ~n13731;
  assign n12413 = ~n12410 | ~n12409;
  assign n12411 = ~n16442 | ~n12413;
  assign P2_U3464 = ~n12412 | ~n12411;
  assign n12415 = ~P2_REG0_REG_5__SCAN_IN | ~n16439;
  assign n12414 = ~n16438 | ~n12413;
  assign P2_U3405 = ~n12415 | ~n12414;
  assign n12419 = ~n12417 & ~n12416;
  assign ADD_1068_U58 = n12419 ^ n12418;
  assign n12423 = ~n15355 | ~n12420;
  assign n12422 = ~n15604 | ~n12421;
  assign n12428 = ~n12423 | ~n12422;
  assign n12426 = ~P2_REG3_REG_1__SCAN_IN | ~n12424;
  assign n12425 = ~n15342 | ~n16479;
  assign n12427 = ~n12426 | ~n12425;
  assign n12433 = ~n12428 & ~n12427;
  assign n12431 = n12430 ^ ~n12429;
  assign n12432 = ~n15596 | ~n12431;
  assign P2_U3162 = ~n12433 | ~n12432;
  assign n12436 = ~n12434;
  assign n12438 = ~n12436 | ~n12435;
  assign n12443 = ~n12438 | ~n12437;
  assign n12441 = ~n12439;
  assign n12442 = ~n12441 & ~n12440;
  assign n12444 = n12443 ^ ~n12442;
  assign n12457 = ~n12444 | ~n15511;
  assign n12446 = ~n15439 | ~n15751;
  assign n12445 = ~n15521 | ~n15739;
  assign n12455 = ~n12446 | ~n12445;
  assign n12453 = ~n15428 | ~n12447;
  assign n12451 = ~n12448;
  assign n12450 = ~n12449 | ~n15516;
  assign n12452 = n12451 & n12450;
  assign n12454 = ~n12453 | ~n12452;
  assign n12456 = ~n12455 & ~n12454;
  assign P1_U3239 = ~n12457 | ~n12456;
  assign n12460 = n12459 ^ n12458;
  assign n12464 = ~n12460 & ~n15617;
  assign n12462 = ~n15355 | ~n16506;
  assign n12461 = ~n15342 | ~n12662;
  assign n12463 = ~n12462 | ~n12461;
  assign n12466 = ~n12464 & ~n12463;
  assign n12469 = ~n12466 | ~n12465;
  assign n12468 = ~n15146 & ~n12467;
  assign n12471 = ~n12469 & ~n12468;
  assign n12470 = ~n15602 | ~n12659;
  assign P2_U3170 = ~n12471 | ~n12470;
  assign n12476 = ~n15074 & ~n12472;
  assign n12474 = ~n15323 | ~P1_REG2_REG_2__SCAN_IN;
  assign n12473 = ~P1_REG3_REG_2__SCAN_IN | ~n15654;
  assign n12475 = ~n12474 | ~n12473;
  assign n12489 = ~n12476 & ~n12475;
  assign n15653 = ~n13226 | ~n12477;
  assign n12487 = ~n15653 & ~n12478;
  assign n12481 = ~n12480 & ~n13221;
  assign n12483 = n12482 | n12481;
  assign n12485 = ~n12484 & ~n12483;
  assign n12486 = ~n12485 & ~n15323;
  assign n12488 = ~n12487 & ~n12486;
  assign P1_U3291 = ~n12489 | ~n12488;
  assign n12495 = ~n12652 | ~n14154;
  assign n12493 = ~n16324 & ~P1_U3086;
  assign n12492 = ~n14157 & ~n12491;
  assign n12494 = ~n12493 & ~n12492;
  assign P1_U3335 = ~n12495 | ~n12494;
  assign n12498 = ~n15521 | ~n12496;
  assign n12497 = ~n15439 | ~n15722;
  assign n12505 = ~n12498 | ~n12497;
  assign n12503 = ~n15428 | ~n15714;
  assign n12501 = ~n12499;
  assign n13502 = ~n15516;
  assign n12500 = ~n13502 & ~P1_REG3_REG_3__SCAN_IN;
  assign n12502 = ~n12501 & ~n12500;
  assign n12504 = ~n12503 | ~n12502;
  assign n12512 = ~n12505 & ~n12504;
  assign n12508 = ~n12507 & ~n12506;
  assign n12510 = n12509 ^ n12508;
  assign n12511 = ~n12510 | ~n15511;
  assign P1_U3218 = ~n12512 | ~n12511;
  assign n12514 = ~n15398 | ~P2_ADDR_REG_10__SCAN_IN;
  assign n12513 = ~n13041 | ~n15396;
  assign n12526 = ~n12514 | ~n12513;
  assign n12519 = ~n12517;
  assign n12520 = ~n12519 | ~n12518;
  assign n12523 = ~n15386 | ~P2_REG2_REG_10__SCAN_IN;
  assign n12522 = ~n15388 | ~P2_REG1_REG_10__SCAN_IN;
  assign n12524 = n13039 ^ n13038;
  assign n12525 = ~n12524 & ~n15268;
  assign n12527 = ~n12526 & ~n12525;
  assign n13415 = ~P2_REG3_REG_10__SCAN_IN | ~P2_U3151;
  assign n12534 = ~n12527 | ~n13415;
  assign n12532 = n13029 ^ n13030;
  assign n12533 = ~n12532 & ~n15182;
  assign n12542 = ~n12534 & ~n12533;
  assign n12540 = n13054 ^ ~n13053;
  assign n12541 = ~n12540 | ~n15378;
  assign P2_U3192 = ~n12542 | ~n12541;
  assign n12544 = ~n15355 | ~n12769;
  assign n12543 = ~n15342 | ~n16551;
  assign n12555 = ~n12544 | ~n12543;
  assign n12546 = ~n15146 & ~n12990;
  assign n12553 = ~n12546 & ~n12545;
  assign n12549 = ~n12548 | ~n12547;
  assign n12551 = ~n12549 | ~n15596;
  assign n12552 = n12551 | n12550;
  assign n12554 = ~n12553 | ~n12552;
  assign n12557 = ~n12555 & ~n12554;
  assign n12556 = ~n12825 | ~n15602;
  assign P2_U3153 = ~n12557 | ~n12556;
  assign n12559 = ~n12571 | ~P1_REG1_REG_13__SCAN_IN;
  assign n12563 = ~n12561 & ~n12560;
  assign n12562 = ~n13488 | ~n8934;
  assign n12570 = ~n12563 & ~n12562;
  assign n12566 = ~n14450 & ~n12564;
  assign n12568 = ~n12566 & ~n12565;
  assign n12567 = ~n15122 | ~P1_ADDR_REG_14__SCAN_IN;
  assign n12569 = ~n12568 | ~n12567;
  assign n12577 = ~n12570 & ~n12569;
  assign n13482 = ~n13487 & ~P1_REG2_REG_14__SCAN_IN;
  assign n13481 = n13487 & P1_REG2_REG_14__SCAN_IN;
  assign n12574 = ~n13482 & ~n13481;
  assign n12573 = ~n12571 | ~P1_REG2_REG_13__SCAN_IN;
  assign n12575 = n12574 ^ n13480;
  assign n12576 = ~n12575 | ~n15137;
  assign P1_U3257 = ~n12577 | ~n12576;
  assign n12603 = ~P1_REG1_REG_8__SCAN_IN | ~n16383;
  assign n12893 = ~n15772 | ~n15777;
  assign n12578 = ~n12893;
  assign n12579 = ~n15754 | ~n15759;
  assign n12581 = ~n15750 | ~n15751;
  assign n12634 = n16173 ^ n12744;
  assign n12584 = ~n12634 & ~n12892;
  assign n12583 = ~n15776 & ~n15536;
  assign n12601 = ~n12584 & ~n12583;
  assign n12739 = ~n12585 & ~n16077;
  assign n12586 = ~n12739 & ~n15479;
  assign n12591 = n12586 | n16173;
  assign n12589 = ~n12588 | ~n12587;
  assign n12590 = ~n12589 | ~n16173;
  assign n12595 = ~n12591 | ~n12590;
  assign n12593 = ~n15759 & ~n15639;
  assign n12592 = ~n12900 & ~n14935;
  assign n12594 = ~n12593 & ~n12592;
  assign n12597 = ~n12596 & ~n15750;
  assign n12598 = n15776 | n12597;
  assign n12633 = ~n12598 | ~n12747;
  assign n12599 = ~n12633 & ~n15534;
  assign n12600 = ~n12636 & ~n12599;
  assign n12602 = ~n16381 | ~n12604;
  assign P1_U3530 = ~n12603 | ~n12602;
  assign n12606 = ~P1_REG0_REG_8__SCAN_IN | ~n16378;
  assign n12605 = ~n16377 | ~n12604;
  assign P1_U3477 = ~n12606 | ~n12605;
  assign n12608 = ~n12607 & ~n16540;
  assign n12774 = ~n12608 & ~n16542;
  assign n12642 = n16859 ^ n12774;
  assign n16423 = ~n16419 | ~n12609;
  assign n12613 = ~n12642 & ~n16423;
  assign n12611 = ~n15240 | ~P2_REG2_REG_6__SCAN_IN;
  assign n12610 = ~n16424 | ~n12765;
  assign n12612 = ~n12611 | ~n12610;
  assign n12628 = ~n12613 & ~n12612;
  assign n12625 = ~n16358 | ~n12684;
  assign n12615 = n12642 | n15455;
  assign n12614 = ~n12675 | ~n16345;
  assign n12624 = ~n12615 | ~n12614;
  assign n12619 = ~n12617 & ~n12616;
  assign n12618 = ~n12793 & ~n12675;
  assign n12764 = ~n12619 & ~n12618;
  assign n12620 = n16859 ^ n12764;
  assign n12622 = ~n12620 | ~n15557;
  assign n12621 = ~n13015 | ~n16346;
  assign n12623 = ~n12622 | ~n12621;
  assign n12646 = ~n12624 & ~n12623;
  assign n12626 = ~n12625 | ~n12646;
  assign n12627 = ~n12626 | ~n16419;
  assign P2_U3227 = ~n12628 | ~n12627;
  assign n12630 = ~n15323 | ~P1_REG2_REG_8__SCAN_IN;
  assign n12629 = ~n12879 | ~n15654;
  assign n12632 = ~n12630 | ~n12629;
  assign n12631 = ~n15497 & ~n15776;
  assign n12641 = ~n12632 & ~n12631;
  assign n12639 = ~n12633 & ~n15074;
  assign n12635 = ~n12634 & ~n12952;
  assign n12637 = ~n12636 & ~n12635;
  assign n12638 = ~n15323 & ~n12637;
  assign n12640 = ~n12639 & ~n12638;
  assign P1_U3285 = ~n12641 | ~n12640;
  assign n12648 = ~P2_REG0_REG_6__SCAN_IN | ~n16439;
  assign n12644 = ~n12642 & ~n16431;
  assign n12643 = ~n12762 & ~n16433;
  assign n12645 = ~n12644 & ~n12643;
  assign n12647 = ~n16438 | ~n12649;
  assign P2_U3408 = ~n12648 | ~n12647;
  assign n12651 = ~P2_REG1_REG_6__SCAN_IN | ~n16444;
  assign n12650 = ~n16442 | ~n12649;
  assign P2_U3465 = ~n12651 | ~n12650;
  assign n12656 = n12654 & n12653;
  assign n12655 = ~n13683 | ~P1_DATAO_REG_20__SCAN_IN;
  assign P2_U3275 = ~n12656 | ~n12655;
  assign n12658 = ~P2_DATAO_REG_26__SCAN_IN | ~n13429;
  assign n12657 = ~P2_U3893 | ~n15572;
  assign P2_U3517 = ~n12658 | ~n12657;
  assign n12661 = ~n15240 | ~P2_REG2_REG_4__SCAN_IN;
  assign n12660 = ~n16358 | ~n12659;
  assign n12667 = ~n12661 | ~n12660;
  assign n12665 = ~n16424 | ~n12662;
  assign n12664 = n12663 | n16423;
  assign n12666 = ~n12665 | ~n12664;
  assign n12670 = ~n12667 & ~n12666;
  assign n12669 = ~n12668 | ~n16419;
  assign P2_U3229 = ~n12670 | ~n12669;
  assign n12672 = n12671 ^ ~n12769;
  assign n12674 = n12673 ^ ~n12672;
  assign n12679 = ~n12674 & ~n15617;
  assign n12677 = ~n15355 | ~n12675;
  assign n12676 = ~n15342 | ~n12765;
  assign n12678 = ~n12677 | ~n12676;
  assign n12681 = ~n12679 & ~n12678;
  assign n12683 = ~n12681 | ~n12680;
  assign n12682 = ~n15146 & ~n16550;
  assign n12686 = ~n12683 & ~n12682;
  assign n12685 = ~n15602 | ~n12684;
  assign P2_U3179 = ~n12686 | ~n12685;
  assign n12690 = ~n12688 & ~n12687;
  assign ADD_1068_U57 = n12690 ^ n12689;
  assign n12692 = ~n15660 | ~n15750;
  assign n12691 = ~n15323 | ~P1_REG2_REG_7__SCAN_IN;
  assign n12703 = ~n12692 | ~n12691;
  assign n12695 = ~n12694 | ~n12693;
  assign n12701 = ~n12695 | ~n13226;
  assign n12699 = ~n12696 & ~n15653;
  assign n12698 = ~n15074 & ~n12697;
  assign n12700 = ~n12699 & ~n12698;
  assign n12702 = ~n12701 | ~n12700;
  assign n12705 = ~n12703 & ~n12702;
  assign n12704 = ~n15654 | ~n12850;
  assign P1_U3286 = ~n12705 | ~n12704;
  assign n12715 = ~n12706 & ~n15653;
  assign n12709 = ~n15660 | ~n15738;
  assign n12708 = ~n15654 | ~n12707;
  assign n12711 = ~n12709 | ~n12708;
  assign n12710 = ~n15502 & ~n12847;
  assign n12713 = ~n12711 & ~n12710;
  assign n12712 = ~n15323 | ~P1_REG2_REG_5__SCAN_IN;
  assign n12714 = ~n12713 | ~n12712;
  assign n12721 = ~n12715 & ~n12714;
  assign n12719 = ~n15323 & ~n12716;
  assign n12718 = n15659 & n12717;
  assign n12720 = ~n12719 & ~n12718;
  assign P1_U3288 = ~n12721 | ~n12720;
  assign n12723 = ~n16358 | ~P2_REG3_REG_1__SCAN_IN;
  assign n12722 = ~n15240 | ~P2_REG2_REG_1__SCAN_IN;
  assign n12728 = ~n12723 | ~n12722;
  assign n12726 = ~n16424 | ~n16479;
  assign n12725 = ~n13390 | ~n12724;
  assign n12727 = ~n12726 | ~n12725;
  assign n12731 = ~n12728 & ~n12727;
  assign n12730 = ~n12729 | ~n16419;
  assign P2_U3232 = ~n12731 | ~n12730;
  assign n12732 = ~n12785;
  assign n12737 = ~n12732 | ~n14154;
  assign n16218 = ~n16236;
  assign n12735 = ~n16218 & ~P1_U3086;
  assign n12734 = ~n14157 & ~n12733;
  assign n12736 = ~n12735 & ~n12734;
  assign P1_U3334 = ~n12737 | ~n12736;
  assign n12757 = ~P1_REG1_REG_9__SCAN_IN | ~n16383;
  assign n12738 = ~n16078;
  assign n12896 = ~n12739 | ~n12738;
  assign n12741 = n12740 ^ ~n16175;
  assign n12743 = ~n12741 & ~n15479;
  assign n12742 = ~n15777 & ~n15639;
  assign n12745 = ~n15772 & ~n15773;
  assign n12890 = ~n12746 & ~n12745;
  assign n12919 = n16175 ^ ~n12890;
  assign n12754 = ~n12919 & ~n12892;
  assign n12907 = ~n15788 & ~n12747;
  assign n12906 = ~n12907;
  assign n12748 = ~n15788 | ~n12747;
  assign n12930 = ~n12906 | ~n12748;
  assign n12752 = n12930 | n15534;
  assign n12750 = ~n12889 & ~n15536;
  assign n12749 = ~n15803 & ~n14935;
  assign n12751 = ~n12750 & ~n12749;
  assign n12753 = ~n12752 | ~n12751;
  assign n12755 = ~n12754 & ~n12753;
  assign n12756 = ~n16381 | ~n12758;
  assign P1_U3531 = ~n12757 | ~n12756;
  assign n12760 = ~P1_REG0_REG_9__SCAN_IN | ~n16378;
  assign n12759 = ~n16377 | ~n12758;
  assign P1_U3480 = ~n12760 | ~n12759;
  assign n12781 = ~P2_REG1_REG_7__SCAN_IN | ~n16444;
  assign n16861 = n16551 ^ n16550;
  assign n12763 = ~n12762 | ~n12761;
  assign n12767 = ~n12764 | ~n12763;
  assign n12766 = ~n12765 | ~n12769;
  assign n12812 = ~n12767 | ~n12766;
  assign n12768 = n16861 ^ n12812;
  assign n12773 = ~n12768 & ~n11752;
  assign n12771 = ~n12769 | ~n16345;
  assign n12770 = ~n12997 | ~n16346;
  assign n12772 = ~n12771 | ~n12770;
  assign n12777 = ~n12773 & ~n12772;
  assign n12775 = ~n12774 | ~n16548;
  assign n12804 = ~n12775 | ~n16553;
  assign n12824 = n16861 ^ n12804;
  assign n12776 = ~n12824 | ~n16410;
  assign n12826 = ~n12810 & ~n16433;
  assign n12779 = ~n12830 & ~n12826;
  assign n12778 = ~n12824 | ~n13731;
  assign n12780 = ~n16442 | ~n12782;
  assign P2_U3466 = ~n12781 | ~n12780;
  assign n12784 = ~P2_REG0_REG_7__SCAN_IN | ~n16439;
  assign n12783 = ~n16438 | ~n12782;
  assign P2_U3411 = ~n12784 | ~n12783;
  assign n12787 = ~n12785 & ~n13679;
  assign n12786 = ~n16939 & ~P2_U3151;
  assign n12789 = ~n12787 & ~n12786;
  assign n12788 = ~n13683 | ~P1_DATAO_REG_21__SCAN_IN;
  assign P2_U3274 = ~n12789 | ~n12788;
  assign n12792 = ~P2_REG2_REG_5__SCAN_IN | ~n15240;
  assign n12791 = ~n16358 | ~n12790;
  assign n12798 = ~n12792 | ~n12791;
  assign n12796 = ~n16424 | ~n12793;
  assign n12795 = ~n12794 | ~n13390;
  assign n12797 = ~n12796 | ~n12795;
  assign n12801 = ~n12798 & ~n12797;
  assign n12800 = ~n12799 | ~n16419;
  assign P2_U3228 = ~n12801 | ~n12800;
  assign n12803 = ~P2_REG2_REG_8__SCAN_IN | ~n15240;
  assign n12802 = ~n16358 | ~n13026;
  assign n12809 = ~n12803 | ~n12802;
  assign n12807 = ~n16424 | ~n13016;
  assign n12805 = ~n12804 | ~n16861;
  assign n12984 = ~n12805 | ~n16560;
  assign n12806 = ~n12939 | ~n13390;
  assign n12808 = ~n12807 | ~n12806;
  assign n12823 = ~n12809 & ~n12808;
  assign n12811 = ~n12810 | ~n16550;
  assign n12813 = ~n16551 | ~n13015;
  assign n12993 = ~n12814 | ~n12813;
  assign n12815 = n16863 ^ ~n12993;
  assign n12819 = ~n12815 & ~n11752;
  assign n12817 = ~n13410 | ~n16346;
  assign n12816 = ~n13015 | ~n16345;
  assign n12818 = ~n12817 | ~n12816;
  assign n12821 = ~n12819 & ~n12818;
  assign n12820 = ~n12939 | ~n16410;
  assign n12822 = ~n12938 | ~n16419;
  assign P2_U3225 = ~n12823 | ~n12822;
  assign n12833 = n12824 & n13390;
  assign n12828 = ~n16358 | ~n12825;
  assign n12827 = ~n12826 | ~n13871;
  assign n12829 = ~n12828 | ~n12827;
  assign n12831 = ~n12830 & ~n12829;
  assign n12832 = ~n12831 & ~n15240;
  assign n12835 = ~n12833 & ~n12832;
  assign n12834 = ~n15240 | ~P2_REG2_REG_7__SCAN_IN;
  assign P2_U3226 = ~n12835 | ~n12834;
  assign n12838 = ~n12837 | ~n12836;
  assign n12840 = n12839 ^ ~n12838;
  assign n12844 = ~n12840 & ~n15426;
  assign n12842 = ~n15439 | ~n15773;
  assign n12841 = ~n15428 | ~n15750;
  assign n12843 = ~n12842 | ~n12841;
  assign n12846 = ~n12844 & ~n12843;
  assign n12849 = ~n12846 | ~n12845;
  assign n12848 = ~n15094 & ~n12847;
  assign n12852 = ~n12849 & ~n12848;
  assign n12851 = ~n12850 | ~n15516;
  assign P1_U3213 = ~n12852 | ~n12851;
  assign n12854 = ~n15521 | ~n15773;
  assign n12856 = ~n12854 | ~n12853;
  assign n12855 = ~n15515 & ~n15803;
  assign n12865 = ~n12856 & ~n12855;
  assign n12859 = n12858 ^ n12857;
  assign n12863 = ~n12859 & ~n15426;
  assign n12861 = ~n15516 | ~n12920;
  assign n12860 = ~n15428 | ~n15788;
  assign n12862 = ~n12861 | ~n12860;
  assign n12864 = ~n12863 & ~n12862;
  assign P1_U3231 = ~n12865 | ~n12864;
  assign n12867 = ~n15439 | ~n15789;
  assign n12866 = ~n15428 | ~n15772;
  assign n12878 = ~n12867 | ~n12866;
  assign n12869 = ~n15094 & ~n15759;
  assign n12876 = ~n12869 & ~n12868;
  assign n12874 = n12873 ^ ~n12872;
  assign n12881 = ~n12878 & ~n12877;
  assign n12880 = ~n12879 | ~n15516;
  assign P1_U3221 = ~n12881 | ~n12880;
  assign n12885 = ~n16332 & ~P1_U3086;
  assign n12884 = ~n14157 & ~n12883;
  assign n12886 = ~n12885 & ~n12884;
  assign P1_U3333 = ~n12887 | ~n12886;
  assign n12914 = ~P1_REG0_REG_10__SCAN_IN | ~n16378;
  assign n16177 = ~n12888 & ~n16076;
  assign n13063 = ~n12891 | ~n15792;
  assign n12905 = ~n12953 & ~n12892;
  assign n12894 = ~n15788 | ~n12900;
  assign n16083 = ~n12894 | ~n12893;
  assign n12895 = ~n16083;
  assign n12898 = ~n12896 | ~n12895;
  assign n16075 = ~n15788 & ~n12900;
  assign n12897 = ~n16075;
  assign n12899 = n16177 ^ n13073;
  assign n12902 = ~n12900 & ~n15639;
  assign n12901 = ~n13283 & ~n14935;
  assign n12903 = ~n12902 & ~n12901;
  assign n12908 = ~n13293 | ~n12906;
  assign n12951 = ~n12908 | ~n13141;
  assign n12910 = ~n12951 & ~n15534;
  assign n12909 = ~n15802 & ~n15536;
  assign n12911 = ~n12910 & ~n12909;
  assign P1_U3483 = ~n12914 | ~n12913;
  assign n12917 = ~P1_REG1_REG_10__SCAN_IN | ~n16383;
  assign n12916 = ~n16381 | ~n12915;
  assign P1_U3532 = ~n12917 | ~n12916;
  assign n12928 = ~n12919 & ~n12918;
  assign n12922 = ~n15323 | ~P1_REG2_REG_9__SCAN_IN;
  assign n12921 = ~n12920 | ~n15654;
  assign n12926 = ~n12922 | ~n12921;
  assign n15083 = ~n15502;
  assign n12924 = ~n15083 | ~n13503;
  assign n12923 = ~n15660 | ~n15788;
  assign n12925 = ~n12924 | ~n12923;
  assign n12927 = n12926 | n12925;
  assign n12934 = ~n12928 & ~n12927;
  assign n12932 = ~n15323 & ~n12929;
  assign n12931 = ~n12930 & ~n15074;
  assign n12933 = ~n12932 & ~n12931;
  assign P1_U3284 = ~n12934 | ~n12933;
  assign n12936 = ~P2_DATAO_REG_27__SCAN_IN | ~n13429;
  assign n12935 = ~P2_U3893 | ~n16779;
  assign P2_U3518 = ~n12936 | ~n12935;
  assign n12943 = ~P2_REG0_REG_8__SCAN_IN | ~n16439;
  assign n12991 = ~n13016;
  assign n12937 = ~n12991 & ~n16433;
  assign n12941 = ~n12938 & ~n12937;
  assign n12940 = ~n12939 | ~n13731;
  assign n12942 = ~n16438 | ~n12944;
  assign P2_U3414 = ~n12943 | ~n12942;
  assign n12946 = ~P2_REG1_REG_8__SCAN_IN | ~n16444;
  assign n12945 = ~n16442 | ~n12944;
  assign P2_U3467 = ~n12946 | ~n12945;
  assign n12948 = ~n15323 | ~P1_REG2_REG_10__SCAN_IN;
  assign n12947 = ~n13298 | ~n15654;
  assign n12950 = ~n12948 | ~n12947;
  assign n12949 = ~n15497 & ~n15802;
  assign n12960 = ~n12950 & ~n12949;
  assign n12958 = ~n12951 & ~n15074;
  assign n12954 = ~n12953 & ~n12952;
  assign n12956 = ~n12955 & ~n12954;
  assign n12957 = ~n15323 & ~n12956;
  assign n12959 = ~n12958 & ~n12957;
  assign P1_U3283 = ~n12960 | ~n12959;
  assign n12962 = ~n15355 | ~n12997;
  assign n12961 = ~n15342 | ~n13315;
  assign n12973 = ~n12962 | ~n12961;
  assign n12964 = ~n15146 & ~n13101;
  assign n12971 = ~n12964 & ~n12963;
  assign n12967 = ~n12966 | ~n12965;
  assign n12969 = ~n12967 | ~n15596;
  assign n12970 = n12969 | n12968;
  assign n12975 = ~n12973 & ~n12972;
  assign n12974 = ~n12981 | ~n15602;
  assign P2_U3171 = ~n12975 | ~n12974;
  assign n12977 = ~n16961 & ~P2_U3151;
  assign n12980 = ~n12978 & ~n12977;
  assign n12979 = ~n13683 | ~P1_DATAO_REG_22__SCAN_IN;
  assign P2_U3273 = ~n12980 | ~n12979;
  assign n12983 = ~P2_REG2_REG_9__SCAN_IN | ~n15240;
  assign n12982 = ~n16358 | ~n12981;
  assign n12989 = ~n12983 | ~n12982;
  assign n12987 = ~n16424 | ~n13315;
  assign n12985 = ~n12984 | ~n16574;
  assign n13102 = ~n12985 | ~n16570;
  assign n12986 = ~n13132 | ~n13390;
  assign n12988 = ~n12987 | ~n12986;
  assign n13005 = ~n12989 & ~n12988;
  assign n12992 = ~n12991 | ~n12990;
  assign n12995 = ~n12993 | ~n12992;
  assign n12996 = n16866 ^ n13314;
  assign n13001 = ~n12996 & ~n11752;
  assign n12999 = ~n13325 | ~n16346;
  assign n12998 = ~n12997 | ~n16345;
  assign n13000 = ~n12999 | ~n12998;
  assign n13003 = ~n13001 & ~n13000;
  assign n13002 = ~n13132 | ~n16410;
  assign n13004 = ~n13131 | ~n16419;
  assign P2_U3224 = ~n13005 | ~n13004;
  assign n13009 = ~n13007 & ~n13006;
  assign ADD_1068_U56 = n13009 ^ n13008;
  assign n13012 = ~n13011 & ~n13010;
  assign n13014 = n13013 ^ n13012;
  assign n13020 = ~n13014 & ~n15617;
  assign n13018 = ~n15355 | ~n13015;
  assign n13017 = ~n15342 | ~n13016;
  assign n13019 = ~n13018 | ~n13017;
  assign n13022 = ~n13020 & ~n13019;
  assign n13025 = ~n13022 | ~n13021;
  assign n13024 = ~n15146 & ~n13023;
  assign n13028 = ~n13025 & ~n13024;
  assign n13027 = ~n15602 | ~n13026;
  assign P2_U3161 = ~n13028 | ~n13027;
  assign n13033 = P2_REG1_REG_11__SCAN_IN ^ n13269;
  assign n13051 = ~n13033 & ~n15182;
  assign n13035 = ~n15398 | ~P2_ADDR_REG_11__SCAN_IN;
  assign n13034 = ~n13258 | ~n15396;
  assign n13036 = ~n13035 | ~n13034;
  assign n13049 = ~n13037 & ~n13036;
  assign n13042 = ~n13040;
  assign n13043 = ~n13042 | ~n13041;
  assign n13046 = ~n15386 | ~P2_REG2_REG_11__SCAN_IN;
  assign n13045 = ~n15388 | ~P2_REG1_REG_11__SCAN_IN;
  assign n13047 = n13256 ^ ~n13255;
  assign n13048 = ~n13047 | ~n15394;
  assign n13050 = ~n13049 | ~n13048;
  assign n13059 = ~n13051 & ~n13050;
  assign n13057 = P2_REG2_REG_11__SCAN_IN ^ ~n13277;
  assign n13058 = ~n15378 | ~n13057;
  assign P2_U3193 = ~n13059 | ~n13058;
  assign n13072 = P1_REG2_REG_12__SCAN_IN & n15323;
  assign n13070 = ~n15654 | ~n13060;
  assign n16181 = ~n13061 & ~n16274;
  assign n13062 = ~n15802 | ~n15803;
  assign n13140 = ~n13065 | ~n13064;
  assign n13068 = ~n13140 | ~n13066;
  assign n13187 = ~n13068 | ~n13067;
  assign n13098 = ~n13072 & ~n13071;
  assign n13075 = ~n13073 | ~n16177;
  assign n13074 = ~n16076;
  assign n13149 = ~n13075 | ~n13074;
  assign n13077 = ~n13149;
  assign n13079 = ~n13077 | ~n16088;
  assign n13195 = ~n13078 | ~n13079;
  assign n13083 = n13195 & n15637;
  assign n13081 = ~n13079 | ~n16270;
  assign n13080 = ~n16181;
  assign n13085 = ~n15840 & ~n14935;
  assign n13084 = ~n13283 & ~n15639;
  assign n13086 = ~n13085 & ~n13084;
  assign n13095 = ~n13245;
  assign n13090 = ~n15819 | ~n13143;
  assign n13091 = ~n13090 | ~n16367;
  assign n13246 = n13091 | n13202;
  assign n13093 = ~n13246 & ~n16322;
  assign n13092 = ~n15826 & ~n13221;
  assign n13094 = ~n13093 & ~n13092;
  assign n13096 = ~n13095 | ~n13094;
  assign n13097 = ~n13096 | ~n13226;
  assign P1_U3281 = ~n13098 | ~n13097;
  assign n13100 = ~P2_REG2_REG_10__SCAN_IN | ~n15240;
  assign n13099 = ~n16358 | ~n13419;
  assign n13107 = ~n13100 | ~n13099;
  assign n13105 = ~n13409 | ~n16424;
  assign n13330 = ~n13103 & ~n16582;
  assign n13104 = ~n13390 | ~n13233;
  assign n13106 = ~n13105 | ~n13104;
  assign n13118 = ~n13107 & ~n13106;
  assign n13108 = ~n13314 & ~n16866;
  assign n13318 = ~n13315 & ~n13410;
  assign n13109 = ~n13108 & ~n13318;
  assign n13110 = n13109 ^ ~n16868;
  assign n13114 = ~n13110 & ~n11752;
  assign n13112 = ~n13410 | ~n16345;
  assign n13111 = ~n16605 | ~n16346;
  assign n13113 = ~n13112 | ~n13111;
  assign n13116 = ~n13114 & ~n13113;
  assign n13117 = ~n13232 | ~n16419;
  assign P2_U3223 = ~n13118 | ~n13117;
  assign n16962 = ~n13119 & ~P2_U3151;
  assign n13121 = ~n13683 | ~P1_DATAO_REG_23__SCAN_IN;
  assign P2_U3272 = ~n13122 | ~n13121;
  assign n13126 = ~n14157 & ~n13125;
  assign P1_U3332 = ~n13128 | ~n16328;
  assign n13136 = ~P2_REG1_REG_9__SCAN_IN | ~n16444;
  assign n13130 = ~n13129 & ~n16433;
  assign n13134 = ~n13131 & ~n13130;
  assign n13133 = ~n13132 | ~n13731;
  assign n13135 = ~n16442 | ~n13137;
  assign P2_U3468 = ~n13136 | ~n13135;
  assign n13139 = ~P2_REG0_REG_9__SCAN_IN | ~n16439;
  assign n13138 = ~n16438 | ~n13137;
  assign P2_U3417 = ~n13139 | ~n13138;
  assign n13146 = ~n13170 & ~n13560;
  assign n13142 = ~n13517 | ~n13141;
  assign n13144 = n13142 & n16367;
  assign n13172 = ~n13144 | ~n13143;
  assign n13145 = ~n13172 & ~n16322;
  assign n13155 = ~n13146 & ~n13145;
  assign n13148 = n13170 | n11663;
  assign n13147 = ~n15820 | ~n15533;
  assign n13150 = n16179 ^ ~n13149;
  assign n13151 = ~n13503 | ~n15484;
  assign n13160 = ~n14874 & ~n13501;
  assign n13158 = ~n13517 | ~n15660;
  assign n13157 = ~n15323 | ~P1_REG2_REG_11__SCAN_IN;
  assign n13159 = ~n13158 | ~n13157;
  assign n13161 = ~n13160 & ~n13159;
  assign P1_U3282 = ~n13162 | ~n13161;
  assign n13164 = ~P2_DATAO_REG_28__SCAN_IN | ~n13429;
  assign P2_U3519 = ~n13164 | ~n13163;
  assign n13167 = ~n13165 & ~P1_U3086;
  assign n13166 = n13309 & P2_DATAO_REG_24__SCAN_IN;
  assign n13168 = ~n13167 & ~n13166;
  assign P1_U3331 = ~n13169 | ~n13168;
  assign n13178 = ~P1_REG0_REG_11__SCAN_IN | ~n16378;
  assign n13171 = ~n13517 | ~n16369;
  assign n13173 = ~n13172 | ~n13171;
  assign P1_U3486 = ~n13178 | ~n13177;
  assign n13181 = ~P1_REG1_REG_11__SCAN_IN | ~n16383;
  assign P1_U3533 = ~n13181 | ~n13180;
  assign n13185 = ~n13183 | ~n13182;
  assign ADD_1068_U55 = n13185 ^ ~n13184;
  assign n13209 = ~P1_REG1_REG_13__SCAN_IN | ~n16383;
  assign n13188 = ~n15819 | ~n15820;
  assign n13191 = ~n13189 | ~n13188;
  assign n13194 = ~n16274;
  assign n13549 = ~n13195 | ~n13194;
  assign n13198 = ~n13571 & ~n14935;
  assign n13197 = ~n15829 & ~n15639;
  assign n13199 = ~n13198 & ~n13197;
  assign n13201 = ~n15839 & ~n13202;
  assign n13203 = ~n13201 & ~n15534;
  assign n13220 = ~n13203 | ~n13541;
  assign n13204 = ~n15835 | ~n16369;
  assign n13205 = ~n13220 | ~n13204;
  assign P1_U3535 = ~n13209 | ~n13208;
  assign n13212 = ~P1_REG0_REG_13__SCAN_IN | ~n16378;
  assign P1_U3492 = ~n13212 | ~n13211;
  assign n13218 = ~n14874 & ~n13213;
  assign n13216 = ~P1_REG2_REG_13__SCAN_IN | ~n15323;
  assign n13229 = ~n13218 & ~n13217;
  assign n13225 = ~n13219;
  assign n13223 = ~n13220 & ~n16322;
  assign n13222 = ~n15839 & ~n13221;
  assign n13224 = ~n13223 & ~n13222;
  assign n13228 = ~n13227 | ~n13226;
  assign P1_U3280 = ~n13229 | ~n13228;
  assign n13237 = ~P2_REG0_REG_10__SCAN_IN | ~n16439;
  assign n13231 = ~n13230 & ~n16433;
  assign P2_U3420 = ~n13237 | ~n13236;
  assign n13240 = ~P2_REG1_REG_10__SCAN_IN | ~n16444;
  assign P2_U3469 = ~n13240 | ~n13239;
  assign n13249 = ~P1_REG0_REG_12__SCAN_IN | ~n16378;
  assign n13242 = ~n15819 | ~n16369;
  assign P1_U3489 = ~n13249 | ~n13248;
  assign n13252 = ~P1_REG1_REG_12__SCAN_IN | ~n16383;
  assign P1_U3534 = ~n13252 | ~n13251;
  assign n13254 = ~n15398 | ~P2_ADDR_REG_12__SCAN_IN;
  assign n13253 = ~n13779 | ~n15396;
  assign n13266 = ~n13254 | ~n13253;
  assign n13259 = ~n13257;
  assign n13260 = ~n13259 | ~n13258;
  assign n13263 = ~n15386 | ~P2_REG2_REG_12__SCAN_IN;
  assign n13262 = ~n15388 | ~P2_REG1_REG_12__SCAN_IN;
  assign n13777 = ~n13263 | ~n13262;
  assign n13264 = n13776 ^ n13775;
  assign n13265 = ~n13264 & ~n15268;
  assign n13267 = ~n13266 & ~n13265;
  assign n13342 = ~P2_REG3_REG_12__SCAN_IN | ~P2_U3151;
  assign n13274 = ~n13267 | ~n13342;
  assign n13766 = ~n13271 | ~n13270;
  assign n13272 = n13766 ^ n13767;
  assign n13273 = ~n13272 & ~n15182;
  assign n13282 = ~n13274 & ~n13273;
  assign n13790 = ~n13279 | ~n13278;
  assign n13280 = n13791 ^ ~n13790;
  assign n13281 = ~n13280 | ~n15378;
  assign P2_U3194 = ~n13282 | ~n13281;
  assign n13285 = ~n15515 & ~n13283;
  assign n13287 = ~n13285 & ~n13284;
  assign n13286 = ~n15521 | ~n15789;
  assign n13297 = ~n13287 | ~n13286;
  assign n13291 = ~n13289 | ~n13288;
  assign n13294 = ~n13293 | ~n15428;
  assign n13299 = ~n13298 | ~n15516;
  assign P1_U3217 = ~n13300 | ~n13299;
  assign n13304 = ~n13303 & ~P2_U3151;
  assign n13306 = ~n13683 | ~P1_DATAO_REG_24__SCAN_IN;
  assign P2_U3271 = ~n13307 | ~n13306;
  assign n13311 = ~n13308 & ~P1_U3086;
  assign n13310 = n13309 & P2_DATAO_REG_25__SCAN_IN;
  assign n13312 = ~n13311 & ~n13310;
  assign P1_U3330 = ~n13313 | ~n13312;
  assign n13338 = ~P2_REG0_REG_11__SCAN_IN | ~n16439;
  assign n13317 = ~n13314;
  assign n13316 = ~n13315 | ~n13410;
  assign n13321 = ~n13317 | ~n13316;
  assign n13319 = ~n13409 & ~n13325;
  assign n13323 = ~n13321 | ~n13320;
  assign n13377 = ~n13323 | ~n13322;
  assign n13324 = n16870 ^ n13377;
  assign n13329 = ~n13324 & ~n11752;
  assign n13327 = ~n13325 | ~n16345;
  assign n13326 = ~n16466 | ~n16346;
  assign n13328 = ~n13327 | ~n13326;
  assign n13361 = ~n13330 | ~n16592;
  assign n13331 = ~n13361 | ~n16586;
  assign n13334 = ~n16610 | ~n14685;
  assign n13339 = n13387 | n13336;
  assign P2_U3423 = ~n13338 | ~n13337;
  assign n13341 = ~P2_REG1_REG_11__SCAN_IN | ~n16444;
  assign P2_U3470 = ~n13341 | ~n13340;
  assign n13345 = ~n15603 & ~n16608;
  assign n13343 = ~n15604 | ~n13859;
  assign n13344 = ~n13343 | ~n13342;
  assign n13355 = ~n13345 & ~n13344;
  assign n13347 = n13346 ^ ~n16466;
  assign n13351 = ~n15602 | ~n13356;
  assign n13350 = ~n13635 | ~n15342;
  assign n13352 = ~n13351 | ~n13350;
  assign P2_U3164 = ~n13355 | ~n13354;
  assign n13358 = ~n15240 | ~P2_REG2_REG_12__SCAN_IN;
  assign n13357 = ~n16358 | ~n13356;
  assign n13371 = ~n13358 | ~n13357;
  assign n13359 = ~n16586;
  assign n13363 = ~n13361 | ~n16597;
  assign n13365 = ~n13363 | ~n13362;
  assign n13636 = ~n13365 | ~n13380;
  assign n13366 = ~n13365 & ~n13380;
  assign n13369 = n13442 | n16423;
  assign n13368 = ~n13635 | ~n16424;
  assign n13385 = ~n13371 & ~n13370;
  assign n13373 = ~n16605 | ~n16345;
  assign n13372 = ~n13859 | ~n16346;
  assign n13374 = ~n13373 | ~n13372;
  assign n13379 = ~n13377 & ~n13376;
  assign n13647 = ~n13379 & ~n13378;
  assign n13384 = ~n13441 | ~n16419;
  assign P2_U3221 = ~n13385 | ~n13384;
  assign n13386 = ~n16607 & ~n15564;
  assign n13388 = ~n13387 & ~n13386;
  assign n13394 = ~n15240 & ~n13388;
  assign n13392 = ~P2_REG2_REG_11__SCAN_IN | ~n15240;
  assign n13391 = ~n13390 | ~n13389;
  assign n13396 = ~n16358 | ~n13395;
  assign P2_U3222 = ~n13397 | ~n13396;
  assign n13405 = ~P2_DATAO_REG_30__SCAN_IN | ~n13429;
  assign n13399 = ~n13430 | ~P2_REG0_REG_30__SCAN_IN;
  assign n13398 = ~n13431 | ~P2_REG1_REG_30__SCAN_IN;
  assign n13403 = n13399 & n13398;
  assign n13436 = ~n8930 | ~n14429;
  assign n13401 = ~n13434 | ~P2_REG2_REG_30__SCAN_IN;
  assign n13404 = ~P2_U3893 | ~n16905;
  assign P2_U3521 = ~n13405 | ~n13404;
  assign n13408 = n13407 ^ n13406;
  assign n13414 = ~n13408 & ~n15617;
  assign n13412 = ~n13409 | ~n15342;
  assign n13411 = ~n15355 | ~n13410;
  assign n13413 = ~n13412 | ~n13411;
  assign n13416 = ~n13414 & ~n13413;
  assign n13417 = ~n15146 & ~n16608;
  assign n13421 = ~n13418 & ~n13417;
  assign n13420 = ~n15602 | ~n13419;
  assign P2_U3157 = ~n13421 | ~n13420;
  assign n13428 = ~P2_DATAO_REG_29__SCAN_IN | ~n13429;
  assign n13423 = ~n13431 | ~P2_REG1_REG_29__SCAN_IN;
  assign n13422 = ~n13430 | ~P2_REG0_REG_29__SCAN_IN;
  assign n13426 = n13423 & n13422;
  assign n13424 = ~n13434 | ~P2_REG2_REG_29__SCAN_IN;
  assign n16801 = ~n13426 | ~n13425;
  assign n13427 = ~P2_U3893 | ~n16801;
  assign P2_U3520 = ~n13428 | ~n13427;
  assign n13440 = ~P2_DATAO_REG_31__SCAN_IN | ~n13429;
  assign n13433 = ~n13430 | ~P2_REG0_REG_31__SCAN_IN;
  assign n13432 = ~n13431 | ~P2_REG1_REG_31__SCAN_IN;
  assign n13438 = n13433 & n13432;
  assign n13435 = ~n13434 | ~P2_REG2_REG_31__SCAN_IN;
  assign n16933 = ~n13438 | ~n13437;
  assign n13439 = ~P2_U3893 | ~n16933;
  assign P2_U3522 = ~n13440 | ~n13439;
  assign n13448 = ~P2_REG0_REG_12__SCAN_IN | ~n16439;
  assign n13443 = ~n16467 & ~n16433;
  assign P2_U3426 = ~n13448 | ~n13447;
  assign n13451 = ~P2_REG1_REG_12__SCAN_IN | ~n16444;
  assign P2_U3471 = ~n13451 | ~n13450;
  assign n13455 = ~n13454 & ~P2_U3151;
  assign n13457 = ~n13683 | ~P1_DATAO_REG_25__SCAN_IN;
  assign P2_U3270 = ~n13458 | ~n13457;
  assign n13463 = ~n13460 & ~P1_U3086;
  assign n13462 = ~n14157 & ~n13461;
  assign n13464 = ~n13463 & ~n13462;
  assign P1_U3329 = ~n13465 | ~n13464;
  assign n13467 = n13466 ^ ~n13859;
  assign n13475 = ~n13714 | ~n15342;
  assign n13471 = ~n15146 & ~n13730;
  assign n13774 = ~P2_STATE_REG_SCAN_IN & ~n13470;
  assign n13473 = n13471 | n13774;
  assign n13472 = ~n15603 & ~n13634;
  assign n13474 = ~n13473 & ~n13472;
  assign n13476 = ~n13475 | ~n13474;
  assign n13478 = ~n13653 | ~n15602;
  assign P2_U3174 = ~n13479 | ~n13478;
  assign n13498 = ~n14450 & ~n13490;
  assign n13486 = ~n13484 & ~P1_REG2_REG_15__SCAN_IN;
  assign n13485 = ~n15137 | ~n13833;
  assign n13495 = ~n13486 & ~n13485;
  assign n13489 = ~n13487 | ~P1_REG1_REG_14__SCAN_IN;
  assign n13493 = ~n13491 & ~P1_REG1_REG_15__SCAN_IN;
  assign n13492 = ~n13841 | ~n8934;
  assign n13494 = ~n13493 & ~n13492;
  assign n13496 = ~n13495 & ~n13494;
  assign n14114 = ~P1_REG3_REG_15__SCAN_IN | ~P1_U3086;
  assign n13500 = ~n13498 & ~n13497;
  assign n13499 = ~n15122 | ~P1_ADDR_REG_15__SCAN_IN;
  assign P1_U3258 = ~n13500 | ~n13499;
  assign n13516 = ~n13502 & ~n13501;
  assign n13505 = ~n15521 | ~n13503;
  assign n13507 = ~n13505 | ~n13504;
  assign n13506 = ~n15515 & ~n15829;
  assign n13514 = ~n13507 & ~n13506;
  assign n13510 = n13509 ^ ~n13508;
  assign n13518 = ~n13517 | ~n15428;
  assign P1_U3236 = ~n13519 | ~n13518;
  assign n13535 = ~n15516 | ~n13520;
  assign n13531 = ~n15835 | ~n15428;
  assign n13527 = ~n15439 | ~n15850;
  assign n13529 = ~n13527 | ~n13526;
  assign n13528 = ~n15094 & ~n15829;
  assign n13530 = ~n13529 & ~n13528;
  assign n13532 = ~n13531 | ~n13530;
  assign P1_U3234 = ~n13535 | ~n13534;
  assign n13538 = ~n15323 | ~P1_REG2_REG_14__SCAN_IN;
  assign n13537 = ~n13536 | ~n15654;
  assign n13540 = ~n13538 | ~n13537;
  assign n13539 = ~n13604 & ~n15497;
  assign n13566 = ~n13540 & ~n13539;
  assign n13543 = ~n13581;
  assign n13542 = ~n15849 | ~n13541;
  assign n13564 = ~n13603 & ~n15074;
  assign n16185 = ~n13545 & ~n13544;
  assign n13567 = ~n13547 & ~n13546;
  assign n13551 = ~n13550 | ~n16061;
  assign n13569 = ~n13551 | ~n16185;
  assign n13555 = ~n13694 & ~n14935;
  assign n13554 = ~n15840 & ~n15639;
  assign n13556 = ~n13555 & ~n13554;
  assign n13608 = n13559 | n13558;
  assign P1_U3279 = ~n13566 | ~n13565;
  assign n16187 = ~n16282 | ~n16060;
  assign n13687 = ~n13568 | ~n15853;
  assign n13691 = ~n13569 | ~n16062;
  assign n13572 = ~n13571 & ~n15639;
  assign n13576 = ~n15654 | ~n14112;
  assign n13577 = ~n13226 | ~n13576;
  assign n13578 = ~n13226 & ~P1_REG2_REG_15__SCAN_IN;
  assign n13590 = n13579 | n13578;
  assign n13582 = ~n13619 & ~n13581;
  assign n13586 = ~n13618 | ~n15659;
  assign n13584 = ~n13619 & ~n15497;
  assign n13583 = ~n15502 & ~n14116;
  assign n13585 = ~n13584 & ~n13583;
  assign n13587 = ~n13586 | ~n13585;
  assign P1_U3278 = ~n13590 | ~n13589;
  assign n13593 = ~n15603 & ~n16462;
  assign n13591 = ~n15604 | ~n16645;
  assign n14024 = ~P2_REG3_REG_14__SCAN_IN | ~P2_U3151;
  assign n13592 = ~n13591 | ~n14024;
  assign n13602 = ~n13593 & ~n13592;
  assign n13598 = ~n15602 | ~n13869;
  assign n13597 = ~n16628 | ~n15342;
  assign n13599 = ~n13598 | ~n13597;
  assign P2_U3155 = ~n13602 | ~n13601;
  assign n13613 = ~P1_REG1_REG_14__SCAN_IN | ~n16383;
  assign n13606 = ~n13603 & ~n15534;
  assign n13605 = ~n13604 & ~n15536;
  assign P1_U3536 = ~n13613 | ~n13612;
  assign n13616 = ~P1_REG0_REG_14__SCAN_IN | ~n16378;
  assign P1_U3495 = ~n13616 | ~n13615;
  assign n13630 = ~P1_REG1_REG_15__SCAN_IN | ~n16383;
  assign n13623 = ~n13618 | ~n16367;
  assign n13621 = ~n13619 & ~n15536;
  assign n13620 = ~n14116 & ~n14935;
  assign n13622 = ~n13621 & ~n13620;
  assign P1_U3537 = ~n13630 | ~n13629;
  assign n13633 = ~P1_REG0_REG_15__SCAN_IN | ~n16378;
  assign P1_U3498 = ~n13633 | ~n13632;
  assign n13638 = ~n13636 | ~n16604;
  assign n16874 = ~n13637 & ~n13727;
  assign n13729 = ~n13638 | ~n16874;
  assign n13640 = ~n13729;
  assign n13639 = ~n13638 & ~n16874;
  assign n13659 = ~n13664 & ~n16423;
  assign n13642 = ~n16631 | ~n16346;
  assign n13641 = ~n16466 | ~n16345;
  assign n13643 = ~n13642 | ~n13641;
  assign n13649 = ~n13647 | ~n13646;
  assign n13716 = ~n13649 | ~n13648;
  assign n13655 = ~n16358 | ~n13653;
  assign n13662 = ~n16461 & ~n16433;
  assign n13654 = ~n13662 | ~n13871;
  assign n13656 = ~n13655 | ~n13654;
  assign n13660 = ~n15240 | ~P2_REG2_REG_13__SCAN_IN;
  assign P2_U3220 = ~n13661 | ~n13660;
  assign n13668 = ~P2_REG0_REG_13__SCAN_IN | ~n16439;
  assign n13665 = n13664 | n16431;
  assign P2_U3429 = ~n13668 | ~n13667;
  assign n13671 = ~P2_REG1_REG_13__SCAN_IN | ~n16444;
  assign P2_U3472 = ~n13671 | ~n13670;
  assign n13676 = ~n13673 & ~P1_U3086;
  assign n13675 = ~n14157 & ~n13674;
  assign n13677 = ~n13676 & ~n13675;
  assign P1_U3328 = ~n13678 | ~n13677;
  assign n13681 = ~n15388 & ~P2_U3151;
  assign n13684 = ~n13683 | ~P1_DATAO_REG_27__SCAN_IN;
  assign P2_U3268 = ~n13685 | ~n13684;
  assign n13689 = ~n13687 & ~n13690;
  assign n13799 = ~n13689 & ~n13688;
  assign n13806 = ~n13692 | ~n16282;
  assign n13696 = ~n15885 & ~n14935;
  assign n13695 = ~n13694 & ~n15639;
  assign n13697 = ~n13696 & ~n13695;
  assign n13701 = ~P1_REG2_REG_16__SCAN_IN;
  assign n13702 = ~n15323 | ~n13701;
  assign n13705 = ~n13797 & ~n13704;
  assign n13709 = ~n13754 | ~n15659;
  assign n13707 = ~n13797 & ~n15497;
  assign n13706 = n15654 & n14134;
  assign n13708 = ~n13707 & ~n13706;
  assign n13710 = ~n13709 | ~n13708;
  assign P1_U3277 = ~n13713 | ~n13712;
  assign n13864 = ~n13718 | ~n13717;
  assign n13721 = ~n13864 | ~n13719;
  assign n13951 = ~n13721 | ~n13720;
  assign n13724 = ~n14079 | ~n16346;
  assign n13723 = ~n16631 | ~n16345;
  assign n13725 = ~n13724 | ~n13723;
  assign n13856 = ~n13729 | ~n13728;
  assign n16456 = ~n16628 | ~n13730;
  assign n13855 = ~n13856 | ~n13865;
  assign n13959 = ~n13855 | ~n16456;
  assign n16386 = ~n16410 & ~n13731;
  assign n13732 = ~n16637 & ~n16433;
  assign n13735 = ~n16444 | ~P2_REG1_REG_15__SCAN_IN;
  assign P2_U3474 = ~n13736 | ~n13735;
  assign n13738 = ~n16439 | ~P2_REG0_REG_15__SCAN_IN;
  assign P2_U3435 = ~n13739 | ~n13738;
  assign n13742 = ~n15240 | ~n13741;
  assign n13748 = ~n16642 | ~n16424;
  assign n13747 = ~n16358 | ~n13746;
  assign n13749 = ~n13748 | ~n13747;
  assign P2_U3218 = ~n13752 | ~n13751;
  assign n13755 = ~n14135 | ~n16369;
  assign n13761 = ~n16383 | ~P1_REG1_REG_16__SCAN_IN;
  assign P1_U3538 = ~n13762 | ~n13761;
  assign n13764 = ~n16378 | ~P1_REG0_REG_16__SCAN_IN;
  assign P1_U3501 = ~n13765 | ~n13764;
  assign n14026 = ~n13769 | ~n13768;
  assign n13770 = P2_REG1_REG_13__SCAN_IN ^ n14027;
  assign n13788 = ~n13770 & ~n15182;
  assign n13772 = ~n15398 | ~P2_ADDR_REG_13__SCAN_IN;
  assign n13771 = ~n14015 | ~n15396;
  assign n13773 = ~n13772 | ~n13771;
  assign n13786 = ~n13774 & ~n13773;
  assign n13778 = ~n13777;
  assign n13780 = ~n13779 | ~n13778;
  assign n13783 = ~n15386 | ~P2_REG2_REG_13__SCAN_IN;
  assign n13782 = ~n15388 | ~P2_REG1_REG_13__SCAN_IN;
  assign n13784 = n14013 ^ ~n14012;
  assign n13785 = ~n13784 | ~n15394;
  assign n13787 = ~n13786 | ~n13785;
  assign n14033 = ~n13793 | ~n13792;
  assign n13794 = P2_REG2_REG_13__SCAN_IN ^ ~n14035;
  assign n13795 = ~n15378 | ~n13794;
  assign P2_U3195 = ~n13796 | ~n13795;
  assign n16229 = ~n14178 & ~n15883;
  assign n16230 = ~n15880 & ~n14177;
  assign n14185 = ~n16229 & ~n16230;
  assign n13911 = ~n13801 | ~n13800;
  assign n14180 = ~n13804 | ~n13803;
  assign n13807 = ~n13806 & ~n13805;
  assign n13913 = ~n13807 & ~n16056;
  assign n13916 = ~n13913 | ~n13912;
  assign n14186 = ~n13916 | ~n15887;
  assign n13812 = ~n14610 & ~n14935;
  assign n13811 = ~n15885 & ~n15639;
  assign n13813 = ~n13812 & ~n13811;
  assign n13815 = ~n13226 & ~P1_REG2_REG_18__SCAN_IN;
  assign n13818 = n15880 & n13927;
  assign n14212 = ~n15880 & ~n13927;
  assign n13823 = ~n13985 | ~n15659;
  assign n13821 = ~n14178 & ~n15497;
  assign n13820 = n15654 & n13819;
  assign n13822 = ~n13821 & ~n13820;
  assign P1_U3275 = ~n13827 | ~n13826;
  assign n13831 = ~n14450 & ~n13828;
  assign n13829 = ~n15122 | ~P1_ADDR_REG_16__SCAN_IN;
  assign n14137 = ~P1_REG3_REG_16__SCAN_IN | ~P1_U3086;
  assign n13830 = ~n13829 | ~n14137;
  assign n13850 = ~n13831 & ~n13830;
  assign n13836 = P1_REG2_REG_16__SCAN_IN ^ n14457;
  assign n13838 = ~n13836 & ~n13835;
  assign n13837 = ~n15137 | ~n14451;
  assign n13848 = ~n13838 & ~n13837;
  assign n13844 = P1_REG1_REG_16__SCAN_IN ^ n14457;
  assign n13846 = ~n13844 & ~n13843;
  assign n13845 = ~n14458 | ~n8934;
  assign n13847 = ~n13846 & ~n13845;
  assign n13849 = ~n13848 & ~n13847;
  assign P1_U3259 = ~n13850 | ~n13849;
  assign n13852 = ~n16958 & ~P2_U3151;
  assign n15586 = ~P1_DATAO_REG_28__SCAN_IN;
  assign n13851 = ~n14356 & ~n15586;
  assign n13853 = ~n13852 & ~n13851;
  assign P2_U3267 = ~n13854 | ~n13853;
  assign n13858 = ~n13855;
  assign n13857 = ~n13856 & ~n13865;
  assign n13861 = ~n16645 | ~n16346;
  assign n13860 = ~n13859 | ~n16345;
  assign n13862 = ~n13861 | ~n13860;
  assign n13873 = ~n16358 | ~n13869;
  assign n13872 = ~n13887 | ~n13871;
  assign n13874 = ~n13873 | ~n13872;
  assign n13878 = ~n15240 | ~P2_REG2_REG_14__SCAN_IN;
  assign P2_U3219 = ~n13879 | ~n13878;
  assign n13884 = ~n13881 & ~P1_U3086;
  assign n13883 = ~n14157 & ~n13882;
  assign n13885 = ~n13884 & ~n13883;
  assign P1_U3327 = ~n13886 | ~n13885;
  assign n13893 = ~P2_REG0_REG_14__SCAN_IN | ~n16439;
  assign n13890 = n13889 | n16431;
  assign P2_U3432 = ~n13893 | ~n13892;
  assign n13896 = ~P2_REG1_REG_14__SCAN_IN | ~n16444;
  assign P2_U3473 = ~n13896 | ~n13895;
  assign n13899 = ~n13898 & ~n13897;
  assign n13908 = n15602 & n13977;
  assign n13904 = ~n14075 & ~n15601;
  assign n13902 = ~n15355 | ~n16645;
  assign n14707 = ~P2_REG3_REG_16__SCAN_IN | ~P2_U3151;
  assign n13903 = ~n13902 | ~n14707;
  assign n13906 = ~n13904 & ~n13903;
  assign n13905 = ~n16665 | ~n15604;
  assign n13907 = ~n13906 | ~n13905;
  assign n13909 = ~n13908 & ~n13907;
  assign P2_U3166 = ~n13910 | ~n13909;
  assign n13918 = ~n14116 & ~n15639;
  assign n13917 = ~n14177 & ~n14935;
  assign n13919 = ~n13918 & ~n13917;
  assign n13923 = ~P1_REG2_REG_17__SCAN_IN;
  assign n13924 = ~n15323 | ~n13923;
  assign n13928 = ~n14059 | ~n13926;
  assign n13932 = ~n13938 | ~n15659;
  assign n13930 = ~n15888 & ~n15497;
  assign n13929 = n15654 & n14058;
  assign n13931 = ~n13930 & ~n13929;
  assign P1_U3276 = ~n13936 | ~n13935;
  assign n13945 = ~n16378 | ~P1_REG0_REG_17__SCAN_IN;
  assign P1_U3504 = ~n13946 | ~n13945;
  assign n13948 = ~n16383 | ~P1_REG1_REG_17__SCAN_IN;
  assign P1_U3539 = ~n13949 | ~n13948;
  assign n16650 = ~n14071 | ~n14074;
  assign n16651 = ~n14075 | ~n14079;
  assign n13953 = ~n13951 | ~n13950;
  assign n14070 = ~n13953 | ~n13952;
  assign n13956 = ~n16669 & ~n15559;
  assign n13955 = ~n13960 & ~n16411;
  assign n13957 = ~n13956 & ~n13955;
  assign n13961 = ~n13959 | ~n16878;
  assign n14084 = ~n13961 | ~n16636;
  assign n13964 = ~n14075 & ~n16433;
  assign n13967 = ~n16444 | ~P2_REG1_REG_16__SCAN_IN;
  assign P2_U3475 = ~n13968 | ~n13967;
  assign n13970 = ~n16439 | ~P2_REG0_REG_16__SCAN_IN;
  assign P2_U3438 = ~n13971 | ~n13970;
  assign n13975 = ~n13972 | ~n16419;
  assign n13974 = ~n15240 | ~n13973;
  assign n13979 = ~n14071 | ~n16424;
  assign n13978 = ~n13977 | ~n16358;
  assign n13980 = ~n13979 | ~n13978;
  assign P2_U3217 = ~n13983 | ~n13982;
  assign n13992 = ~n16383 | ~P1_REG1_REG_18__SCAN_IN;
  assign P1_U3540 = ~n13993 | ~n13992;
  assign n13995 = ~n16378 | ~P1_REG0_REG_18__SCAN_IN;
  assign P1_U3507 = ~n13996 | ~n13995;
  assign n14002 = ~n13999 & ~P2_U3151;
  assign n14001 = ~n14356 & ~n14000;
  assign n14003 = ~n14002 & ~n14001;
  assign P2_U3266 = ~n14004 | ~n14003;
  assign n14007 = ~n14005 & ~P1_U3086;
  assign n14895 = ~P2_DATAO_REG_29__SCAN_IN;
  assign n14006 = ~n14157 & ~n14895;
  assign n14008 = ~n14007 & ~n14006;
  assign P1_U3326 = ~n14009 | ~n14008;
  assign n14011 = ~n15398 | ~P2_ADDR_REG_14__SCAN_IN;
  assign n14010 = ~n14587 | ~n15396;
  assign n14023 = ~n14011 | ~n14010;
  assign n14016 = ~n14014;
  assign n14017 = ~n14016 | ~n14015;
  assign n14020 = ~n15386 | ~P2_REG2_REG_14__SCAN_IN;
  assign n14019 = ~n15388 | ~P2_REG1_REG_14__SCAN_IN;
  assign n14586 = ~n14020 | ~n14019;
  assign n14021 = n14585 ^ n14584;
  assign n14022 = ~n14021 & ~n15268;
  assign n14025 = ~n14023 & ~n14022;
  assign n14575 = ~n14029 | ~n14028;
  assign n14030 = n14575 ^ n14576;
  assign n14031 = ~n14030 & ~n15182;
  assign n14599 = ~n14037 | ~n14036;
  assign n14038 = n14600 ^ ~n14599;
  assign P2_U3196 = ~n14040 | ~n14039;
  assign n14046 = ~n15355 | ~n14079;
  assign n14045 = ~n15604 | ~n16680;
  assign n14052 = ~n14046 | ~n14045;
  assign n14050 = ~n15602 | ~n14101;
  assign n14048 = ~n16658 & ~n15601;
  assign n15188 = ~P2_STATE_REG_SCAN_IN & ~n14047;
  assign n14049 = ~n14048 & ~n15188;
  assign n14051 = ~n14050 | ~n14049;
  assign n14053 = ~n14052 & ~n14051;
  assign P2_U3168 = ~n14054 | ~n14053;
  assign n14067 = n15516 & n14058;
  assign n14065 = ~n14059 | ~n15428;
  assign n14061 = ~n15521 | ~n14060;
  assign n14466 = ~P1_REG3_REG_17__SCAN_IN | ~P1_U3086;
  assign n14063 = ~n14061 | ~n14466;
  assign n14062 = ~n15515 & ~n14177;
  assign n14064 = ~n14063 & ~n14062;
  assign n14066 = ~n14065 | ~n14064;
  assign n14068 = ~n14067 & ~n14066;
  assign P1_U3228 = ~n14069 | ~n14068;
  assign n14073 = ~n14070;
  assign n14077 = ~n14073 | ~n14072;
  assign n14274 = ~n14077 | ~n14076;
  assign n14081 = ~n16680 | ~n16346;
  assign n14080 = ~n14079 | ~n16345;
  assign n14082 = ~n14081 | ~n14080;
  assign n14085 = ~n14084 & ~n16666;
  assign n14283 = ~n14374 | ~n16882;
  assign n14086 = ~n14374 & ~n16882;
  assign n14091 = ~n16439 | ~P2_REG0_REG_17__SCAN_IN;
  assign P2_U3441 = ~n14092 | ~n14091;
  assign n14094 = ~n16444 | ~P2_REG1_REG_17__SCAN_IN;
  assign P2_U3476 = ~n14095 | ~n14094;
  assign n14099 = ~n14096 | ~n16419;
  assign n14097 = ~P2_REG2_REG_17__SCAN_IN;
  assign n14098 = ~n15240 | ~n14097;
  assign n14103 = ~n16659 | ~n16424;
  assign n14102 = ~n14101 | ~n16358;
  assign n14104 = ~n14103 | ~n14102;
  assign P2_U3216 = ~n14107 | ~n14106;
  assign n14127 = n14109 & n14108;
  assign n14126 = ~n14109 & ~n14108;
  assign n14122 = n15516 & n14112;
  assign n14120 = ~n14113 | ~n15428;
  assign n14115 = ~n15521 | ~n15850;
  assign n14118 = ~n14115 | ~n14114;
  assign n14117 = ~n15515 & ~n14116;
  assign n14119 = ~n14118 & ~n14117;
  assign n14121 = ~n14120 | ~n14119;
  assign n14123 = ~n14122 & ~n14121;
  assign P1_U3241 = ~n14124 | ~n14123;
  assign n14144 = n15516 & n14134;
  assign n14142 = ~n14135 | ~n15428;
  assign n14138 = ~n15521 | ~n14136;
  assign n14140 = ~n14138 | ~n14137;
  assign n14139 = ~n15515 & ~n15885;
  assign n14141 = ~n14140 & ~n14139;
  assign n14143 = ~n14142 | ~n14141;
  assign n14145 = ~n14144 & ~n14143;
  assign P1_U3226 = ~n14146 | ~n14145;
  assign n14151 = ~n14149 & ~P2_U3151;
  assign n14423 = ~P1_DATAO_REG_30__SCAN_IN;
  assign n14150 = ~n14356 & ~n14423;
  assign n14152 = ~n14151 & ~n14150;
  assign P2_U3265 = ~n14153 | ~n14152;
  assign n14159 = ~n14156 & ~P1_U3086;
  assign n14891 = ~P2_DATAO_REG_30__SCAN_IN;
  assign n14158 = ~n14157 & ~n14891;
  assign n14160 = ~n14159 & ~n14158;
  assign P1_U3325 = ~n14161 | ~n14160;
  assign n14166 = ~n14300;
  assign n14174 = ~n14167 & ~n14166;
  assign n14170 = ~n16675 & ~n15601;
  assign n14168 = ~n16665 | ~n15355;
  assign n15274 = ~P2_U3151 | ~P2_REG3_REG_18__SCAN_IN;
  assign n14169 = ~n14168 | ~n15274;
  assign n14172 = ~n14170 & ~n14169;
  assign n14171 = ~n14492 | ~n15604;
  assign P2_U3178 = ~n14176 | ~n14175;
  assign n14228 = ~n14182 | ~n14181;
  assign n16192 = ~n16289 & ~n16291;
  assign n14183 = n14228 | n16192;
  assign n14188 = ~n14186 | ~n14185;
  assign n14206 = ~n14188 | ~n16099;
  assign n14189 = ~n14206 | ~n16192;
  assign n14236 = ~n14189 | ~n15908;
  assign n14191 = ~n15901 | ~n15484;
  assign n14193 = ~n13226 & ~P1_REG2_REG_20__SCAN_IN;
  assign n14214 = n15902 & n14212;
  assign n14243 = n14337 & n14214;
  assign n14199 = ~n14337 & ~n15497;
  assign n14197 = ~n14609 | ~n15654;
  assign n14196 = ~n15083 | ~n14611;
  assign n14198 = ~n14197 | ~n14196;
  assign n14200 = ~n14199 & ~n14198;
  assign P1_U3273 = ~n14205 | ~n14204;
  assign n14208 = ~n15883 | ~n15484;
  assign n14216 = ~n15902 & ~n15536;
  assign n14215 = ~n14737 & ~n14935;
  assign n14217 = ~n14216 & ~n14215;
  assign n14222 = ~n16378 | ~P1_REG0_REG_19__SCAN_IN;
  assign P1_U3509 = ~n14223 | ~n14222;
  assign n14225 = ~n16383 | ~P1_REG1_REG_19__SCAN_IN;
  assign P1_U3541 = ~n14226 | ~n14225;
  assign n16106 = ~n14736 & ~n14914;
  assign n16196 = ~n15927 & ~n16106;
  assign n14234 = ~n14232 | ~n14231;
  assign n14399 = ~n14234 | ~n14233;
  assign n14403 = ~n14236 | ~n14235;
  assign n14240 = ~n15916 | ~n15484;
  assign n14245 = n14311 | n16322;
  assign n14247 = ~n13226 & ~P1_REG2_REG_21__SCAN_IN;
  assign n14250 = ~n15502 & ~n15937;
  assign n14249 = n15654 & n14735;
  assign n14251 = ~n14250 & ~n14249;
  assign P1_U3272 = ~n14256 | ~n14255;
  assign n14258 = n13226 | P1_REG2_REG_19__SCAN_IN;
  assign n14264 = ~n14262 | ~n15660;
  assign n14263 = ~n14439 | ~n15654;
  assign n14266 = ~n14264 | ~n14263;
  assign n14265 = ~n14737 & ~n15502;
  assign n14267 = ~n14266 & ~n14265;
  assign P1_U3274 = ~n14272 | ~n14271;
  assign n14276 = ~n14274 | ~n14273;
  assign n14362 = ~n14276 | ~n14275;
  assign n14279 = ~n16696 & ~n15559;
  assign n14278 = ~n16669 & ~n16411;
  assign n14280 = ~n14279 & ~n14278;
  assign n14290 = ~n16444 | ~P2_REG1_REG_18__SCAN_IN;
  assign P2_U3477 = ~n14291 | ~n14290;
  assign n14293 = ~n16439 | ~P2_REG0_REG_18__SCAN_IN;
  assign P2_U3444 = ~n14294 | ~n14293;
  assign n14297 = ~n15240 | ~n14296;
  assign n14302 = ~n16679 | ~n16424;
  assign n14301 = ~n14300 | ~n16358;
  assign n14303 = ~n14302 | ~n14301;
  assign P2_U3215 = ~n14306 | ~n14305;
  assign n14308 = ~n15937 & ~n14935;
  assign n14316 = ~n16378 | ~P1_REG0_REG_21__SCAN_IN;
  assign P1_U3511 = ~n14317 | ~n14316;
  assign n14319 = ~n16383 | ~P1_REG1_REG_21__SCAN_IN;
  assign P1_U3543 = ~n14320 | ~n14319;
  assign n14326 = ~n15355 | ~n16680;
  assign n14325 = ~n15604 | ~n14641;
  assign n14332 = ~n14326 | ~n14325;
  assign n14330 = ~n15602 | ~n14381;
  assign n14328 = ~n16695 & ~n15601;
  assign n15399 = ~P2_U3151 | ~P2_REG3_REG_19__SCAN_IN;
  assign n14327 = ~n15399;
  assign n14329 = ~n14328 & ~n14327;
  assign P2_U3159 = ~n14334 | ~n14333;
  assign n14339 = ~n14337 & ~n15536;
  assign n14338 = ~n14914 & ~n14935;
  assign n14346 = ~n16383 | ~P1_REG1_REG_20__SCAN_IN;
  assign P1_U3542 = ~n14347 | ~n14346;
  assign n14349 = ~n16378 | ~P1_REG0_REG_20__SCAN_IN;
  assign P1_U3510 = ~n14350 | ~n14349;
  assign n14353 = ~P2_IR_REG_30__SCAN_IN & ~P2_U3151;
  assign n14354 = ~P2_IR_REG_31__SCAN_IN | ~n14353;
  assign n14358 = ~n14355 & ~n14354;
  assign n14568 = ~P1_DATAO_REG_31__SCAN_IN;
  assign n14357 = ~n14356 & ~n14568;
  assign n14359 = ~n14358 & ~n14357;
  assign P2_U3264 = ~n14360 | ~n14359;
  assign n14364 = ~n14362 | ~n14361;
  assign n14488 = ~n14364 | ~n14363;
  assign n14367 = ~n14641 | ~n16346;
  assign n14366 = ~n16680 | ~n16345;
  assign n14368 = ~n14367 | ~n14366;
  assign n14370 = n16419 | P2_REG2_REG_19__SCAN_IN;
  assign n14380 = ~n14374 | ~n14373;
  assign n14494 = ~n14380 | ~n14379;
  assign n14383 = ~n14495 | ~n16424;
  assign n14382 = ~n14381 | ~n16358;
  assign P2_U3214 = ~n14387 | ~n14386;
  assign n14393 = ~n16444 | ~P2_REG1_REG_19__SCAN_IN;
  assign P2_U3478 = ~n14394 | ~n14393;
  assign n14396 = ~n16439 | ~P2_REG0_REG_19__SCAN_IN;
  assign P2_U3446 = ~n14397 | ~n14396;
  assign n16198 = ~n16294 | ~n14398;
  assign n14548 = ~n14404 | ~n16109;
  assign n14407 = ~n15953 & ~n14935;
  assign n14406 = ~n14914 & ~n15639;
  assign n14408 = ~n14407 & ~n14406;
  assign n14410 = ~n13226 & ~P1_REG2_REG_22__SCAN_IN;
  assign n14416 = ~n15936 & ~n15497;
  assign n14415 = n15654 & n14919;
  assign n14417 = ~n14416 & ~n14415;
  assign P1_U3271 = ~n14422 | ~n14421;
  assign n14424 = ~n8933 & ~n14423;
  assign n16906 = ~n14425 & ~n14424;
  assign n16926 = ~n16906;
  assign n14427 = ~n14426 | ~P2_B_REG_SCAN_IN;
  assign n14430 = n15240 | n14686;
  assign n14431 = n15240 & P2_REG2_REG_30__SCAN_IN;
  assign P2_U3203 = ~n14433 | ~n14432;
  assign n14446 = n15516 & n14439;
  assign n14442 = ~n15902 & ~n15518;
  assign n14440 = ~n15521 | ~n15883;
  assign n15120 = ~P1_REG3_REG_19__SCAN_IN | ~P1_U3086;
  assign n14441 = ~n14440 | ~n15120;
  assign n14443 = ~n15916 | ~n15439;
  assign P1_U3219 = ~n14448 | ~n14447;
  assign n14469 = ~n14450 & ~n14449;
  assign n14454 = P1_REG2_REG_17__SCAN_IN ^ n14755;
  assign n14452 = ~n14457 | ~P1_REG2_REG_16__SCAN_IN;
  assign n14456 = ~n14454 & ~n14453;
  assign n14455 = ~n15137 | ~n14748;
  assign n14465 = ~n14456 & ~n14455;
  assign n14461 = P1_REG1_REG_17__SCAN_IN ^ n14755;
  assign n14459 = ~n14457 | ~P1_REG1_REG_16__SCAN_IN;
  assign n14463 = ~n14461 & ~n14460;
  assign n14462 = ~n14756 | ~n8934;
  assign n14464 = ~n14463 & ~n14462;
  assign n14470 = ~n15122 | ~P1_ADDR_REG_17__SCAN_IN;
  assign P1_U3260 = ~n14471 | ~n14470;
  assign n14478 = ~n15355 | ~n14492;
  assign n14477 = ~P2_REG3_REG_20__SCAN_IN | ~P2_U3151;
  assign n14484 = ~n14478 | ~n14477;
  assign n14482 = ~n15602 | ~n14507;
  assign n14480 = ~n16702 & ~n15601;
  assign n14479 = ~n16721 & ~n15146;
  assign n14481 = ~n14480 & ~n14479;
  assign P2_U3173 = ~n14486 | ~n14485;
  assign n16888 = ~n14637 & ~n16714;
  assign n14490 = ~n14488 & ~n14487;
  assign n14497 = ~n14494 | ~n14493;
  assign n14648 = ~n14497 | ~n14496;
  assign n14499 = ~n16721 & ~n15559;
  assign n14498 = ~n16696 & ~n16411;
  assign n14500 = ~n14499 & ~n14498;
  assign n14504 = n16419 | P2_REG2_REG_20__SCAN_IN;
  assign n14508 = ~n14507 | ~n16358;
  assign P2_U3213 = ~n14513 | ~n14512;
  assign n14519 = ~n16444 | ~P2_REG1_REG_20__SCAN_IN;
  assign P2_U3479 = ~n14520 | ~n14519;
  assign n14522 = ~n16439 | ~P2_REG0_REG_20__SCAN_IN;
  assign P2_U3447 = ~n14523 | ~n14522;
  assign n14532 = ~n16378 | ~P1_REG0_REG_22__SCAN_IN;
  assign P1_U3512 = ~n14533 | ~n14532;
  assign n14535 = ~n16383 | ~P1_REG1_REG_22__SCAN_IN;
  assign P1_U3544 = ~n14536 | ~n14535;
  assign n14538 = ~n16444 | ~P2_REG1_REG_30__SCAN_IN;
  assign P2_U3489 = ~n14539 | ~n14538;
  assign n14541 = ~n16439 | ~P2_REG0_REG_30__SCAN_IN;
  assign P2_U3457 = ~n14542 | ~n14541;
  assign n14818 = ~n14546 & ~n14545;
  assign n14549 = ~n14548 & ~n16198;
  assign n14822 = ~n14549 & ~n16113;
  assign n14551 = ~n15933 | ~n15484;
  assign n14553 = ~n13226 & ~P1_REG2_REG_23__SCAN_IN;
  assign n14563 = ~n14671 | ~n15659;
  assign n14559 = ~n15083 | ~n15964;
  assign n14558 = ~n15654 | ~n15091;
  assign n14560 = ~n14559 | ~n14558;
  assign P1_U3270 = ~n14567 | ~n14566;
  assign n14569 = ~n8933 & ~n14568;
  assign n16912 = ~n14570 & ~n14569;
  assign n14571 = n15240 & P2_REG2_REG_31__SCAN_IN;
  assign P2_U3202 = ~n14574 | ~n14573;
  assign n14709 = ~n14578 | ~n14577;
  assign n14581 = ~n15398 | ~P2_ADDR_REG_15__SCAN_IN;
  assign n14580 = ~n14698 | ~n15396;
  assign n14582 = ~n14581 | ~n14580;
  assign n14595 = ~n14583 & ~n14582;
  assign n14588 = ~n14586;
  assign n14589 = ~n14588 | ~n14587;
  assign n14592 = ~n15386 | ~P2_REG2_REG_15__SCAN_IN;
  assign n14591 = ~n15388 | ~P2_REG1_REG_15__SCAN_IN;
  assign n14697 = ~n14592 | ~n14591;
  assign n14593 = n14696 ^ ~n14695;
  assign n14716 = ~n14602 | ~n14601;
  assign P2_U3197 = ~n14605 | ~n14604;
  assign n14619 = n15516 & n14609;
  assign n14615 = ~n14610 & ~n15094;
  assign n14613 = ~n15439 | ~n14611;
  assign n14612 = ~P1_REG3_REG_20__SCAN_IN | ~P1_U3086;
  assign n14614 = ~n14613 | ~n14612;
  assign n14616 = ~n14615 & ~n14614;
  assign P1_U3233 = ~n14621 | ~n14620;
  assign n14633 = n15602 & n14652;
  assign n14629 = ~n16703 & ~n15603;
  assign n14627 = ~n15604 | ~n16734;
  assign n14626 = ~P2_REG3_REG_21__SCAN_IN | ~P2_U3151;
  assign n14628 = ~n14627 | ~n14626;
  assign n14630 = ~n14629 & ~n14628;
  assign P2_U3163 = ~n14635 | ~n14634;
  assign n14639 = ~n14638 & ~n14637;
  assign n14772 = ~n14639 & ~n16714;
  assign n14643 = ~n14641 | ~n16345;
  assign n14642 = ~n16734 | ~n16346;
  assign n14646 = n16419 | P2_REG2_REG_21__SCAN_IN;
  assign n14651 = ~n14648 & ~n16888;
  assign n14653 = ~n14652 | ~n16358;
  assign P2_U3212 = ~n14658 | ~n14657;
  assign n14664 = ~n16444 | ~P2_REG1_REG_21__SCAN_IN;
  assign P2_U3480 = ~n14665 | ~n14664;
  assign n14667 = ~n16439 | ~P2_REG0_REG_21__SCAN_IN;
  assign P2_U3448 = ~n14668 | ~n14667;
  assign n14673 = ~n15952 & ~n15536;
  assign n14672 = ~n15045 & ~n14935;
  assign n14682 = ~n14679 | ~n14678;
  assign n14680 = ~n16383 | ~P1_REG1_REG_23__SCAN_IN;
  assign P1_U3545 = ~n14681 | ~n14680;
  assign n14683 = ~n16378 | ~P1_REG0_REG_23__SCAN_IN;
  assign P1_U3513 = ~n14684 | ~n14683;
  assign n14690 = ~n14687 | ~n14686;
  assign n14688 = ~n16439 | ~P2_REG0_REG_31__SCAN_IN;
  assign P2_U3458 = ~n14689 | ~n14688;
  assign n14691 = ~n16444 | ~P2_REG1_REG_31__SCAN_IN;
  assign P2_U3490 = ~n14692 | ~n14691;
  assign n14694 = ~n15398 | ~P2_ADDR_REG_16__SCAN_IN;
  assign n14693 = ~n15192 | ~n15396;
  assign n14706 = ~n14694 | ~n14693;
  assign n14699 = ~n14697;
  assign n14700 = ~n14699 | ~n14698;
  assign n14703 = ~n15386 | ~P2_REG2_REG_16__SCAN_IN;
  assign n14702 = ~n15388 | ~P2_REG1_REG_16__SCAN_IN;
  assign n15191 = ~n14703 | ~n14702;
  assign n15178 = ~n14712 | ~n14711;
  assign n15207 = ~n14720 | ~n14719;
  assign P2_U3198 = ~n14723 | ~n14722;
  assign n14745 = n15516 & n14735;
  assign n14741 = ~n14737 & ~n15094;
  assign n14739 = ~n15439 | ~n15933;
  assign n14738 = ~P1_REG3_REG_21__SCAN_IN | ~P1_U3086;
  assign n14740 = ~n14739 | ~n14738;
  assign n14742 = ~n14741 & ~n14740;
  assign P1_U3223 = ~n14747 | ~n14746;
  assign n14751 = P1_REG2_REG_18__SCAN_IN ^ ~n14754;
  assign n14749 = ~P1_REG2_REG_17__SCAN_IN | ~n14755;
  assign n14753 = ~n14751 & ~n14750;
  assign n14752 = ~n15137 | ~n15134;
  assign n14759 = P1_REG1_REG_18__SCAN_IN ^ ~n14754;
  assign n14757 = ~P1_REG1_REG_17__SCAN_IN | ~n14755;
  assign n14761 = ~n14759 & ~n14758;
  assign n14764 = ~n15119 | ~n15132;
  assign n14768 = ~n15122 | ~P1_ADDR_REG_18__SCAN_IN;
  assign P1_U3261 = ~n14769 | ~n14768;
  assign n14774 = ~n14772 | ~n14771;
  assign n14776 = ~n14774 | ~n14773;
  assign n16892 = ~n14775 | ~n14854;
  assign n14845 = ~n14776 | ~n16892;
  assign n14777 = n14776 | n16892;
  assign n14798 = ~n14782 & ~n14781;
  assign n14783 = n16419 | P2_REG2_REG_22__SCAN_IN;
  assign n14853 = ~n14787 | ~n14786;
  assign n14788 = ~n16358 | ~n14808;
  assign P2_U3211 = ~n14793 | ~n14792;
  assign n14795 = ~n16730 & ~n16433;
  assign n14799 = ~n16439 | ~P2_REG0_REG_22__SCAN_IN;
  assign P2_U3449 = ~n14800 | ~n14799;
  assign n14802 = ~n16444 | ~P2_REG1_REG_22__SCAN_IN;
  assign P2_U3481 = ~n14803 | ~n14802;
  assign n14807 = ~n15355 | ~n16724;
  assign n14806 = ~P2_REG3_REG_22__SCAN_IN | ~P2_U3151;
  assign n14814 = ~n14807 | ~n14806;
  assign n14812 = ~n16454 & ~n15146;
  assign n14813 = n14812 | n14811;
  assign P2_U3175 = ~n14816 | ~n14815;
  assign n16117 = ~n15965 | ~n15045;
  assign n16202 = ~n16051 | ~n16117;
  assign n14820 = ~n14818 | ~n14817;
  assign n14930 = ~n14824 | ~n14823;
  assign n14898 = ~n15965 & ~n14830;
  assign n14841 = n14877 | n14838;
  assign n14839 = ~n16378 | ~P1_REG0_REG_24__SCAN_IN;
  assign P1_U3514 = ~n14840 | ~n14839;
  assign n14842 = ~n16383 | ~P1_REG1_REG_24__SCAN_IN;
  assign P1_U3546 = ~n14843 | ~n14842;
  assign n14990 = ~n14845 | ~n16740;
  assign n14848 = ~n15334 | ~n16346;
  assign n14847 = ~n16734 | ~n16345;
  assign n14867 = ~n14850 & ~n14849;
  assign n14851 = n16419 | P2_REG2_REG_23__SCAN_IN;
  assign n14856 = ~n14853 & ~n16892;
  assign n14858 = ~n14991 | ~n16424;
  assign n14857 = ~n15218 | ~n16358;
  assign P2_U3210 = ~n14862 | ~n14861;
  assign n14870 = ~n14867 | ~n14866;
  assign n14868 = ~n16444 | ~P2_REG1_REG_23__SCAN_IN;
  assign P2_U3482 = ~n14869 | ~n14868;
  assign n14871 = ~n16439 | ~P2_REG0_REG_23__SCAN_IN;
  assign P2_U3450 = ~n14872 | ~n14871;
  assign n14876 = ~n15502 & ~n15983;
  assign n14875 = ~n14874 & ~n14873;
  assign n14889 = ~n14876 & ~n14875;
  assign n14882 = ~n15166 & ~n15497;
  assign P1_U3269 = ~n14889 | ~n14888;
  assign n14893 = ~n14890 & ~n14967;
  assign n14896 = ~n14970 & ~n14895;
  assign n16011 = ~n14897 & ~n14896;
  assign n15072 = ~n15984 | ~n14898;
  assign n15071 = ~n15429 & ~n15072;
  assign n15656 = n15670 & n14899;
  assign n16038 = ~n16133;
  assign n14901 = ~n14900 | ~P1_B_REG_SCAN_IN;
  assign n15640 = ~n15533 | ~n14901;
  assign n14976 = ~n13226 | ~n15028;
  assign n14902 = ~n15323 | ~P1_REG2_REG_30__SCAN_IN;
  assign n14903 = ~n14976 | ~n14902;
  assign P1_U3264 = ~n14906 | ~n14905;
  assign n14910 = ~n14908 | ~n14907;
  assign n14913 = ~n15439 | ~n15949;
  assign n14912 = ~P1_REG3_REG_22__SCAN_IN | ~P1_U3086;
  assign n14916 = ~n14913 | ~n14912;
  assign n14915 = ~n15094 & ~n14914;
  assign n14917 = ~n14916 & ~n14915;
  assign n14920 = n15516 & n14919;
  assign P1_U3235 = ~n14923 | ~n14922;
  assign n16204 = ~n14924 & ~n16054;
  assign n15055 = ~n14928 & ~n14927;
  assign n14933 = n14931 & n16117;
  assign n15059 = ~n14933 | ~n16204;
  assign n14937 = ~n15045 & ~n15639;
  assign n14936 = ~n15308 & ~n14935;
  assign n14938 = ~n14937 & ~n14936;
  assign n14961 = ~n14941 & ~n14940;
  assign n14942 = n13226 | P1_REG2_REG_25__SCAN_IN;
  assign n14947 = ~n15984 & ~n15497;
  assign n14946 = n15654 & n15042;
  assign P1_U3268 = ~n14953 | ~n14952;
  assign n14956 = ~n15968 | ~n16369;
  assign n14964 = ~n14961 | ~n14960;
  assign n14962 = ~n16383 | ~P1_REG1_REG_25__SCAN_IN;
  assign P1_U3547 = ~n14963 | ~n14962;
  assign n14965 = ~n16378 | ~P1_REG0_REG_25__SCAN_IN;
  assign P1_U3515 = ~n14966 | ~n14965;
  assign n14972 = ~n14968 & ~n14967;
  assign n14969 = ~P2_DATAO_REG_31__SCAN_IN;
  assign n16037 = ~n14972 & ~n14971;
  assign n14975 = ~n15323 | ~P1_REG2_REG_31__SCAN_IN;
  assign n14977 = ~n14976 | ~n14975;
  assign P1_U3263 = ~n14980 | ~n14979;
  assign n14987 = ~n14984 | ~n14983;
  assign n14985 = ~n16383 | ~P1_REG1_REG_30__SCAN_IN;
  assign P1_U3552 = ~n14986 | ~n14985;
  assign n14988 = ~n16378 | ~P1_REG0_REG_30__SCAN_IN;
  assign P1_U3520 = ~n14989 | ~n14988;
  assign n14993 = ~n14990 | ~n16895;
  assign n16753 = ~n15234 | ~n15343;
  assign n16901 = ~n14995 & ~n14994;
  assign n14996 = ~n14997 | ~n16901;
  assign n15002 = n14998 | n15229;
  assign n15000 = ~n15446 & ~n15559;
  assign n14999 = ~n16454 & ~n16411;
  assign n15006 = ~n15003 & ~n16895;
  assign n15247 = ~n15006 & ~n15005;
  assign n15021 = ~n15008 & ~n15007;
  assign n15009 = n16419 | P2_REG2_REG_24__SCAN_IN;
  assign n15012 = ~n15341 | ~n16358;
  assign n15011 = ~n15343 | ~n16424;
  assign P2_U3209 = ~n15016 | ~n15015;
  assign n15024 = ~n15021 | ~n15020;
  assign n15022 = ~n16439 | ~P2_REG0_REG_24__SCAN_IN;
  assign P2_U3451 = ~n15023 | ~n15022;
  assign n15025 = ~n16444 | ~P2_REG1_REG_24__SCAN_IN;
  assign P2_U3483 = ~n15026 | ~n15025;
  assign n15034 = ~n15031 | ~n15030;
  assign n15032 = ~n16378 | ~P1_REG0_REG_31__SCAN_IN;
  assign P1_U3521 = ~n15033 | ~n15032;
  assign n15035 = ~n16383 | ~P1_REG1_REG_31__SCAN_IN;
  assign P1_U3553 = ~n15036 | ~n15035;
  assign n15040 = n15038 | n15037;
  assign n15041 = ~n15040 | ~n15039;
  assign n15049 = ~n15516 | ~n15042;
  assign n15044 = ~n15439 | ~n15520;
  assign n15043 = ~P1_REG3_REG_25__SCAN_IN | ~P1_U3086;
  assign n15047 = ~n15044 | ~n15043;
  assign n15046 = ~n15094 & ~n15045;
  assign n15048 = ~n15047 & ~n15046;
  assign n15050 = ~n15049 | ~n15048;
  assign P1_U3225 = ~n15053 | ~n15052;
  assign n16299 = ~n15429 & ~n15308;
  assign n15056 = ~n15055 | ~n15054;
  assign n15307 = ~n15056 | ~n15982;
  assign n15062 = ~n15059 | ~n15058;
  assign n15314 = ~n15062 | ~n15061;
  assign n15064 = ~n15969 | ~n15484;
  assign n15111 = ~n15067 | ~n15066;
  assign n15076 = ~n15429 | ~n15660;
  assign n15075 = ~n15654 | ~n15430;
  assign n15084 = ~n15999 | ~n15083;
  assign P1_U3267 = ~n15085 | ~n15084;
  assign n15157 = n15087 & n15086;
  assign n15156 = ~n15087 & ~n15086;
  assign n15098 = ~n15516 | ~n15091;
  assign n15093 = ~n15439 | ~n15964;
  assign n15092 = ~P1_REG3_REG_23__SCAN_IN | ~P1_U3086;
  assign n15096 = ~n15093 | ~n15092;
  assign n15095 = ~n15094 & ~n15937;
  assign n15097 = ~n15096 & ~n15095;
  assign n15099 = ~n15098 | ~n15097;
  assign P1_U3216 = ~n15102 | ~n15101;
  assign n15113 = ~n15111 & ~n15110;
  assign n15116 = ~n15113 | ~n15112;
  assign n15114 = ~n16383 | ~P1_REG1_REG_26__SCAN_IN;
  assign P1_U3548 = ~n15115 | ~n15114;
  assign n15117 = ~n16378 | ~P1_REG0_REG_26__SCAN_IN;
  assign P1_U3516 = ~n15118 | ~n15117;
  assign n15121 = ~n15119 | ~n16322;
  assign n15131 = ~n15121 | ~n15120;
  assign n15129 = ~P1_ADDR_REG_19__SCAN_IN | ~n15122;
  assign n15124 = ~P1_REG1_REG_18__SCAN_IN | ~n15132;
  assign n15133 = ~P1_REG2_REG_18__SCAN_IN | ~n15132;
  assign P1_U3262 = ~n15140 | ~n15139;
  assign n15145 = ~n15355 | ~n15334;
  assign n15144 = ~P2_REG3_REG_25__SCAN_IN | ~P2_U3151;
  assign n15152 = ~n15145 | ~n15144;
  assign n15442 = ~n16760;
  assign n15147 = ~n15146 & ~n15575;
  assign P2_U3165 = ~n15154 | ~n15153;
  assign n15173 = ~n15516 | ~n15167;
  assign n15169 = ~n15521 | ~n15949;
  assign n15168 = ~P1_REG3_REG_24__SCAN_IN | ~P1_U3086;
  assign n15171 = ~n15169 | ~n15168;
  assign n15170 = ~n15515 & ~n15983;
  assign n15172 = ~n15171 & ~n15170;
  assign n15174 = ~n15173 | ~n15172;
  assign P1_U3229 = ~n15177 | ~n15176;
  assign n15280 = ~n15181 | ~n15180;
  assign n15186 = ~n15398 | ~P2_ADDR_REG_17__SCAN_IN;
  assign n15185 = ~n15184 | ~n15396;
  assign n15187 = ~n15186 | ~n15185;
  assign n15203 = ~n15188 & ~n15187;
  assign n15193 = ~n15191;
  assign n15194 = ~n15193 | ~n15192;
  assign n15197 = ~n15386 | ~P2_REG2_REG_17__SCAN_IN;
  assign n15196 = ~n15388 | ~P2_REG1_REG_17__SCAN_IN;
  assign n15257 = ~n15197 | ~n15196;
  assign n15200 = n15199 | n15198;
  assign n15210 = ~P2_REG2_REG_16__SCAN_IN | ~n15206;
  assign P2_U3199 = ~n15213 | ~n15212;
  assign n15217 = ~n15355 | ~n16734;
  assign n15216 = ~P2_REG3_REG_23__SCAN_IN | ~P2_U3151;
  assign n15224 = ~n15217 | ~n15216;
  assign n15220 = n15218 & n15602;
  assign P2_U3156 = ~n15226 | ~n15225;
  assign n15231 = ~n15229 & ~n15228;
  assign n15453 = ~n15446 & ~n16760;
  assign n16910 = ~n15453 & ~n15230;
  assign n15232 = n15231 | n15452;
  assign n15444 = ~n15231 | ~n15452;
  assign n15233 = ~n15232 | ~n15444;
  assign n15236 = ~n15234 & ~n16411;
  assign n15243 = ~n15239 | ~n16358;
  assign n15245 = ~n16419 & ~P2_REG2_REG_25__SCAN_IN;
  assign n15250 = n15246 | n15245;
  assign n15248 = ~n15247 | ~n16901;
  assign n15451 = ~n15248 | ~n16753;
  assign P2_U3208 = ~n15250 | ~n15249;
  assign n15261 = ~n15257 & ~n15281;
  assign n15259 = ~n15386 & ~P2_REG1_REG_18__SCAN_IN;
  assign n15258 = ~n15388 & ~P2_REG2_REG_18__SCAN_IN;
  assign n15262 = ~n15259 & ~n15258;
  assign n15263 = ~n15261;
  assign n15264 = ~n15263 | ~n15262;
  assign n15266 = ~n15396 & ~n15381;
  assign n15270 = ~n15381;
  assign n15275 = ~n15398 | ~P2_ADDR_REG_18__SCAN_IN;
  assign n15276 = ~n15275 | ~n15274;
  assign P2_U3200 = ~n15287 | ~n15286;
  assign n15295 = ~n15292 | ~n15291;
  assign n15293 = ~n16439 | ~P2_REG0_REG_25__SCAN_IN;
  assign P2_U3452 = ~n15294 | ~n15293;
  assign n15296 = ~n16444 | ~P2_REG1_REG_25__SCAN_IN;
  assign P2_U3484 = ~n15297 | ~n15296;
  assign n15305 = ~n15669 & ~n15502;
  assign n15303 = ~n15517 | ~n15654;
  assign n15313 = n15305 | n15304;
  assign n16212 = ~n15489 | ~n15488;
  assign n15487 = ~n15311 & ~n15310;
  assign n15316 = ~n15314 | ~n15975;
  assign n15478 = ~n16212 | ~n15316;
  assign n15417 = ~n15321 & ~n15320;
  assign P1_U3266 = ~n15327 | ~n15326;
  assign n15331 = ~n15330 & ~n15329;
  assign n15340 = ~n15355 | ~n15338;
  assign n15339 = ~P2_REG3_REG_24__SCAN_IN | ~P2_U3151;
  assign n15349 = ~n15340 | ~n15339;
  assign n15345 = ~n15341 | ~n15602;
  assign P2_U3169 = ~n15351 | ~n15350;
  assign n15357 = ~n15355 | ~n16759;
  assign n15356 = ~P2_REG3_REG_26__SCAN_IN | ~P2_U3151;
  assign n15359 = ~n15602 | ~n15460;
  assign n15358 = ~n15604 | ~n16779;
  assign n15362 = n15361 | n15360;
  assign P2_U3180 = ~n15365 | ~n15364;
  assign n15379 = ~n15378;
  assign n15387 = ~n15385;
  assign n15391 = ~n15387 | ~n15386;
  assign n15390 = ~n15389 | ~n15388;
  assign n15392 = ~n15391 | ~n15390;
  assign n15397 = ~n15396;
  assign n15402 = ~n15397 & ~n8925;
  assign n15400 = ~n15398 | ~P2_ADDR_REG_19__SCAN_IN;
  assign n15401 = ~n15400 | ~n15399;
  assign n15403 = ~n15402 & ~n15401;
  assign P2_U3201 = ~n15408 | ~n15407;
  assign n15421 = ~n15418 | ~n15417;
  assign n15419 = ~n16383 | ~P1_REG1_REG_27__SCAN_IN;
  assign P1_U3549 = ~n15420 | ~n15419;
  assign n15422 = ~n16378 | ~P1_REG0_REG_27__SCAN_IN;
  assign P1_U3517 = ~n15423 | ~n15422;
  assign n15434 = n15516 & n15430;
  assign n15432 = ~n15521 | ~n15969;
  assign n15431 = ~P1_REG3_REG_26__SCAN_IN | ~P1_U3086;
  assign n15433 = ~n15432 | ~n15431;
  assign n15435 = ~n15434 & ~n15433;
  assign n15440 = ~n15999 | ~n15439;
  assign P1_U3240 = ~n15441 | ~n15440;
  assign n16894 = ~n15552 | ~n15550;
  assign n15551 = ~n15444 | ~n15443;
  assign n15448 = ~n15446 & ~n16411;
  assign n15454 = ~n15452 & ~n15451;
  assign n15471 = ~n15457 & ~n15456;
  assign n15458 = n16419 | P2_REG2_REG_26__SCAN_IN;
  assign n15462 = ~n15576 | ~n16424;
  assign n15461 = ~n16358 | ~n15460;
  assign P2_U3207 = ~n15466 | ~n15465;
  assign n15474 = ~n15471 | ~n15470;
  assign n15472 = ~n16439 | ~P2_REG0_REG_26__SCAN_IN;
  assign P2_U3453 = ~n15473 | ~n15472;
  assign n15475 = ~n16444 | ~P2_REG1_REG_26__SCAN_IN;
  assign P2_U3485 = ~n15476 | ~n15475;
  assign n16128 = ~n15669 & ~n15674;
  assign n15481 = ~n15478 | ~n16227;
  assign n15635 = ~n15482 | ~n15481;
  assign n15490 = ~n15488 | ~n15487;
  assign n15645 = ~n15490 | ~n15489;
  assign n15544 = ~n15492 & ~n15491;
  assign n15493 = n13226 | P1_REG2_REG_28__SCAN_IN;
  assign n15503 = ~n16130 & ~n15502;
  assign n15505 = n15504 | n15503;
  assign P1_U3265 = ~n15508 | ~n15507;
  assign n15512 = ~n15510 | ~n15509;
  assign n15531 = n15514 | n15513;
  assign n15529 = ~n15669 & ~n15515;
  assign n15523 = ~n15521 | ~n15520;
  assign n15522 = ~P1_REG3_REG_27__SCAN_IN | ~P1_U3086;
  assign P1_U3214 = ~n15531 | ~n15530;
  assign n15543 = ~n15542 & ~n15541;
  assign n15547 = ~n15544 | ~n15543;
  assign n15545 = ~n16378 | ~P1_REG0_REG_28__SCAN_IN;
  assign P1_U3518 = ~n15546 | ~n15545;
  assign n15548 = ~n16383 | ~P1_REG1_REG_28__SCAN_IN;
  assign P1_U3550 = ~n15549 | ~n15548;
  assign n15553 = ~n15551 | ~n15550;
  assign n15555 = ~n15553 | ~n15552;
  assign n16340 = ~n15555 | ~n15578;
  assign n15624 = ~n15563 | ~n15562;
  assign n15566 = ~n16358 | ~n15565;
  assign n15567 = ~n16419 | ~n15566;
  assign n15569 = n15568 | n15567;
  assign n15570 = ~n16419 & ~P2_REG2_REG_27__SCAN_IN;
  assign n15581 = n15571 | n15570;
  assign n16782 = ~n15573 | ~n15572;
  assign n16353 = ~n15577 | ~n16783;
  assign P2_U3206 = ~n15581 | ~n15580;
  assign n15620 = ~n15583 & ~n15582;
  assign n15587 = ~n8933 & ~n15586;
  assign n16808 = ~n15588 & ~n15587;
  assign n16397 = ~n16407 & ~n15589;
  assign n15592 = ~n15595 | ~n16775;
  assign n15597 = ~n15596 | ~n16775;
  assign n15610 = ~n15602 | ~n16357;
  assign n15608 = ~n15603 & ~n16775;
  assign n15606 = ~n15604 | ~n16801;
  assign n15605 = ~P2_REG3_REG_28__SCAN_IN | ~P2_U3151;
  assign n15607 = ~n15606 | ~n15605;
  assign n15609 = ~n15608 & ~n15607;
  assign P2_U3160 = ~n15622 | ~n15621;
  assign n15631 = ~n15628 | ~n15627;
  assign n15629 = ~n16439 | ~P2_REG0_REG_27__SCAN_IN;
  assign P2_U3454 = ~n15630 | ~n15629;
  assign n15632 = ~n16444 | ~P2_REG1_REG_27__SCAN_IN;
  assign P2_U3486 = ~n15633 | ~n15632;
  assign n15636 = ~n15635 | ~n15634;
  assign n16370 = ~n16011;
  assign n15638 = n15636 ^ n16215;
  assign n15644 = ~n15638 | ~n15637;
  assign n15642 = ~n15669 & ~n15639;
  assign n15641 = ~n16313 & ~n15640;
  assign n15650 = ~n15644 | ~n15643;
  assign n15647 = ~n16214 | ~n15645;
  assign n16366 = n15648 ^ ~n16215;
  assign n15652 = ~n16376 | ~n13226;
  assign n15651 = n13226 | P1_REG2_REG_29__SCAN_IN;
  assign n15668 = ~n15652 | ~n15651;
  assign n15666 = ~n16366 & ~n15653;
  assign n15664 = n15655 & n15654;
  assign n15665 = n15664 | n15663;
  assign P1_U3356 = ~n15668 | ~n15667;
  assign n15672 = ~n15669 | ~n16045;
  assign n15671 = ~n15670 | ~n15816;
  assign n15676 = ~n15673 & ~n16045;
  assign n15675 = ~n15674 & ~n15816;
  assign n15677 = ~n16299 & ~n16045;
  assign n15678 = ~n16301 | ~n16045;
  assign n16001 = ~n15997 | ~n16045;
  assign n15682 = ~n15680 & ~n16045;
  assign n15681 = ~n16242 & ~n15816;
  assign n15689 = ~n15682 & ~n15681;
  assign n15686 = ~n15683 | ~n16045;
  assign n15685 = ~n15684 | ~n15816;
  assign n15702 = ~n15686 | ~n15685;
  assign n15688 = ~n15702 & ~n15687;
  assign n15706 = ~n15689 & ~n15688;
  assign n15692 = ~n15702 | ~n15690;
  assign n15693 = ~n15692 | ~n15691;
  assign n15699 = ~n15706 | ~n15693;
  assign n15695 = ~n15715 & ~n15816;
  assign n15694 = ~n15714 & ~n16045;
  assign n15717 = ~n15695 & ~n15694;
  assign n15697 = ~n15717 & ~n15696;
  assign n15698 = ~n15697 & ~n16242;
  assign n15700 = ~n15699 | ~n15698;
  assign n15713 = ~n15700 | ~n16021;
  assign n15704 = ~n15702 | ~n15701;
  assign n15705 = ~n15704 | ~n15703;
  assign n15710 = ~n15706 | ~n15705;
  assign n15708 = ~n15707 | ~n15714;
  assign n15709 = n15708 & n16245;
  assign n15711 = ~n15710 | ~n15709;
  assign n15712 = ~n15711 | ~n16045;
  assign n15719 = ~n15713 | ~n15712;
  assign n15716 = ~n15715 | ~n15714;
  assign n15718 = ~n15717 | ~n15716;
  assign n15729 = ~n15719 | ~n15718;
  assign n15721 = ~n15722 & ~n15816;
  assign n15720 = ~n15723 & ~n16045;
  assign n15728 = ~n15721 & ~n15720;
  assign n15727 = ~n15729 & ~n15728;
  assign n15725 = ~n15722 & ~n16045;
  assign n15724 = ~n15723 & ~n15816;
  assign n15726 = ~n15725 & ~n15724;
  assign n15737 = ~n15727 & ~n15726;
  assign n15735 = ~n15729 | ~n15728;
  assign n15733 = ~n15730 | ~n16045;
  assign n15732 = ~n15731 | ~n16021;
  assign n15734 = ~n15733 | ~n15732;
  assign n15736 = ~n15735 | ~n15734;
  assign n15745 = ~n15737 & ~n15736;
  assign n15741 = ~n15738 & ~n16045;
  assign n15740 = ~n15739 & ~n15816;
  assign n15743 = ~n15741 & ~n15740;
  assign n15744 = ~n15743 & ~n15742;
  assign n15749 = ~n15745 & ~n15744;
  assign n15747 = ~n16166 & ~n16045;
  assign n15746 = ~n16259 & ~n15816;
  assign n15748 = ~n15747 & ~n15746;
  assign n15768 = ~n15749 & ~n15748;
  assign n15753 = ~n15750 & ~n16021;
  assign n15752 = ~n15751 & ~n16045;
  assign n15769 = ~n15753 & ~n15752;
  assign n15757 = ~n15768 & ~n15769;
  assign n15766 = ~n16259;
  assign n15755 = ~n15757 | ~n15766;
  assign n15756 = ~n15755 | ~n15754;
  assign n15765 = ~n15756 | ~n16021;
  assign n15758 = ~n15757;
  assign n15763 = ~n15758 | ~n15759;
  assign n15760 = ~n15769 & ~n15759;
  assign n15761 = ~n15760 & ~n16256;
  assign n15762 = ~n15761 & ~n15816;
  assign n15764 = ~n15763 | ~n15762;
  assign n15783 = ~n15765 | ~n15764;
  assign n15767 = ~n15766 & ~n16045;
  assign n15771 = ~n15768 & ~n15767;
  assign n15770 = ~n15769;
  assign n15775 = ~n15772 & ~n16045;
  assign n15774 = ~n15773 & ~n15816;
  assign n15785 = ~n15775 & ~n15774;
  assign n15779 = ~n15776 | ~n16045;
  assign n15778 = ~n15777 | ~n16021;
  assign n15784 = ~n15779 | ~n15778;
  assign n15780 = ~n15785 & ~n15784;
  assign n15787 = ~n15783 | ~n15782;
  assign n15786 = ~n15785 | ~n15784;
  assign n15794 = ~n15787 | ~n15786;
  assign n15791 = ~n15788 & ~n15816;
  assign n15790 = ~n15789 & ~n16045;
  assign n15795 = ~n15791 & ~n15790;
  assign n15793 = ~n15795 | ~n15792;
  assign n15799 = ~n15794 | ~n15793;
  assign n15797 = ~n15795;
  assign n15798 = ~n15797 | ~n15796;
  assign n15809 = ~n15799 | ~n15798;
  assign n15801 = ~n15802 | ~n16045;
  assign n15800 = ~n15803 | ~n16021;
  assign n15808 = ~n15801 | ~n15800;
  assign n15807 = ~n15809 & ~n15808;
  assign n15805 = ~n15802 & ~n16045;
  assign n15804 = ~n15803 & ~n15816;
  assign n15806 = ~n15805 & ~n15804;
  assign n15815 = ~n15807 & ~n15806;
  assign n15813 = ~n15809 | ~n15808;
  assign n15811 = ~n16088 | ~n16045;
  assign n15810 = ~n16270 | ~n16021;
  assign n15812 = ~n15811 | ~n15810;
  assign n15814 = ~n15813 | ~n15812;
  assign n15825 = ~n15815 & ~n15814;
  assign n15818 = ~n15819 & ~n15816;
  assign n15817 = ~n15820 & ~n16045;
  assign n15824 = ~n15825 & ~n15830;
  assign n15822 = ~n15819 & ~n16045;
  assign n15821 = ~n15820 & ~n16021;
  assign n15823 = ~n15822 & ~n15821;
  assign n15848 = ~n15824 & ~n15823;
  assign n15846 = ~n15825 | ~n15830;
  assign n15827 = ~n15830 & ~n15826;
  assign n15828 = ~n15827 & ~n16088;
  assign n15834 = ~n15828 & ~n16045;
  assign n15831 = ~n15830 & ~n15829;
  assign n15832 = ~n15831 & ~n16270;
  assign n15844 = ~n15834 & ~n15833;
  assign n15838 = ~n15835 & ~n16045;
  assign n15837 = ~n15836 & ~n16021;
  assign n15842 = ~n15839 | ~n16045;
  assign n15841 = ~n15840 | ~n16021;
  assign n15854 = ~n15842 | ~n15841;
  assign n15843 = ~n15855 & ~n15854;
  assign n15845 = ~n15844 & ~n15843;
  assign n15847 = ~n15846 | ~n15845;
  assign n15859 = ~n15848 & ~n15847;
  assign n15852 = ~n15849 & ~n16045;
  assign n15851 = ~n15850 & ~n16021;
  assign n15862 = ~n15852 & ~n15851;
  assign n15857 = ~n15862 | ~n15853;
  assign n15856 = ~n15855 | ~n15854;
  assign n15858 = ~n15857 | ~n15856;
  assign n15868 = ~n15859 & ~n15858;
  assign n15861 = ~n16282 | ~n16021;
  assign n15860 = ~n16060 | ~n16045;
  assign n15866 = ~n15861 | ~n15860;
  assign n15864 = ~n15862;
  assign n15865 = ~n15864 | ~n15863;
  assign n15870 = ~n15868 & ~n15867;
  assign n15869 = ~n16282 & ~n16021;
  assign n15871 = ~n15870 & ~n15869;
  assign n15877 = ~n15871 & ~n16056;
  assign n15872 = ~n16060 | ~n16021;
  assign n15875 = ~n16056 & ~n15872;
  assign n15874 = ~n15873 & ~n16021;
  assign n15876 = ~n15875 & ~n15874;
  assign n15879 = ~n15877 & ~n15876;
  assign n15878 = ~n16156 & ~n16045;
  assign n15894 = ~n15879 & ~n15878;
  assign n15881 = ~n15880 & ~n16045;
  assign n15884 = ~n15883 | ~n16021;
  assign n15892 = ~n15895 | ~n15884;
  assign n15886 = ~n15885 | ~n16021;
  assign n15890 = ~n15887 | ~n15886;
  assign n15889 = ~n15888 | ~n16021;
  assign n15891 = ~n15890 | ~n15889;
  assign n15906 = ~n15894 & ~n15893;
  assign n15897 = ~n16229 & ~n16021;
  assign n15899 = ~n16099 | ~n16021;
  assign n15903 = n15902 ^ n15901;
  assign n15914 = ~n15906 & ~n15905;
  assign n15907 = ~n16101 | ~n16021;
  assign n15909 = ~n15908 | ~n16045;
  assign n15911 = ~n15910 & ~n15909;
  assign n15922 = ~n15914 & ~n15913;
  assign n15918 = ~n15915 & ~n16045;
  assign n15917 = ~n15916 & ~n16021;
  assign n15920 = ~n15918 & ~n15917;
  assign n15926 = ~n15922 & ~n15921;
  assign n15924 = ~n15927 & ~n16045;
  assign n15931 = ~n15926 & ~n15925;
  assign n15929 = ~n15927 & ~n16021;
  assign n15928 = ~n16106 & ~n16045;
  assign n15941 = ~n15931 & ~n15930;
  assign n15934 = ~n15933 & ~n16045;
  assign n15939 = ~n15936 | ~n15816;
  assign n15938 = ~n15937 | ~n16045;
  assign n15947 = ~n15941 | ~n15940;
  assign n15945 = ~n15942;
  assign n15957 = ~n15947 | ~n15946;
  assign n15950 = ~n15949 & ~n16045;
  assign n15955 = ~n15952 | ~n15816;
  assign n15954 = ~n15953 | ~n16045;
  assign n15963 = ~n15957 & ~n15956;
  assign n15961 = ~n15958;
  assign n15960 = ~n15959;
  assign n15967 = ~n15963 & ~n15962;
  assign n15966 = n15965 ^ ~n15964;
  assign n15974 = ~n15967 | ~n15966;
  assign n15971 = ~n15968 & ~n16045;
  assign n15970 = ~n15969 & ~n16021;
  assign n15979 = n15974 | n15973;
  assign n15977 = ~n15975 | ~n16045;
  assign n15976 = ~n16301 | ~n15816;
  assign n15992 = ~n15979 | ~n15978;
  assign n15981 = ~n16051 | ~n16045;
  assign n15980 = ~n16117 | ~n15816;
  assign n15990 = n15985 | n15982;
  assign n15993 = ~n15992 & ~n15991;
  assign n15995 = ~n15994 & ~n15993;
  assign n16004 = ~n15996 | ~n15995;
  assign n16000 = ~n15999 | ~n16045;
  assign n16003 = ~n16002 | ~n16001;
  assign n16005 = ~n16004 | ~n16003;
  assign n16016 = ~n16006 & ~n16005;
  assign n16010 = ~n16130 | ~n16045;
  assign n16009 = ~n16011 | ~n15816;
  assign n16012 = ~n16130 | ~n16011;
  assign n16030 = ~n16016 & ~n16015;
  assign n16024 = ~n16134 & ~n16021;
  assign n16022 = ~n16313;
  assign n16138 = ~n16022 | ~n16133;
  assign n16023 = ~n16138 & ~n16045;
  assign n16031 = ~n16024 & ~n16023;
  assign n16035 = ~n16314 | ~n15816;
  assign n16025 = ~n16138;
  assign n16032 = ~n16025 | ~n16045;
  assign n16042 = ~n16030 & ~n16029;
  assign n16317 = ~n16037 | ~n16133;
  assign n16208 = ~n16039 | ~n16038;
  assign n16043 = ~n16317 & ~n16045;
  assign n16148 = ~n16320 | ~n16045;
  assign n16046 = ~n16152 | ~n16148;
  assign n16145 = ~n16046 | ~n16322;
  assign n16052 = ~n16117 | ~n16050;
  assign n16053 = ~n16052 | ~n16051;
  assign n16057 = ~n16228 & ~n16056;
  assign n16096 = ~n16156 | ~n16282;
  assign n16281 = ~n16060 | ~n16059;
  assign n16279 = ~n16062 | ~n16061;
  assign n16066 = ~n16064 & ~n16063;
  assign n16068 = ~n16066 & ~n16065;
  assign n16069 = ~n16068 & ~n16067;
  assign n16070 = ~n16069 & ~n16252;
  assign n16071 = ~n16070 & ~n16254;
  assign n16072 = ~n16071 & ~n16166;
  assign n16074 = ~n16072 & ~n16259;
  assign n16080 = ~n16074 & ~n16073;
  assign n16084 = ~n16076 & ~n16075;
  assign n16079 = ~n16078 & ~n16077;
  assign n16264 = ~n16084 | ~n16079;
  assign n16082 = ~n16080 & ~n16264;
  assign n16081 = ~n16270;
  assign n16087 = ~n16082 & ~n16081;
  assign n16086 = ~n16084 | ~n16083;
  assign n16265 = n16086 & n16085;
  assign n16090 = ~n16087 | ~n16265;
  assign n16268 = ~n16088;
  assign n16089 = ~n16274 & ~n16268;
  assign n16091 = ~n16090 | ~n16089;
  assign n16092 = ~n16091 | ~n16271;
  assign n16093 = ~n16092 & ~n16276;
  assign n16094 = ~n16279 & ~n16093;
  assign n16095 = ~n16281 & ~n16094;
  assign n16097 = ~n16096 & ~n16095;
  assign n16098 = ~n16286 & ~n16097;
  assign n16100 = ~n16291 & ~n16098;
  assign n16102 = ~n16100 | ~n16099;
  assign n16103 = ~n16102 | ~n16101;
  assign n16104 = ~n16294 | ~n16103;
  assign n16105 = n16296 | n16104;
  assign n16123 = ~n16105 | ~n16301;
  assign n16108 = ~n16106;
  assign n16114 = ~n16112 & ~n16111;
  assign n16118 = ~n16116 & ~n16115;
  assign n16119 = ~n16118 | ~n16117;
  assign n16127 = ~n16130 & ~n16370;
  assign n16147 = ~n16145 | ~n16144;
  assign n16223 = ~n16147 | ~n16146;
  assign n16151 = ~n16150 & ~n16149;
  assign n16153 = ~n16152 | ~n16151;
  assign n16157 = ~n16155;
  assign n16163 = ~n16159 | ~n16158;
  assign n16162 = ~n16161 | ~n16160;
  assign n16165 = ~n16163 & ~n16162;
  assign n16167 = ~n16165 | ~n16164;
  assign n16169 = ~n16167 & ~n16166;
  assign n16171 = ~n16169 | ~n16168;
  assign n16172 = ~n16171 & ~n16170;
  assign n16174 = ~n16173 | ~n16172;
  assign n16176 = ~n16175 & ~n16174;
  assign n16178 = ~n16177 | ~n16176;
  assign n16180 = ~n16179 & ~n16178;
  assign n16182 = ~n16181 | ~n16180;
  assign n16184 = ~n16183 & ~n16182;
  assign n16186 = ~n16185 | ~n16184;
  assign n16188 = ~n16187 & ~n16186;
  assign n16191 = ~n16232 & ~n16190;
  assign n16193 = ~n16192 | ~n16191;
  assign n16195 = ~n16194 & ~n16193;
  assign n16197 = ~n16196 | ~n16195;
  assign n16199 = ~n16198 & ~n16197;
  assign n16203 = ~n16202 & ~n16201;
  assign n16216 = ~n16214 & ~n16213;
  assign n16217 = ~n16216 | ~n16215;
  assign n16225 = ~n16223 | ~n16222;
  assign n16327 = ~n16225 | ~n16224;
  assign n16305 = ~n16227;
  assign n16231 = ~n16229 & ~n16228;
  assign n16234 = ~n16231 & ~n16230;
  assign n16233 = ~n16232;
  assign n16288 = ~n16234 & ~n16233;
  assign n16241 = ~n16235;
  assign n16239 = ~n16237 | ~n16236;
  assign n16240 = ~n16239 & ~n16238;
  assign n16243 = ~n16241 & ~n16240;
  assign n16247 = ~n16243 & ~n16242;
  assign n16246 = ~n16245 | ~n16244;
  assign n16251 = ~n16247 & ~n16246;
  assign n16250 = ~n16249 | ~n16248;
  assign n16253 = ~n16251 & ~n16250;
  assign n16255 = ~n16253 & ~n16252;
  assign n16258 = ~n16255 & ~n16254;
  assign n16257 = ~n16260 | ~n16256;
  assign n16262 = n16258 | n16257;
  assign n16261 = ~n16260 | ~n16259;
  assign n16263 = ~n16262 | ~n16261;
  assign n16267 = ~n16264 & ~n16263;
  assign n16266 = ~n16265;
  assign n16269 = ~n16267 & ~n16266;
  assign n16273 = ~n16269 & ~n16268;
  assign n16272 = ~n16271 | ~n16270;
  assign n16275 = ~n16273 & ~n16272;
  assign n16277 = ~n16275 & ~n16274;
  assign n16278 = ~n16277 & ~n16276;
  assign n16280 = ~n16279 & ~n16278;
  assign n16284 = ~n16281 & ~n16280;
  assign n16283 = ~n16282;
  assign n16285 = ~n16284 & ~n16283;
  assign n16287 = ~n16286 & ~n16285;
  assign n16290 = ~n16288 & ~n16287;
  assign n16292 = ~n16290 & ~n16289;
  assign n16293 = ~n16292 & ~n16291;
  assign n16295 = ~n16294 | ~n16293;
  assign n16298 = ~n16296 & ~n16295;
  assign n16302 = ~n16301;
  assign n16329 = ~n16327 | ~n16326;
  assign n16338 = ~n16329 | ~n16333;
  assign n16336 = ~n16331 & ~n16330;
  assign n16334 = ~n16333 | ~n16332;
  assign n16335 = ~n16334 | ~P1_B_REG_SCAN_IN;
  assign n16337 = n16336 | n16335;
  assign P1_U3242 = ~n16338 | ~n16337;
  assign n16341 = ~n16340 | ~n16339;
  assign n16399 = ~n16341 | ~n16900;
  assign n16344 = ~n16343 & ~n16342;
  assign n16350 = ~n16344 & ~n11752;
  assign n16391 = ~n16350 & ~n16349;
  assign n16351 = n16419 | P2_REG2_REG_28__SCAN_IN;
  assign n16355 = ~n16353 | ~n16898;
  assign n16406 = ~n16355 | ~n16354;
  assign P2_U3205 = ~n16364 | ~n16363;
  assign n16374 = ~n16366 & ~n16365;
  assign n16375 = ~n16374 & ~n16373;
  assign n16380 = ~n16382 | ~n16377;
  assign n16379 = ~n16378 | ~P1_REG0_REG_29__SCAN_IN;
  assign P1_U3519 = ~n16380 | ~n16379;
  assign n16385 = ~n16382 | ~n16381;
  assign n16384 = ~n16383 | ~P1_REG1_REG_29__SCAN_IN;
  assign P1_U3551 = ~n16385 | ~n16384;
  assign n16394 = ~n16391 | ~n16390;
  assign n16392 = ~n16439 | ~P2_REG0_REG_28__SCAN_IN;
  assign P2_U3455 = ~n16393 | ~n16392;
  assign n16395 = ~n16444 | ~P2_REG1_REG_28__SCAN_IN;
  assign P2_U3487 = ~n16396 | ~n16395;
  assign n16402 = ~n16401 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n16802 = ~n16403 | ~n16402;
  assign n16903 = ~n16927 | ~n16923;
  assign n16418 = ~n16405 & ~n11752;
  assign n16422 = n16924 ^ n16903;
  assign n16414 = ~n16809 & ~n16411;
  assign n16413 = ~n16913 & ~n16412;
  assign n16417 = ~n16416 | ~n16415;
  assign n16420 = n16419 | P2_REG2_REG_29__SCAN_IN;
  assign P2_U3204 = ~n16430 | ~n16429;
  assign n16435 = ~n16432 & ~n16431;
  assign n16436 = ~n16435 & ~n16434;
  assign n16443 = ~n16437 | ~n16436;
  assign n16440 = ~n16439 | ~P2_REG0_REG_29__SCAN_IN;
  assign P2_U3456 = ~n16441 | ~n16440;
  assign n16445 = ~n16444 | ~P2_REG1_REG_29__SCAN_IN;
  assign P2_U3488 = ~n16446 | ~n16445;
  assign n16448 = ~n16759 & ~n16798;
  assign n16447 = ~n16760 & ~n16591;
  assign n16450 = ~n16753 | ~n16798;
  assign n16449 = ~n16754 | ~n16591;
  assign n16452 = ~n16454 | ~n16798;
  assign n16451 = ~n16453 | ~n16774;
  assign n16455 = ~n16454 & ~n16453;
  assign n16464 = ~n16461 | ~n16798;
  assign n16463 = ~n16462 | ~n16774;
  assign n16469 = ~n16615 | ~n16774;
  assign n16468 = ~n16604 | ~n16798;
  assign n16483 = ~n16471 & ~n16470;
  assign n16474 = ~n16483 & ~n16939;
  assign n16473 = ~n16472 | ~n16798;
  assign n16481 = ~n16474 & ~n16473;
  assign n16478 = ~n16475 | ~n16798;
  assign n16477 = ~n16476 | ~n16591;
  assign n16488 = ~n16478 | ~n16477;
  assign n16480 = ~n16488 | ~n16479;
  assign n16484 = ~n16483 & ~n16798;
  assign n16491 = ~n16505;
  assign n16490 = ~n16488;
  assign n16493 = ~n16495 | ~n16591;
  assign n16492 = ~n16496 | ~n16798;
  assign n16500 = ~n16494 | ~n16501;
  assign n16498 = ~n16495 | ~n16798;
  assign n16497 = ~n16496 | ~n16774;
  assign n16499 = ~n16498 | ~n16497;
  assign n16591 = n16774;
  assign n16509 = ~n16506 & ~n16591;
  assign n16508 = ~n16507 & ~n16798;
  assign n16515 = ~n16509 & ~n16508;
  assign n16511 = ~n16515 & ~n16510;
  assign n16530 = ~n16514 | ~n16513;
  assign n16519 = ~n16515;
  assign n16518 = ~n16517 & ~n16516;
  assign n16528 = ~n16519 & ~n16518;
  assign n16521 = ~n16522 | ~n16591;
  assign n16520 = ~n16523 | ~n16798;
  assign n16534 = ~n16521 | ~n16520;
  assign n16526 = ~n16534;
  assign n16525 = ~n16522 | ~n16798;
  assign n16524 = ~n16523 | ~n16774;
  assign n16527 = ~n16526 & ~n16533;
  assign n16529 = ~n16528 & ~n16527;
  assign n16532 = ~n16540 & ~n16798;
  assign n16531 = ~n16542 & ~n16774;
  assign n16537 = ~n16532 & ~n16531;
  assign n16535 = ~n16533;
  assign n16536 = ~n16535 & ~n16534;
  assign n16538 = ~n16537 & ~n16536;
  assign n16547 = ~n16539 | ~n16538;
  assign n16541 = ~n16540 & ~n16591;
  assign n16545 = ~n16553 | ~n16541;
  assign n16543 = ~n16542 & ~n16798;
  assign n16544 = ~n16548 | ~n16543;
  assign n16546 = ~n16545 | ~n16544;
  assign n16559 = ~n16547 | ~n16546;
  assign n16549 = ~n16548;
  assign n16552 = ~n16549 & ~n16774;
  assign n16563 = ~n16551 | ~n16550;
  assign n16557 = ~n16552 | ~n16563;
  assign n16555 = ~n16554 & ~n16798;
  assign n16569 = ~n16559 | ~n16558;
  assign n16561 = ~n16560;
  assign n16562 = ~n16561 & ~n16591;
  assign n16567 = ~n16570 | ~n16562;
  assign n16565 = ~n16564 & ~n16798;
  assign n16566 = ~n16574 | ~n16565;
  assign n16581 = ~n16569 | ~n16568;
  assign n16572 = ~n16571 & ~n16798;
  assign n16579 = ~n16573 | ~n16572;
  assign n16577 = ~n16575 & ~n16591;
  assign n16578 = ~n16577 | ~n16576;
  assign n16580 = ~n16579 | ~n16578;
  assign n16590 = ~n16581 | ~n16580;
  assign n16583 = ~n16582 & ~n16798;
  assign n16588 = ~n16592 | ~n16583;
  assign n16585 = ~n16584 & ~n16774;
  assign n16596 = ~n16590 | ~n16589;
  assign n16593 = ~n16592 & ~n16591;
  assign n16595 = ~n16594 & ~n16593;
  assign n16599 = ~n16596 | ~n16595;
  assign n16598 = ~n16597 & ~n16798;
  assign n16600 = ~n16599 & ~n16598;
  assign n16601 = ~n16617 | ~n16600;
  assign n16602 = ~n16620 & ~n16601;
  assign n16606 = ~n16605 & ~n16798;
  assign n16612 = ~n16607 & ~n16606;
  assign n16609 = ~n16608 & ~n16774;
  assign n16611 = ~n16610 & ~n16609;
  assign n16613 = ~n16612 & ~n16611;
  assign n16618 = ~n16616 | ~n16615;
  assign n16635 = ~n16627 | ~n16626;
  assign n16629 = ~n16628 | ~n16798;
  assign n16632 = ~n16631 | ~n16798;
  assign n16641 = ~n16635 | ~n16634;
  assign n16639 = ~n16636 | ~n16774;
  assign n16643 = ~n16637 | ~n16645;
  assign n16638 = ~n16643 | ~n16798;
  assign n16649 = ~n16641 | ~n16640;
  assign n16644 = ~n16642 | ~n16798;
  assign n16646 = ~n16645 | ~n16798;
  assign n16655 = ~n16649 | ~n16648;
  assign n16653 = ~n16650 | ~n16774;
  assign n16652 = ~n16651 | ~n16798;
  assign n16684 = ~n16655 | ~n16654;
  assign n16656 = ~n16669 | ~n16774;
  assign n16683 = ~n16657 | ~n16656;
  assign n16670 = ~n16684 | ~n16683;
  assign n16664 = ~n16670 | ~n16658;
  assign n16663 = n16662 & n16774;
  assign n16674 = ~n16664 | ~n16663;
  assign n16667 = ~n16683 | ~n16665;
  assign n16672 = n16668 & n16798;
  assign n16671 = ~n16670 | ~n16669;
  assign n16673 = ~n16672 | ~n16671;
  assign n16688 = ~n16674 | ~n16673;
  assign n16678 = ~n16675 | ~n16798;
  assign n16677 = ~n16676 | ~n16774;
  assign n16690 = ~n16678 | ~n16677;
  assign n16682 = ~n16679 & ~n16798;
  assign n16681 = ~n16680 & ~n16774;
  assign n16685 = ~n16684 & ~n16683;
  assign n16692 = ~n16688 | ~n16687;
  assign n16691 = ~n16690 | ~n16689;
  assign n16701 = ~n16692 | ~n16691;
  assign n16694 = ~n16695 | ~n16798;
  assign n16693 = ~n16696 | ~n16774;
  assign n16698 = ~n16695 | ~n16774;
  assign n16697 = ~n16696 | ~n16798;
  assign n16713 = n16701 & n16700;
  assign n16705 = ~n16702 | ~n16798;
  assign n16704 = ~n16703 | ~n16774;
  assign n16710 = ~n16709 | ~n16708;
  assign n16717 = ~n16713 & ~n16712;
  assign n16716 = ~n16715 & ~n16714;
  assign n16719 = ~n16717 & ~n16716;
  assign n16729 = ~n16719 & ~n16718;
  assign n16722 = ~n16720 & ~n16798;
  assign n16725 = ~n16723 & ~n16774;
  assign n16739 = ~n16729 & ~n16728;
  assign n16733 = ~n16730 | ~n16798;
  assign n16732 = ~n16731 | ~n16774;
  assign n16736 = ~n16735 | ~n16734;
  assign n16742 = ~n16741 | ~n16740;
  assign n16750 = ~n16745 & ~n16744;
  assign n16751 = ~n16750 & ~n16749;
  assign n16758 = ~n16752 | ~n16751;
  assign n16756 = ~n16753 | ~n16591;
  assign n16755 = ~n16754 | ~n16798;
  assign n16765 = n16758 & n16757;
  assign n16764 = ~n16766 & ~n16765;
  assign n16762 = ~n16759 & ~n16591;
  assign n16761 = ~n16760 & ~n16798;
  assign n16772 = ~n16764 & ~n16763;
  assign n16770 = ~n16766 | ~n16765;
  assign n16768 = ~n16782 | ~n16591;
  assign n16767 = ~n16783 | ~n16798;
  assign n16771 = ~n16770 | ~n16769;
  assign n16789 = ~n16772 & ~n16771;
  assign n16777 = ~n16773 | ~n16798;
  assign n16776 = ~n16775 | ~n16591;
  assign n16781 = ~n16778 & ~n16798;
  assign n16780 = ~n16779 & ~n16591;
  assign n16787 = ~n16791 | ~n16790;
  assign n16785 = ~n16782 | ~n16798;
  assign n16784 = ~n16783 | ~n16591;
  assign n16793 = ~n16789 & ~n16788;
  assign n16807 = ~n16793 & ~n16792;
  assign n16794 = ~n16809 | ~n16591;
  assign n16805 = ~n16797 | ~n16796;
  assign n16799 = ~n16801 & ~n16798;
  assign n16816 = ~n16800 & ~n16799;
  assign n16803 = ~n16802 | ~n16801;
  assign n16815 = n16805 & n16804;
  assign n16811 = ~n16808 | ~n16591;
  assign n16810 = ~n16809 | ~n16798;
  assign n16823 = ~n16828 | ~n16830;
  assign n16827 = ~n16823 | ~n16829;
  assign n16840 = ~n16827 | ~n16826;
  assign n16838 = ~n16833 & ~n16832;
  assign n16839 = ~n16838 & ~n16837;
  assign n16844 = ~n16840 | ~n16839;
  assign n16846 = ~n16844 | ~n16843;
  assign n16852 = ~n16850 | ~n16849;
  assign n16858 = ~n16852 & ~n16851;
  assign n16856 = ~n16854 | ~n16853;
  assign n16857 = ~n16856 & ~n16855;
  assign n16860 = ~n16858 | ~n16857;
  assign n16862 = ~n16860 & ~n16859;
  assign n16864 = ~n16862 | ~n16861;
  assign n16865 = ~n16864 & ~n16863;
  assign n16867 = ~n16866 | ~n16865;
  assign n16869 = ~n16868 & ~n16867;
  assign n16871 = ~n16870 | ~n16869;
  assign n16873 = ~n16872 & ~n16871;
  assign n16876 = ~n16874 | ~n16873;
  assign n16877 = ~n16876 & ~n16875;
  assign n16879 = ~n16878 | ~n16877;
  assign n16881 = ~n16880 & ~n16879;
  assign n16883 = ~n16882 | ~n16881;
  assign n16885 = ~n16884 & ~n16883;
  assign n16893 = ~n16892 & ~n16891;
  assign n16942 = ~n16916 & ~n16930;
  assign n16919 = ~n8926 & ~n16917;
  assign n16955 = ~n16922 | ~n16921;
  assign n16932 = ~n16924 | ~n16923;
  assign n16950 = ~n16932 | ~n16931;
  assign n16938 = ~n16950 | ~n16946;
  assign n16937 = ~n16947;
  assign n16945 = ~n16938 | ~n16937;
  assign n16941 = ~n8922 | ~n16939;
  assign n16953 = ~n16945 | ~n16944;
  assign n16951 = ~n16950 | ~n16949;
  assign n16954 = ~n16953 | ~n16952;
  assign n16959 = ~n15386 & ~n16958;
  assign n16965 = ~n16960 | ~n16959;
  assign n16963 = ~n16962 | ~n16961;
  assign n16964 = n16963 & P2_B_REG_SCAN_IN;
  assign n16966 = ~n16965 | ~n16964;
  assign n16969 = n16967 & n16966;
  assign n16968 = ~P2_STATE_REG_SCAN_IN & ~P2_B_REG_SCAN_IN;
  assign P2_U3296 = ~n16969 & ~n16968;
endmodule


