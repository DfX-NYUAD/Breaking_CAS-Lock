// Benchmark "b14_C_lock" written by ABC on Thu May 13 23:35:02 2021

module b14_C_lock ( 
    keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
    keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
    keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
    keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
    keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
    keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
    keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
    keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
    keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
    keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
    keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
    keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
    keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
    keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
    keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
    keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
    keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
    keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
    keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
    keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
    keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
    keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
    keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
    keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
    keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
    keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
    keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
    keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
    keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
    keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
    keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
    keyinput_156, keyinput_157, keyinput_158, keyinput_159, DATAI_28_,
    DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
    DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
    DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
    DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
    DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
    REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
    REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
    REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
    REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
    REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
    REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
    REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
    IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
    IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
    IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
    IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
    IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
    IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
    IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
    IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
    IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
    IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
    IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
    D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN,
    D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
    D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
    D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
    D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
    D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
    D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
    D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
    D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
    D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
    REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
    REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
    REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
    REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
    REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
    REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
    REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
    REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
    REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
    REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG1_REG_0__SCAN_IN,
    REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN,
    REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN,
    REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN,
    REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN,
    REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN,
    REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN,
    REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN,
    REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN,
    REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN,
    REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG2_REG_0__SCAN_IN,
    REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
    REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
    REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
    REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
    REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
    REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
    REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
    REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
    REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
    REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, B_REG_SCAN_IN,
    REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
    REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
    REG3_REG_22__SCAN_IN,
    U3217  );
  input  keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4,
    keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9,
    keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14,
    keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19,
    keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24,
    keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29,
    keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34,
    keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39,
    keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44,
    keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49,
    keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54,
    keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59,
    keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64,
    keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69,
    keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74,
    keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79,
    keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84,
    keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89,
    keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94,
    keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99,
    keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104,
    keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109,
    keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114,
    keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119,
    keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124,
    keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129,
    keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134,
    keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139,
    keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144,
    keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149,
    keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154,
    keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159,
    DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
    DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
    DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
    DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
    DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
    REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
    REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
    REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
    REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
    REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
    REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
    REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
    REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
    IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
    IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
    IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
    IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
    IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
    IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
    IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
    IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
    IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
    IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
    D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
    D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN,
    D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN,
    D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN,
    D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN,
    D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN,
    D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN,
    D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN,
    D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN,
    D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN,
    REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN,
    REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN,
    REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN,
    REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN,
    REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN,
    REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN,
    REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN,
    REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN,
    REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN,
    REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN,
    REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
    REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
    REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
    REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
    REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
    REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
    REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
    REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
    REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
    REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
    REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
    REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
    REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
    REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
    REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
    REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
    REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
    REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
    REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
    REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
    B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
    REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
    REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3217;
  wire n4324, n3178, n6252, n4145, n3755, n4879, n6067, n4223, n3421, n3460,
    n3262, n3179, n3180, n3181, n4692, n4928, n6066, n5993, n4701, n3275,
    n3682, n3395, n3229, n3452, n3438, n4675, n3688, n3252, n4402, n4004,
    n4175, n3759, n3223, n3258, n3254, n3692, n3248, n4367, n4067, n3285,
    n3332, n5924, n5700, n3689, n3246, n3242, n3894, n3872, n5536, n4005,
    n3224, n5534, n3888, n4089, n4090, n5673, n3219, n3218, n3410, n3420,
    n3251, n3250, n4169, n3263, n3475, n3467, n3196, n3241, n3951, n3932,
    n3225, n4078, n4152, n3606, n3566, n4552, n5963, n5831, n5471, n5145,
    n3203, n3204, n4361, n4343, n4360, n5407, n5275, n6476, n5600, n3207,
    n5103, n3220, n3334, n3335, n5369, n6288, n3317, n5666, n6020, n6559,
    n4505, n3274, n3273, n6216, n3852, n3685, n3687, n3683, n6208, n3586,
    n3228, n3350, n3388, n3245, n3468, n3466, n4748, n6369, n6248, n6477,
    n6472, n6385, n6299, n6365, n6358, n5943, n5676, n4876, n3436, n3413,
    n3425, n3602, n3264, n4501, n3720, n3719, n4511, n4504, n6215, n6168,
    n3686, n3684, n4495, n6211, n3355, n3186, n6460, n4369, n3187, n3666,
    n3905, n3188, n3216, n3189, n3190, n3459, n3191, n3192, n3193, n3194,
    n3195, n3222, n3197, n3198, n3255, n3199, n3637, n3200, n3201, n5741,
    n3202, n6465, n5869, n3206, n3208, n4932, n3212, n3213, n3214, n3215,
    n4575, n3217, n4220, n4405, n3221, n3718, n3226, n3227, n3588, n3349,
    n3446, n3265, n4084, n6553, n4602, n3237, n4094, n3257, n5186, n3260,
    n6568, n3887, n5870, n3623, n3633, n6300, n5744, n3378, n3482, n3249,
    n4203, n5763, n4339, n3358, n5864, n3593, n5701, n5525, n3401, n4317,
    n4282, n3722, n3756, n4237, n5738, n4213, n4854, n5162, n4398, n5861,
    n5809, n4284, n4506, n3757, n5265, n6563, n5768, n4503, n3400, n3499,
    n3522, n3506, n3539, n3371, n3340, n3316, n3582, n3632, n6243, n3615,
    n4189, n3294, n6473, n3277, n4261, n3658, n3669, n6545, n3244, n3243,
    n3515, n3247, n3253, n3709, n3256, n3259, n3261, n4497, n3272, n3267,
    n3266, n3270, n3268, n3269, n3271, n3469, n3276, n4370, n6428, n3284,
    n3279, n3278, n3282, n3280, n3281, n3283, n6296, n6375, n6314, n3292,
    n3287, n3286, n3290, n3288, n3289, n3291, n3293, n6487, n3301, n3296,
    n3295, n3299, n3297, n3298, n3300, n3302, n6388, n3308, n3310, n3569,
    n6340, n3309, n5647, n4573, n3312, n3311, n3315, n3313, n3314, n3320,
    n5750, n3318, n3319, n3321, n3326, n3337, n3322, n3323, n3324, n5900,
    n3325, n3328, n3327, n3331, n3329, n3330, n5678, n3333, n3336, n3339,
    n5732, n3338, n5465, n5468, n3342, n3341, n3347, n3345, n3343, n3344,
    n3346, n3348, n3354, n3366, n3351, n3352, n5559, n3353, n5594, n3357,
    n3356, n3364, n5607, n3359, n3362, n3360, n3361, n3363, n5460, n3365,
    n3368, n5428, n3367, n5446, n3370, n3369, n3377, n5582, n3372, n3375,
    n3373, n3374, n3376, n5604, n5490, n3380, n3379, n3385, n3383, n3381,
    n3382, n3384, n5441, n3386, n3393, n3387, n3389, n3390, n3391, n5378,
    n3392, n5361, n5483, n3394, n3397, n3491, n4805, n3396, n5045, n3399,
    n3398, n3407, n5097, n3402, n3405, n3403, n3404, n3406, n5152, n3408,
    n3409, n3412, n3411, n3414, n4745, n3417, n3415, n3416, n4777, n3418,
    n3419, n3423, n3422, n3424, n4765, n3426, n3428, n3427, n4778, n5007,
    n3431, n3430, n3432, n3434, n3433, n3435, n3437, n3440, n3439, n5025,
    n4240, n3443, n3442, n3449, n3444, n3447, n3445, n3448, n3450, n3456,
    n3451, n3453, n3454, n4830, n3455, n4880, n4902, n4947, n3458, n3457,
    n3464, n3462, n3461, n3463, n3465, n3471, n4720, n3470, n4912, n4925,
    n3474, n3479, n3476, n3477, n4818, n3478, n3933, n3481, n3480, n3487,
    n5079, n3485, n3483, n3484, n3486, n6019, n3490, n3496, n3492, n3493,
    n3494, n4864, n3495, n5119, n5155, n3498, n3497, n3504, n5142, n3502,
    n3500, n3501, n3503, n5194, n5327, n3508, n3507, n3513, n3511, n3509,
    n3510, n3512, n5271, n3514, n3519, n3529, n3516, n3517, n3547, n5171,
    n3518, n5237, n5340, n3521, n3520, n3527, n5315, n3525, n3523, n3524,
    n3526, n5328, n3528, n3531, n4988, n3530, n5277, n3538, n3537, n3545,
    n5412, n3540, n3543, n3541, n3542, n3544, n5487, n3546, n3551, n3548,
    n3549, n5222, n3550, n6024, n4016, n3562, n3561, n3565, n3563, n3564,
    n3568, n5945, n3567, n5817, n3570, n3571, n3572, n6411, n3575, n3573,
    n3574, n3579, n3577, n3578, n3581, n3580, n3584, n5868, n3583, n3585,
    n3592, n3587, n3589, n3590, n6520, n3591, n5810, n3594, n3601, n3596,
    n3595, n3599, n3597, n3598, n3600, n5865, n3603, n6572, n3605, n3604,
    n5981, n3613, n3608, n3607, n3611, n3609, n3610, n3612, n6260, n3614,
    n4426, n3622, n3617, n3616, n3620, n3618, n3619, n3621, n4449, n6360,
    n3630, n3625, n3624, n3628, n3626, n3627, n3629, n6246, n3631, n6251,
    n3641, n3635, n3634, n3639, n3636, n3638, n3640, n5780, n4346, n3665,
    n3660, n3659, n3663, n3661, n3662, n3664, n4347, n4278, n3670, n3677,
    n3672, n3671, n3675, n3673, n3674, n3676, n6556, n6204, n3695, n3690,
    n3691, n3693, n3694, n4703, n4546, n6106, n3712, n3710, n3711, n3714,
    n3713, n3715, n3717, n3716, n3721, n3723, n3725, n3724, n3731, n4540,
    n4539, n3729, n3727, n3726, n3728, n3730, n3747, n3733, n3732, n3737,
    n3735, n3734, n3736, n3745, n3739, n3738, n3743, n3741, n3740, n3742,
    n3744, n3746, n3752, n3749, n3748, n3750, n3751, n3753, n3754, n4151,
    n4272, n3758, n4176, n4547, n4031, n4080, n6247, n4120, n4328, n3875,
    n3853, n4553, U3149, n3873, n3874, n3876, n3878, n3877, n3893, n4749,
    n3892, n4142, n3880, n4677, n3879, n3886, n4671, n3885, n3883, n3881,
    n3882, n3884, n4672, n3890, n3889, n3891, n3896, n3895, n4235, n3898,
    n3897, n3899, n3903, n3901, n3900, n3902, n3904, n4234, n3907, n3906,
    n3908, n3911, n3910, n3909, n3912, n4885, n3913, n3914, n3926, n3916,
    n3915, n3917, n3920, n3919, n3918, n3921, n3927, n3923, n3922, n3924,
    n4931, n3925, n3928, n5081, n3930, n3929, n3931, n3936, n3935, n3934,
    n3937, n3941, n3939, n3938, n3940, n5080, n3942, n3949, n3944, n3943,
    n3945, n3948, n5095, n3947, n3946, n5094, n3950, n3953, n3952, n3954,
    n3957, n3956, n3955, n3958, n3962, n3960, n3959, n3961, n5146, n3964,
    n3963, n3965, n3968, n3967, n3966, n3969, n3973, n3971, n3970, n3972,
    n5274, n3974, n5332, n3976, n3975, n3977, n3980, n3979, n3978, n3981,
    n3985, n3983, n3982, n3984, n5331, n5335, n3987, n3986, n3988, n3992,
    n3990, n3989, n3991, n5404, n3993, n3995, n3994, n3996, n3999, n3998,
    n3997, n4000, n4002, n4001, n4003, n5491, n4007, n4006, n4008, n4011,
    n4010, n4009, n4012, n5533, n4015, n4014, n4013, n4018, n4017, n4019,
    n4027, n4021, n4020, n4028, n5597, n4023, n4022, n4024, n4036, n4026,
    n4025, n4037, n4403, n4030, n4029, n5598, n4044, n4033, n4032, n4034,
    n4043, n4035, n4039, n4038, n4041, n4040, n4042, n4045, n4047, n4046,
    n5669, n5742, n4049, n4048, n4050, n4053, n4052, n4051, n4054, n4056,
    n4055, n4058, n4371, n4057, n4059, n4062, n4061, n4060, n4063, n4065,
    n4064, n4066, n5947, n4069, n4068, n4070, n4073, n4072, n4071, n4074,
    n4076, n4075, n4077, n4079, n4419, n4082, n4081, n4083, n4088, n4086,
    n4085, n4087, n4420, n4092, n4091, n4093, n4130, n4096, n4095, n4129,
    n6347, n4098, n4097, n4099, n4126, n4101, n4100, n4127, n6350, n4131,
    n6353, n4103, n4102, n4104, n4107, n4106, n4193, n4105, n4108, n4133,
    n4110, n4109, n4111, n4196, n4113, n4112, n4114, n4135, n4116, n4115,
    n4136, n6459, n4118, n4117, n4119, n4123, n4122, n4121, n4124, n6463,
    n4140, n4156, n4125, n4141, n4128, n4132, n6348, n6354, n4183, n4134,
    n4197, n4139, n4137, n4138, n6461, n6467, n4158, n4144, n4143, n4146,
    n4247, n4148, n4147, n4248, n4155, n4150, n4174, n4170, n4172, n4153,
    n4159, n4334, n4162, n6219, n4165, n4166, n6366, n4171, n4173, n4178,
    n4177, n6486, n4249, n4338, n4252, n4251, n4253, n4257, n4255, n4254,
    n4256, n4342, n4336, n4379, n4326, n4325, n4327, n4332, n4330, n4329,
    n4331, n4333, n4362, n4335, n4344, n4337, n4340, n4341, n4364, n4363,
    n4377, n4366, n4365, n4368, n4375, n4373, n4372, n4374, n4376, n4378,
    n4389, n4381, n4380, n4383, n4382, n4387, n4385, n4384, n4386, n4388,
    U3217_Lock, input_0, input_1, AND_1, input_2, AND_2, input_3, AND_3,
    input_4, OR_4, input_5, AND_5, input_6, AND_6, input_7, OR_7, input_8,
    OR_8, input_9, OR_9, input_10, OR_10, input_11, AND_11, input_12,
    OR_12, input_13, OR_13, input_14, OR_14, input_15, AND_15, input_16,
    OR_16, input_17, AND_17, input_18, AND_18, input_19, AND_19, input_20,
    AND_20, input_21, AND_21, input_22, OR_22, input_23, OR_23, input_24,
    AND_24, input_25, OR_25, input_26, AND_26, input_27, AND_27, input_28,
    AND_28, input_29, OR_29, input_30, AND_30, input_31, OR_31, input_32,
    AND_32, input_33, AND_33, input_34, OR_34, input_35, OR_35, input_36,
    AND_36, input_37, AND_37, input_38, OR_38, input_39, AND_39, input_40,
    AND_40, input_41, OR_41, input_42, OR_42, input_43, AND_43, input_44,
    AND_44, input_45, OR_45, input_46, OR_46, input_47, OR_47, input_48,
    AND_48, input_49, OR_49, input_50, AND_50, input_51, OR_51, input_52,
    OR_52, input_53, OR_53, input_54, OR_54, input_55, AND_55, input_56,
    OR_56, input_57, AND_57, input_58, AND_58, input_59, OR_59, input_60,
    OR_60, input_61, OR_61, input_62, AND_62, input_63, OR_63, input_64,
    OR_64, input_65, OR_65, input_66, OR_66, input_67, OR_67, input_68,
    OR_68, input_69, AND_69, input_70, OR_70, input_71, OR_71, input_72,
    AND_72, input_73, OR_73, input_74, OR_74, input_75, AND_75, input_76,
    OR_76, input_77, OR_77, input_78, OR_78, input_79, OR_79, input_80,
    input_81, AND_81, input_82, AND_82, input_83, AND_83, input_84, OR_84,
    input_85, AND_85, input_86, AND_86, input_87, OR_87, input_88, OR_88,
    input_89, OR_89, input_90, OR_90, input_91, AND_91, input_92, OR_92,
    input_93, OR_93, input_94, OR_94, input_95, AND_95, input_96, OR_96,
    input_97, AND_97, input_98, AND_98, input_99, AND_99, input_100,
    AND_100, input_101, AND_101, input_102, OR_102, input_103, OR_103,
    input_104, AND_104, input_105, OR_105, input_106, AND_106, input_107,
    AND_107, input_108, AND_108, input_109, OR_109, input_110, AND_110,
    input_111, OR_111, input_112, AND_112, input_113, AND_113, input_114,
    OR_114, input_115, OR_115, input_116, AND_116, input_117, AND_117,
    input_118, OR_118, input_119, AND_119, input_120, AND_120, input_121,
    OR_121, input_122, OR_122, input_123, AND_123, input_124, AND_124,
    input_125, OR_125, input_126, OR_126, input_127, OR_127, input_128,
    AND_128, input_129, OR_129, input_130, AND_130, input_131, OR_131,
    input_132, OR_132, input_133, OR_133, input_134, OR_134, input_135,
    AND_135, input_136, OR_136, input_137, AND_137, input_138, AND_138,
    input_139, OR_139, input_140, OR_140, input_141, OR_141, input_142,
    AND_142, input_143, OR_143, input_144, OR_144, input_145, OR_145,
    input_146, OR_146, input_147, OR_147, input_148, OR_148, input_149,
    AND_149, input_150, OR_150, input_151, OR_151, input_152, AND_152,
    input_153, OR_153, input_154, OR_154, input_155, AND_155, input_156,
    OR_156, input_157, OR_157, input_158, OR_158, input_159, OR_159,
    OR_159_INV, CASOP;
  assign n4324 = ~n4317 | ~n4175;
  assign n3178 = ~n6465;
  assign n6252 = ~n4170 & ~n4153;
  assign n4145 = ~n4367;
  assign n3755 = ~IR_REG_31__SCAN_IN;
  assign n4879 = ~n3464 | ~n3463;
  assign n6067 = ~n3413 | ~n3189;
  assign n4223 = ~n3264 ^ IR_REG_29__SCAN_IN;
  assign n3421 = n4220 & n4223;
  assign n3460 = ~n4575;
  assign n3262 = ~n4497 | ~IR_REG_31__SCAN_IN;
  assign n3179 = ~n3421;
  assign n3180 = ~n3179;
  assign n3181 = ~n3179;
  assign n4692 = ~n3452 ^ IR_REG_2__SCAN_IN;
  assign n4928 = ~n3449 | ~n3448;
  assign n6066 = ~n4777;
  assign n5993 = ~n3666;
  assign n4701 = ~n3275 ^ n3260;
  assign n3275 = ~n3190 | ~IR_REG_31__SCAN_IN;
  assign n3682 = ~n3251 | ~n3192;
  assign n3395 = ~n3244 & ~n3243;
  assign n3229 = n3186 & n3191;
  assign n3452 = n3755 | n3438;
  assign n3438 = ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN;
  assign n4675 = ~n3274 ^ n3222;
  assign n3688 = ~n3682 & ~n3253;
  assign n3252 = ~IR_REG_19__SCAN_IN & ~IR_REG_20__SCAN_IN;
  assign n4402 = ~n5600 | ~n5597;
  assign n4004 = n3999 | n4000;
  assign n4175 = ~n3759 | ~n4501;
  assign n3759 = n4511 & n4504;
  assign n3223 = ~IR_REG_24__SCAN_IN & ~n3259;
  assign n3258 = ~IR_REG_25__SCAN_IN;
  assign n3254 = ~IR_REG_22__SCAN_IN & ~IR_REG_23__SCAN_IN;
  assign n3692 = ~n3688;
  assign n3248 = ~IR_REG_13__SCAN_IN;
  assign n4367 = ~n4317 | ~n3853;
  assign n4067 = n4062 | n4063;
  assign n3285 = ~n3294 & ~n6473;
  assign n3332 = ~n3340 & ~n4398;
  assign n5924 = ~n6369;
  assign n5700 = ~n3695 & ~n3694;
  assign n3689 = ~IR_REG_22__SCAN_IN;
  assign n3246 = ~IR_REG_10__SCAN_IN & ~IR_REG_11__SCAN_IN;
  assign n3242 = ~IR_REG_5__SCAN_IN;
  assign n3894 = ~n3874 ^ n4367;
  assign n3872 = n6066 | n4324;
  assign n5536 = ~n4005 | ~n4004;
  assign n4005 = ~n3225 | ~n3198;
  assign n3224 = ~n3993;
  assign n5534 = n4014 | n4013;
  assign n3888 = ~n3887 & ~n3886;
  assign n4089 = n4088 | n4087;
  assign n4090 = n4419 | n4420;
  assign n5673 = ~n3219 | ~n3220;
  assign n3219 = n3221 & n3199;
  assign n3218 = n3217 & n4220;
  assign n3410 = n3637 | n3408;
  assign n3420 = n3637 | n3418;
  assign n3251 = ~n3588;
  assign n3250 = ~IR_REG_18__SCAN_IN;
  assign n4169 = ~n4552 & ~n4547;
  assign n3263 = n3256 & n3195;
  assign n3475 = IR_REG_31__SCAN_IN & n3467;
  assign n3467 = IR_REG_3__SCAN_IN | n3466;
  assign n3196 = n4317 | n4213;
  assign n3241 = ~IR_REG_2__SCAN_IN & ~IR_REG_3__SCAN_IN;
  assign n3951 = n5095 | n5094;
  assign n3932 = ~n4324 & ~n3876;
  assign n3225 = ~n5335 | ~n3226;
  assign n4078 = n4073 | n4074;
  assign n4152 = n6168 & n6215;
  assign n3606 = ~n3615 & ~n4189;
  assign n3566 = ~n3316 & ~n3317;
  assign n4552 = n6168 | n6215;
  assign n5963 = ~n4203;
  assign n5831 = ~n5864;
  assign n5471 = ~n5465;
  assign n5145 = ~n3951 | ~n3203;
  assign n3203 = ~n3204 & ~n5146;
  assign n3204 = ~n3950;
  assign n4361 = ~n4344 | ~n4343;
  assign n4343 = n4342 | n4341;
  assign n4360 = ~n4333 & ~n4362;
  assign n5407 = ~n6024;
  assign n5275 = ~n5145 | ~n3962;
  assign n6476 = n5993 | n3302;
  assign n5600 = n4015 & n5534;
  assign n3207 = n3208 & n4067;
  assign n5103 = ~n5045;
  assign n3220 = ~n4405 | ~n4045;
  assign n3334 = n3180 & n3333;
  assign n3335 = n3331 | n3330;
  assign n5369 = ~REG3_REG_12__SCAN_IN;
  assign n6288 = ~n6300;
  assign n3317 = ~REG3_REG_16__SCAN_IN;
  assign n5666 = ~n3326 | ~n3325;
  assign n6020 = ~n3933;
  assign n6559 = ~n4546 | ~n6106;
  assign n4505 = n4503 & n4175;
  assign n3274 = ~n3273 | ~IR_REG_31__SCAN_IN;
  assign n3273 = ~n3256 | ~n3188;
  assign n6216 = IR_REG_23__SCAN_IN ^ n3757;
  assign n3852 = n3756 | n3693;
  assign n3685 = ~IR_REG_21__SCAN_IN;
  assign n3687 = n3683 & IR_REG_31__SCAN_IN;
  assign n3683 = n3682 | IR_REG_19__SCAN_IN;
  assign n6208 = ~n3687 ^ IR_REG_20__SCAN_IN;
  assign n3586 = ~IR_REG_16__SCAN_IN & ~IR_REG_17__SCAN_IN;
  assign n3228 = n3229 & n3249;
  assign n3350 = ~IR_REG_12__SCAN_IN;
  assign n3388 = ~IR_REG_8__SCAN_IN & ~IR_REG_9__SCAN_IN;
  assign n3245 = ~IR_REG_6__SCAN_IN & ~IR_REG_7__SCAN_IN;
  assign n3468 = ~IR_REG_4__SCAN_IN;
  assign n3466 = n3453 & IR_REG_31__SCAN_IN;
  assign n4748 = n3890 & n3889;
  assign n6369 = n5993 | n3631;
  assign n6248 = ~n5809 | ~n4171;
  assign n6477 = ~n6248;
  assign n6472 = ~n4165 | ~n4703;
  assign n6385 = ~n3292 | ~n3291;
  assign n6299 = ~n3301 | ~n3300;
  assign n6365 = ~n3622 | ~n3621;
  assign n6358 = ~n3641 | ~n3640;
  assign n5943 = ~n3320 | ~n3319;
  assign n5676 = ~n3347 | ~n3346;
  assign n4876 = ~n3436 | ~n3435;
  assign n3436 = n3431 & n3430;
  assign n3413 = n3410 & n3409;
  assign n3425 = n3420 & n3419;
  assign n3602 = ~IR_REG_19__SCAN_IN;
  assign n3264 = n3263 | n3755;
  assign n4501 = ~n3720 ^ IR_REG_26__SCAN_IN;
  assign n3720 = ~n3719 | ~IR_REG_31__SCAN_IN;
  assign n3719 = n3718 | IR_REG_25__SCAN_IN;
  assign n4511 = ~n3711 ^ IR_REG_25__SCAN_IN;
  assign n4504 = ~n3712 ^ IR_REG_24__SCAN_IN;
  assign n6215 = ~n3852;
  assign n6168 = ~n3686 ^ n3685;
  assign n3686 = ~n3684 & ~n3755;
  assign n3684 = ~IR_REG_20__SCAN_IN & ~n3687;
  assign n4495 = ~STATE_REG_SCAN_IN;
  assign n6211 = ~n6572;
  assign n3355 = ~n3459;
  assign n3186 = n3388 & n3246;
  assign n6460 = ~n4090 | ~n4089;
  assign n4369 = ~n3196;
  assign n3187 = n3200 & n5947;
  assign n3666 = ~n3469;
  assign n3905 = n3903 | n3902;
  assign n3188 = n3223 & n3260;
  assign n3216 = ~n4223;
  assign n3189 = ~n3412 & ~n3218;
  assign n3190 = ~n3256 | ~n3223;
  assign n3459 = n3265 & n4223;
  assign n3191 = n3248 & n3350;
  assign n3192 = n3586 & n3250;
  assign n3193 = n3221 & n4040;
  assign n3194 = n3905 & n4885;
  assign n3195 = n3188 & n3222;
  assign n3222 = ~IR_REG_28__SCAN_IN;
  assign n3197 = ~n4334 & ~n4342;
  assign n3198 = ~n3224 & ~n5491;
  assign n3255 = ~IR_REG_24__SCAN_IN;
  assign n3199 = n4040 & n5669;
  assign n3637 = ~n3265 | ~n3216;
  assign n3200 = ~n4056 | ~n4055;
  assign n3201 = n4135 ^ n4136;
  assign n5741 = ~n4053 ^ n4054;
  assign n3202 = n3247 & n3229;
  assign n6465 = ~n6252;
  assign n5869 = ~n3206 | ~n3207;
  assign n3206 = ~n5742 | ~n3187;
  assign n3208 = ~n3187 | ~n5741;
  assign n4932 = ~n3212 | ~n3914;
  assign n3212 = ~n3213 | ~n3194;
  assign n3213 = ~n3215 | ~n3214;
  assign n3214 = ~n4234;
  assign n3215 = ~n4235;
  assign n4575 = ~n3216 | ~n4220;
  assign n3217 = ~n4223 & ~n3411;
  assign n4220 = ~n3262 ^ IR_REG_30__SCAN_IN;
  assign n4405 = ~n4402 | ~n4044;
  assign n3221 = ~n4402 | ~n4035;
  assign n3718 = ~n3256 | ~n3255;
  assign n3226 = ~n5404 & ~n3227;
  assign n3227 = ~n3985;
  assign n3588 = ~n3247 | ~n3228;
  assign n3349 = ~n3247 | ~n3186;
  assign n3446 = n4575 | n3445;
  assign n3265 = ~n4220;
  assign n4084 = ~n4094;
  assign n6553 = ~n4602;
  assign n4602 = ~n5700;
  assign n3237 = ~n4133 | ~n4111;
  assign n4094 = ~n3932;
  assign n3257 = ~IR_REG_26__SCAN_IN;
  assign n5186 = ~n5277;
  assign n3260 = ~IR_REG_27__SCAN_IN;
  assign n6568 = ~n4370;
  assign n3887 = ~n3880 | ~n3879;
  assign n5870 = n4078 & n4077;
  assign n3623 = ~n3632 & ~n6243;
  assign n3633 = ~n3355;
  assign n6300 = n5993 | n3293;
  assign n5744 = ~n5647;
  assign n3378 = ~n3539 & ~n5162;
  assign n3482 = REG3_REG_3__SCAN_IN & REG3_REG_4__SCAN_IN;
  assign n3249 = ~IR_REG_14__SCAN_IN & ~IR_REG_15__SCAN_IN;
  assign n4203 = n3469 | n3614;
  assign n5763 = ~n3605 | ~n3604;
  assign n4339 = n4159 | n4158;
  assign n3358 = ~n3371 & ~n5369;
  assign n5864 = ~n3592 | ~n3591;
  assign n3593 = ~n3582 & ~n5861;
  assign n5701 = ~n3575 | ~n3574;
  assign n5525 = ~n5446;
  assign n3401 = ~REG3_REG_6__SCAN_IN;
  assign n4317 = ~n6168 | ~n6208;
  assign n4282 = ~n3725 & ~n3724;
  assign n3722 = ~n4501 & ~n4504;
  assign n3756 = n3690 & n3689;
  assign n4237 = ~n4178 & ~n4177;
  assign n5738 = ~n3335 & ~n3334;
  assign n4213 = ~n4175;
  assign n4854 = ~REG3_REG_8__SCAN_IN;
  assign n5162 = ~REG3_REG_10__SCAN_IN;
  assign n4398 = ~REG3_REG_14__SCAN_IN;
  assign n5861 = ~REG3_REG_18__SCAN_IN;
  assign n5809 = ~n4505 | ~n4169;
  assign n4284 = ~n3723 & ~n3722;
  assign n4506 = ~n3721 | ~n4501;
  assign n3757 = ~n3756 & ~n3755;
  assign n5265 = ~n3272 | ~n3271;
  assign n6563 = ~n3665 | ~n3664;
  assign n5768 = ~n3584 | ~n3583;
  assign n4503 = ~n6216 & ~n4495;
  assign n3400 = ~n3482 | ~REG3_REG_5__SCAN_IN;
  assign n3499 = ~n3400 & ~n3401;
  assign n3522 = ~n3499 | ~REG3_REG_7__SCAN_IN;
  assign n3506 = ~n3522 & ~n4854;
  assign n3539 = ~n3506 | ~REG3_REG_9__SCAN_IN;
  assign n3371 = ~n3378 | ~REG3_REG_11__SCAN_IN;
  assign n3340 = ~n3358 | ~REG3_REG_13__SCAN_IN;
  assign n3316 = ~n3332 | ~REG3_REG_15__SCAN_IN;
  assign n3582 = ~n3566 | ~REG3_REG_17__SCAN_IN;
  assign n3632 = ~n3593 | ~REG3_REG_19__SCAN_IN;
  assign n6243 = ~REG3_REG_20__SCAN_IN;
  assign n3615 = ~n3623 | ~REG3_REG_21__SCAN_IN;
  assign n4189 = ~REG3_REG_22__SCAN_IN;
  assign n3294 = ~n3606 | ~REG3_REG_23__SCAN_IN;
  assign n6473 = ~REG3_REG_24__SCAN_IN;
  assign n3277 = ~n3285 | ~REG3_REG_25__SCAN_IN;
  assign n4261 = ~REG3_REG_26__SCAN_IN;
  assign n3658 = ~n3277 & ~n4261;
  assign n3669 = n3658 & REG3_REG_27__SCAN_IN;
  assign n6545 = REG3_REG_28__SCAN_IN ^ n3669;
  assign n3244 = ~n3438 | ~n3241;
  assign n3243 = ~n3468 | ~n3242;
  assign n3515 = ~n3395 | ~n3245;
  assign n3247 = ~n3515;
  assign n3253 = ~n3252 | ~n3685;
  assign n3709 = ~n3688 | ~n3254;
  assign n3256 = ~n3709;
  assign n3259 = ~n3258 | ~n3257;
  assign n3261 = ~IR_REG_29__SCAN_IN;
  assign n4497 = ~n3263 | ~n3261;
  assign n3272 = ~n6545 | ~n3181;
  assign n3267 = ~n4573 | ~REG0_REG_28__SCAN_IN;
  assign n3266 = ~n3633 | ~REG1_REG_28__SCAN_IN;
  assign n3270 = ~n3267 | ~n3266;
  assign n3268 = ~REG2_REG_28__SCAN_IN;
  assign n3269 = ~n4575 & ~n3268;
  assign n3271 = ~n3270 & ~n3269;
  assign n3469 = n4675 & n4701;
  assign n3276 = ~DATAI_28_;
  assign n4370 = ~n3469 & ~n3276;
  assign n6428 = n4261 ^ n3277;
  assign n3284 = ~n6428 | ~n3181;
  assign n3279 = ~n4573 | ~REG0_REG_26__SCAN_IN;
  assign n3278 = ~n3633 | ~REG1_REG_26__SCAN_IN;
  assign n3282 = ~n3279 | ~n3278;
  assign n3280 = ~REG2_REG_26__SCAN_IN;
  assign n3281 = ~n4575 & ~n3280;
  assign n3283 = ~n3282 & ~n3281;
  assign n6296 = ~n3284 | ~n3283;
  assign n6375 = ~n3666 | ~DATAI_26_;
  assign n6314 = REG3_REG_25__SCAN_IN ^ n3285;
  assign n3292 = ~n6314 | ~n3180;
  assign n3287 = ~n4573 | ~REG0_REG_25__SCAN_IN;
  assign n3286 = ~n3633 | ~REG1_REG_25__SCAN_IN;
  assign n3290 = ~n3287 | ~n3286;
  assign n3288 = ~REG2_REG_25__SCAN_IN;
  assign n3289 = ~n4575 & ~n3288;
  assign n3291 = ~n3290 & ~n3289;
  assign n3293 = ~DATAI_25_;
  assign n6487 = n6473 ^ n3294;
  assign n3301 = ~n6487 | ~n3181;
  assign n3296 = ~n4573 | ~REG0_REG_24__SCAN_IN;
  assign n3295 = ~n3633 | ~REG1_REG_24__SCAN_IN;
  assign n3299 = ~n3296 | ~n3295;
  assign n3297 = ~REG2_REG_24__SCAN_IN;
  assign n3298 = ~n4575 & ~n3297;
  assign n3300 = ~n3299 & ~n3298;
  assign n3302 = ~DATAI_24_;
  assign n6388 = ~n6375;
  assign n3308 = ~DATAI_16_;
  assign n3310 = n3469 | n3308;
  assign n3569 = ~n3588 | ~IR_REG_31__SCAN_IN;
  assign n6340 = ~n3569 ^ IR_REG_16__SCAN_IN;
  assign n3309 = ~n3469 | ~n6340;
  assign n5647 = ~n3310 | ~n3309;
  assign n4573 = ~n3637;
  assign n3312 = ~n4573 | ~REG0_REG_16__SCAN_IN;
  assign n3311 = ~n3633 | ~REG1_REG_16__SCAN_IN;
  assign n3315 = ~n3312 | ~n3311;
  assign n3313 = ~REG2_REG_16__SCAN_IN;
  assign n3314 = ~n4575 & ~n3313;
  assign n3320 = ~n3315 & ~n3314;
  assign n5750 = ~n3317 ^ n3316;
  assign n3318 = ~n5750;
  assign n3319 = ~n3180 | ~n3318;
  assign n3321 = ~DATAI_15_;
  assign n3326 = n5993 | n3321;
  assign n3337 = n3202 | n3755;
  assign n3322 = ~n3337;
  assign n3323 = ~n3322 & ~IR_REG_14__SCAN_IN;
  assign n3324 = ~n3323 & ~n3755;
  assign n5900 = IR_REG_15__SCAN_IN ^ n3324;
  assign n3325 = ~n5993 | ~n5900;
  assign n3328 = ~n4573 | ~REG0_REG_15__SCAN_IN;
  assign n3327 = ~n3633 | ~REG1_REG_15__SCAN_IN;
  assign n3331 = ~n3328 | ~n3327;
  assign n3329 = ~REG2_REG_15__SCAN_IN;
  assign n3330 = ~n4575 & ~n3329;
  assign n5678 = ~REG3_REG_15__SCAN_IN ^ n3332;
  assign n3333 = ~n5678;
  assign n3336 = ~DATAI_14_;
  assign n3339 = n5993 | n3336;
  assign n5732 = ~n3337 ^ IR_REG_14__SCAN_IN;
  assign n3338 = ~n5993 | ~n5732;
  assign n5465 = ~n3339 | ~n3338;
  assign n5468 = n4398 ^ n3340;
  assign n3342 = ~n3181 | ~n5468;
  assign n3341 = ~n4573 | ~REG0_REG_14__SCAN_IN;
  assign n3347 = n3342 & n3341;
  assign n3345 = ~n3633 | ~REG1_REG_14__SCAN_IN;
  assign n3343 = ~REG2_REG_14__SCAN_IN;
  assign n3344 = n4575 | n3343;
  assign n3346 = n3345 & n3344;
  assign n3348 = ~DATAI_13_;
  assign n3354 = n5993 | n3348;
  assign n3366 = ~n3349 | ~IR_REG_31__SCAN_IN;
  assign n3351 = n3366 & n3350;
  assign n3352 = ~n3351 & ~n3755;
  assign n5559 = IR_REG_13__SCAN_IN ^ n3352;
  assign n3353 = ~n5993 | ~n5559;
  assign n5594 = ~n3354 | ~n3353;
  assign n3357 = ~n4573 | ~REG0_REG_13__SCAN_IN;
  assign n3356 = ~n3633 | ~REG1_REG_13__SCAN_IN;
  assign n3364 = n3357 & n3356;
  assign n5607 = ~REG3_REG_13__SCAN_IN ^ n3358;
  assign n3359 = ~n5607;
  assign n3362 = ~n3181 | ~n3359;
  assign n3360 = ~REG2_REG_13__SCAN_IN;
  assign n3361 = n4575 | n3360;
  assign n3363 = n3362 & n3361;
  assign n5460 = ~n3364 | ~n3363;
  assign n3365 = ~DATAI_12_;
  assign n3368 = n5993 | n3365;
  assign n5428 = ~n3366 ^ IR_REG_12__SCAN_IN;
  assign n3367 = ~n5993 | ~n5428;
  assign n5446 = ~n3368 | ~n3367;
  assign n3370 = ~n4573 | ~REG0_REG_12__SCAN_IN;
  assign n3369 = ~n3633 | ~REG1_REG_12__SCAN_IN;
  assign n3377 = n3370 & n3369;
  assign n5582 = ~n5369 ^ n3371;
  assign n3372 = ~n5582;
  assign n3375 = ~n3181 | ~n3372;
  assign n3373 = ~REG2_REG_12__SCAN_IN;
  assign n3374 = n4575 | n3373;
  assign n3376 = n3375 & n3374;
  assign n5604 = ~n3377 | ~n3376;
  assign n5490 = REG3_REG_11__SCAN_IN ^ n3378;
  assign n3380 = ~n3181 | ~n5490;
  assign n3379 = ~n3633 | ~REG1_REG_11__SCAN_IN;
  assign n3385 = n3380 & n3379;
  assign n3383 = ~n4573 | ~REG0_REG_11__SCAN_IN;
  assign n3381 = ~REG2_REG_11__SCAN_IN;
  assign n3382 = n4575 | n3381;
  assign n3384 = n3383 & n3382;
  assign n5441 = ~n3385 | ~n3384;
  assign n3386 = ~DATAI_11_;
  assign n3393 = n5993 | n3386;
  assign n3387 = ~IR_REG_10__SCAN_IN;
  assign n3389 = ~n3388 | ~n3387;
  assign n3390 = n3515 | n3389;
  assign n3391 = ~n3390 | ~IR_REG_31__SCAN_IN;
  assign n5378 = ~n3391 ^ IR_REG_11__SCAN_IN;
  assign n3392 = ~n5993 | ~n5378;
  assign n5361 = ~n3393 | ~n3392;
  assign n5483 = ~n5361;
  assign n3394 = ~DATAI_6_;
  assign n3397 = n5993 | n3394;
  assign n3491 = n3395 | n3755;
  assign n4805 = ~n3491 ^ IR_REG_6__SCAN_IN;
  assign n3396 = ~n5993 | ~n4805;
  assign n5045 = ~n3397 | ~n3396;
  assign n3399 = ~n4573 | ~REG0_REG_6__SCAN_IN;
  assign n3398 = ~n3459 | ~REG1_REG_6__SCAN_IN;
  assign n3407 = n3399 & n3398;
  assign n5097 = ~n3401 ^ n3400;
  assign n3402 = ~n5097;
  assign n3405 = ~n3180 | ~n3402;
  assign n3403 = ~REG2_REG_6__SCAN_IN;
  assign n3404 = n4575 | n3403;
  assign n3406 = n3405 & n3404;
  assign n5152 = ~n3407 | ~n3406;
  assign n3408 = ~REG0_REG_1__SCAN_IN;
  assign n3409 = ~n3459 | ~REG1_REG_1__SCAN_IN;
  assign n3412 = n3421 & REG3_REG_1__SCAN_IN;
  assign n3411 = ~REG2_REG_1__SCAN_IN;
  assign n3414 = ~IR_REG_31__SCAN_IN | ~IR_REG_0__SCAN_IN;
  assign n4745 = ~n3414 ^ IR_REG_1__SCAN_IN;
  assign n3417 = ~n3469 | ~n4745;
  assign n3415 = ~DATAI_1_;
  assign n3416 = n3469 | n3415;
  assign n4777 = ~n3417 | ~n3416;
  assign n3418 = ~REG0_REG_0__SCAN_IN;
  assign n3419 = ~n3459 | ~REG1_REG_0__SCAN_IN;
  assign n3423 = ~n3421 | ~REG3_REG_0__SCAN_IN;
  assign n3422 = ~n3460 | ~REG2_REG_0__SCAN_IN;
  assign n3424 = n3423 & n3422;
  assign n4765 = ~n3425 | ~n3424;
  assign n3426 = ~DATAI_0_;
  assign n3428 = n3469 | n3426;
  assign n3427 = ~n3469 | ~IR_REG_0__SCAN_IN;
  assign n4778 = ~n3428 | ~n3427;
  assign n5007 = ~n4778;
  assign n3431 = ~n3460 | ~REG2_REG_2__SCAN_IN;
  assign n3430 = ~n3459 | ~REG1_REG_2__SCAN_IN;
  assign n3432 = ~REG0_REG_2__SCAN_IN;
  assign n3434 = n3637 | n3432;
  assign n3433 = ~n3421 | ~REG3_REG_2__SCAN_IN;
  assign n3435 = n3434 & n3433;
  assign n3437 = ~DATAI_2_;
  assign n3440 = n3469 | n3437;
  assign n3439 = ~n3469 | ~n4692;
  assign n5025 = ~n3440 | ~n3439;
  assign n4240 = ~n5025;
  assign n3443 = ~n4573 | ~REG0_REG_3__SCAN_IN;
  assign n3442 = ~n3459 | ~REG1_REG_3__SCAN_IN;
  assign n3449 = n3443 & n3442;
  assign n3444 = ~REG3_REG_3__SCAN_IN;
  assign n3447 = ~n3421 | ~n3444;
  assign n3445 = ~REG2_REG_3__SCAN_IN;
  assign n3448 = n3447 & n3446;
  assign n3450 = ~DATAI_3_;
  assign n3456 = n3469 | n3450;
  assign n3451 = ~IR_REG_2__SCAN_IN;
  assign n3453 = ~n3452 | ~n3451;
  assign n3454 = ~IR_REG_3__SCAN_IN;
  assign n4830 = ~n3466 ^ n3454;
  assign n3455 = ~n3469 | ~n4830;
  assign n4880 = ~n3456 | ~n3455;
  assign n4902 = ~n4880;
  assign n4947 = REG3_REG_3__SCAN_IN ^ REG3_REG_4__SCAN_IN;
  assign n3458 = ~n3180 | ~n4947;
  assign n3457 = ~n4573 | ~REG0_REG_4__SCAN_IN;
  assign n3464 = n3458 & n3457;
  assign n3462 = ~n3459 | ~REG1_REG_4__SCAN_IN;
  assign n3461 = ~n3460 | ~REG2_REG_4__SCAN_IN;
  assign n3463 = n3462 & n3461;
  assign n3465 = ~DATAI_4_;
  assign n3471 = n3469 | n3465;
  assign n4720 = ~n3475 ^ n3468;
  assign n3470 = ~n3469 | ~n4720;
  assign n4912 = ~n3471 | ~n3470;
  assign n4925 = ~n4912;
  assign n3474 = ~DATAI_5_;
  assign n3479 = n5993 | n3474;
  assign n3476 = ~IR_REG_4__SCAN_IN & ~n3475;
  assign n3477 = ~n3476 & ~n3755;
  assign n4818 = IR_REG_5__SCAN_IN ^ n3477;
  assign n3478 = ~n5993 | ~n4818;
  assign n3933 = ~n3479 | ~n3478;
  assign n3481 = ~n4573 | ~REG0_REG_5__SCAN_IN;
  assign n3480 = ~n3459 | ~REG1_REG_5__SCAN_IN;
  assign n3487 = n3481 & n3480;
  assign n5079 = REG3_REG_5__SCAN_IN ^ n3482;
  assign n3485 = ~n3421 | ~n5079;
  assign n3483 = ~REG2_REG_5__SCAN_IN;
  assign n3484 = n4575 | n3483;
  assign n3486 = n3485 & n3484;
  assign n6019 = ~n3487 | ~n3486;
  assign n3490 = ~DATAI_7_;
  assign n3496 = n5993 | n3490;
  assign n3492 = ~n3491;
  assign n3493 = ~n3492 & ~IR_REG_6__SCAN_IN;
  assign n3494 = ~n3493 & ~n3755;
  assign n4864 = IR_REG_7__SCAN_IN ^ n3494;
  assign n3495 = ~n5993 | ~n4864;
  assign n5119 = ~n3496 | ~n3495;
  assign n5155 = ~n5119;
  assign n3498 = ~n4573 | ~REG0_REG_7__SCAN_IN;
  assign n3497 = ~n3459 | ~REG1_REG_7__SCAN_IN;
  assign n3504 = n3498 & n3497;
  assign n5142 = REG3_REG_7__SCAN_IN ^ n3499;
  assign n3502 = ~n3181 | ~n5142;
  assign n3500 = ~REG2_REG_7__SCAN_IN;
  assign n3501 = n4575 | n3500;
  assign n3503 = n3502 & n3501;
  assign n5194 = ~n3504 | ~n3503;
  assign n5327 = REG3_REG_9__SCAN_IN ^ n3506;
  assign n3508 = ~n3181 | ~n5327;
  assign n3507 = ~n3633 | ~REG1_REG_9__SCAN_IN;
  assign n3513 = n3508 & n3507;
  assign n3511 = ~n4573 | ~REG0_REG_9__SCAN_IN;
  assign n3509 = ~REG2_REG_9__SCAN_IN;
  assign n3510 = n4575 | n3509;
  assign n3512 = n3511 & n3510;
  assign n5271 = ~n3513 | ~n3512;
  assign n3514 = ~DATAI_9_;
  assign n3519 = n5993 | n3514;
  assign n3529 = ~n3515 | ~IR_REG_31__SCAN_IN;
  assign n3516 = ~n3529;
  assign n3517 = ~n3516 & ~IR_REG_8__SCAN_IN;
  assign n3547 = ~n3517 & ~n3755;
  assign n5171 = IR_REG_9__SCAN_IN ^ n3547;
  assign n3518 = ~n5993 | ~n5171;
  assign n5237 = ~n3519 | ~n3518;
  assign n5340 = ~n5237;
  assign n3521 = ~n4573 | ~REG0_REG_8__SCAN_IN;
  assign n3520 = ~n3633 | ~REG1_REG_8__SCAN_IN;
  assign n3527 = n3521 & n3520;
  assign n5315 = n4854 ^ n3522;
  assign n3525 = ~n3181 | ~n5315;
  assign n3523 = ~REG2_REG_8__SCAN_IN;
  assign n3524 = n4575 | n3523;
  assign n3526 = n3525 & n3524;
  assign n5328 = ~n3527 | ~n3526;
  assign n3528 = ~DATAI_8_;
  assign n3531 = n5993 | n3528;
  assign n4988 = ~n3529 ^ IR_REG_8__SCAN_IN;
  assign n3530 = ~n5993 | ~n4988;
  assign n5277 = ~n3531 | ~n3530;
  assign n3538 = ~n4573 | ~REG0_REG_10__SCAN_IN;
  assign n3537 = ~n3633 | ~REG1_REG_10__SCAN_IN;
  assign n3545 = n3538 & n3537;
  assign n5412 = ~n5162 ^ n3539;
  assign n3540 = ~n5412;
  assign n3543 = ~n3181 | ~n3540;
  assign n3541 = ~REG2_REG_10__SCAN_IN;
  assign n3542 = n4575 | n3541;
  assign n3544 = n3543 & n3542;
  assign n5487 = ~n3545 | ~n3544;
  assign n3546 = ~DATAI_10_;
  assign n3551 = n5993 | n3546;
  assign n3548 = ~IR_REG_9__SCAN_IN & ~n3547;
  assign n3549 = ~n3548 & ~n3755;
  assign n5222 = IR_REG_10__SCAN_IN ^ n3549;
  assign n3550 = ~n5993 | ~n5222;
  assign n6024 = ~n3551 | ~n3550;
  assign n4016 = ~n5594;
  assign n3562 = ~n4573 | ~REG0_REG_17__SCAN_IN;
  assign n3561 = ~n3633 | ~REG1_REG_17__SCAN_IN;
  assign n3565 = ~n3562 | ~n3561;
  assign n3563 = ~REG2_REG_17__SCAN_IN;
  assign n3564 = ~n4575 & ~n3563;
  assign n3568 = ~n3565 & ~n3564;
  assign n5945 = REG3_REG_17__SCAN_IN ^ n3566;
  assign n3567 = ~n5945 | ~n3181;
  assign n5817 = ~n3568 | ~n3567;
  assign n3570 = ~n3569;
  assign n3571 = ~n3570 & ~IR_REG_16__SCAN_IN;
  assign n3572 = ~n3571 & ~n3755;
  assign n6411 = IR_REG_17__SCAN_IN ^ n3572;
  assign n3575 = ~n6411 | ~n3469;
  assign n3573 = ~DATAI_17_;
  assign n3574 = n3469 | n3573;
  assign n3579 = ~n4573 | ~REG0_REG_18__SCAN_IN;
  assign n3577 = ~REG2_REG_18__SCAN_IN;
  assign n3578 = n4575 | n3577;
  assign n3581 = ~n3579 | ~n3578;
  assign n3580 = n3633 & REG1_REG_18__SCAN_IN;
  assign n3584 = ~n3581 & ~n3580;
  assign n5868 = n5861 ^ n3582;
  assign n3583 = ~n5868 | ~n3181;
  assign n3585 = ~DATAI_18_;
  assign n3592 = n3469 | n3585;
  assign n3587 = ~n3586;
  assign n3589 = n3588 | n3587;
  assign n3590 = ~n3589 | ~IR_REG_31__SCAN_IN;
  assign n6520 = ~n3590 ^ IR_REG_18__SCAN_IN;
  assign n3591 = ~n3469 | ~n6520;
  assign n5810 = ~REG3_REG_19__SCAN_IN ^ n3593;
  assign n3594 = ~n5810;
  assign n3601 = ~n3594 | ~n3180;
  assign n3596 = ~n4573 | ~REG0_REG_19__SCAN_IN;
  assign n3595 = ~n3633 | ~REG1_REG_19__SCAN_IN;
  assign n3599 = ~n3596 | ~n3595;
  assign n3597 = ~REG2_REG_19__SCAN_IN;
  assign n3598 = ~n4575 & ~n3597;
  assign n3600 = ~n3599 & ~n3598;
  assign n5865 = ~n3601 | ~n3600;
  assign n3603 = ~n3682 | ~IR_REG_31__SCAN_IN;
  assign n6572 = ~n3603 ^ n3602;
  assign n3605 = ~n3469 | ~n6211;
  assign n3604 = ~n3666 | ~DATAI_19_;
  assign n5981 = REG3_REG_23__SCAN_IN ^ n3606;
  assign n3613 = ~n5981 | ~n3180;
  assign n3608 = ~n4573 | ~REG0_REG_23__SCAN_IN;
  assign n3607 = ~n3633 | ~REG1_REG_23__SCAN_IN;
  assign n3611 = ~n3608 | ~n3607;
  assign n3609 = ~REG2_REG_23__SCAN_IN;
  assign n3610 = ~n4575 & ~n3609;
  assign n3612 = ~n3611 & ~n3610;
  assign n6260 = ~n3613 | ~n3612;
  assign n3614 = ~DATAI_23_;
  assign n4426 = n4189 ^ n3615;
  assign n3622 = ~n4426 | ~n3181;
  assign n3617 = ~n4573 | ~REG0_REG_22__SCAN_IN;
  assign n3616 = ~n3633 | ~REG1_REG_22__SCAN_IN;
  assign n3620 = ~n3617 | ~n3616;
  assign n3618 = ~REG2_REG_22__SCAN_IN;
  assign n3619 = ~n4575 & ~n3618;
  assign n3621 = ~n3620 & ~n3619;
  assign n4449 = ~n3666 | ~DATAI_22_;
  assign n6360 = REG3_REG_21__SCAN_IN ^ n3623;
  assign n3630 = ~n6360 | ~n3181;
  assign n3625 = ~n4573 | ~REG0_REG_21__SCAN_IN;
  assign n3624 = ~n3633 | ~REG1_REG_21__SCAN_IN;
  assign n3628 = ~n3625 | ~n3624;
  assign n3626 = ~REG2_REG_21__SCAN_IN;
  assign n3627 = ~n4575 & ~n3626;
  assign n3629 = ~n3628 & ~n3627;
  assign n6246 = ~n3630 | ~n3629;
  assign n3631 = ~DATAI_21_;
  assign n6251 = n6243 ^ n3632;
  assign n3641 = ~n6251 | ~n3181;
  assign n3635 = ~n3633 | ~REG1_REG_20__SCAN_IN;
  assign n3634 = ~n3460 | ~REG2_REG_20__SCAN_IN;
  assign n3639 = ~n3635 | ~n3634;
  assign n3636 = ~REG0_REG_20__SCAN_IN;
  assign n3638 = ~n3637 & ~n3636;
  assign n3640 = ~n3639 & ~n3638;
  assign n5780 = ~n3666 | ~DATAI_20_;
  assign n4346 = REG3_REG_27__SCAN_IN ^ n3658;
  assign n3665 = ~n4346 | ~n3180;
  assign n3660 = ~n4573 | ~REG0_REG_27__SCAN_IN;
  assign n3659 = ~n3633 | ~REG1_REG_27__SCAN_IN;
  assign n3663 = ~n3660 | ~n3659;
  assign n3661 = ~REG2_REG_27__SCAN_IN;
  assign n3662 = ~n4575 & ~n3661;
  assign n3664 = ~n3663 & ~n3662;
  assign n4347 = ~n3666 | ~DATAI_27_;
  assign n4278 = ~n3669 | ~REG3_REG_28__SCAN_IN;
  assign n3670 = ~n4278;
  assign n3677 = ~n3670 | ~n3180;
  assign n3672 = ~n4573 | ~REG0_REG_29__SCAN_IN;
  assign n3671 = ~n3633 | ~REG1_REG_29__SCAN_IN;
  assign n3675 = ~n3672 | ~n3671;
  assign n3673 = ~REG2_REG_29__SCAN_IN;
  assign n3674 = ~n4575 & ~n3673;
  assign n3676 = ~n3675 & ~n3674;
  assign n6556 = ~n3677 | ~n3676;
  assign n6204 = ~n6168;
  assign n3695 = ~n6204 & ~n6208;
  assign n3690 = ~n3692 | ~IR_REG_31__SCAN_IN;
  assign n3691 = IR_REG_31__SCAN_IN & IR_REG_22__SCAN_IN;
  assign n3693 = n3692 & n3691;
  assign n3694 = ~n6572 & ~n3852;
  assign n4703 = ~n4675;
  assign n4546 = ~n4552;
  assign n6106 = ~n6208;
  assign n3712 = ~n3709 | ~IR_REG_31__SCAN_IN;
  assign n3710 = ~n3712 | ~n3255;
  assign n3711 = ~n3710 | ~IR_REG_31__SCAN_IN;
  assign n3714 = ~n4511;
  assign n3713 = ~n4504;
  assign n3715 = ~n3714 | ~n3713;
  assign n3717 = ~n3715 | ~B_REG_SCAN_IN;
  assign n3716 = n4504 | B_REG_SCAN_IN;
  assign n3721 = ~n3717 | ~n3716;
  assign n3723 = ~D_REG_0__SCAN_IN & ~n4506;
  assign n3725 = ~D_REG_1__SCAN_IN & ~n4506;
  assign n3724 = ~n4501 & ~n4511;
  assign n3731 = ~D_REG_31__SCAN_IN & ~D_REG_29__SCAN_IN;
  assign n4540 = ~D_REG_26__SCAN_IN;
  assign n4539 = ~D_REG_30__SCAN_IN;
  assign n3729 = ~n4540 | ~n4539;
  assign n3727 = ~D_REG_13__SCAN_IN & ~D_REG_12__SCAN_IN;
  assign n3726 = ~D_REG_11__SCAN_IN & ~D_REG_10__SCAN_IN;
  assign n3728 = ~n3727 | ~n3726;
  assign n3730 = ~n3729 & ~n3728;
  assign n3747 = ~n3731 | ~n3730;
  assign n3733 = ~D_REG_19__SCAN_IN & ~D_REG_18__SCAN_IN;
  assign n3732 = ~D_REG_17__SCAN_IN & ~D_REG_16__SCAN_IN;
  assign n3737 = ~n3733 | ~n3732;
  assign n3735 = ~D_REG_21__SCAN_IN & ~D_REG_9__SCAN_IN;
  assign n3734 = ~D_REG_14__SCAN_IN & ~D_REG_20__SCAN_IN;
  assign n3736 = ~n3735 | ~n3734;
  assign n3745 = ~n3737 & ~n3736;
  assign n3739 = ~D_REG_6__SCAN_IN & ~D_REG_5__SCAN_IN;
  assign n3738 = ~D_REG_4__SCAN_IN & ~D_REG_23__SCAN_IN;
  assign n3743 = ~n3739 | ~n3738;
  assign n3741 = ~D_REG_15__SCAN_IN & ~D_REG_3__SCAN_IN;
  assign n3740 = ~D_REG_8__SCAN_IN & ~D_REG_7__SCAN_IN;
  assign n3742 = ~n3741 | ~n3740;
  assign n3744 = ~n3743 & ~n3742;
  assign n3746 = ~n3745 | ~n3744;
  assign n3752 = ~n3747 & ~n3746;
  assign n3749 = ~D_REG_25__SCAN_IN & ~D_REG_24__SCAN_IN;
  assign n3748 = ~D_REG_28__SCAN_IN & ~D_REG_27__SCAN_IN;
  assign n3750 = ~n3749 | ~n3748;
  assign n3751 = ~D_REG_2__SCAN_IN & ~n3750;
  assign n3753 = ~n3752 | ~n3751;
  assign n3754 = ~D_REG_22__SCAN_IN & ~n3753;
  assign n4151 = ~n4506 & ~n3754;
  assign n4272 = ~n4152;
  assign n3758 = ~n6553 & ~n4272;
  assign n4176 = ~n6216 & ~n3758;
  assign n4547 = ~n6208 | ~n6211;
  assign n4031 = ~n5666;
  assign n4080 = ~n5763;
  assign n6247 = ~n5780;
  assign n4120 = ~n6476;
  assign n4328 = ~n4347;
  assign n3875 = ~n6208 | ~n3852;
  assign n3853 = ~n6215 | ~n6572;
  assign n4553 = n4317 | n3853;
  assign U3149 = ~STATE_REG_SCAN_IN;
  assign n3873 = ~n6067 | ~n4369;
  assign n3874 = ~n3873 | ~n3872;
  assign n3876 = ~n3875;
  assign n3878 = ~n6067 | ~n3932;
  assign n3877 = ~n4142 | ~n4777;
  assign n3893 = ~n3878 | ~n3877;
  assign n4749 = ~n3894 ^ n3893;
  assign n3892 = ~n4749;
  assign n4142 = ~n3196;
  assign n3880 = ~n4765 | ~n4142;
  assign n4677 = ~REG1_REG_0__SCAN_IN;
  assign n3879 = n4175 | n4677;
  assign n3886 = ~n4324 & ~n5007;
  assign n4671 = n3887 | n3886;
  assign n3885 = ~n4765 | ~n3932;
  assign n3883 = ~n3196 & ~n5007;
  assign n3881 = ~IR_REG_0__SCAN_IN;
  assign n3882 = ~n4175 & ~n3881;
  assign n3884 = ~n3883 & ~n3882;
  assign n4672 = n3885 & n3884;
  assign n3890 = ~n4671 | ~n4672;
  assign n3889 = ~n3888 | ~n4367;
  assign n3891 = ~n4748;
  assign n3896 = ~n3892 | ~n3891;
  assign n3895 = n3894 | n3893;
  assign n4235 = ~n3896 | ~n3895;
  assign n3898 = ~n4876 | ~n4142;
  assign n3897 = n4240 | n4324;
  assign n3899 = ~n3898 | ~n3897;
  assign n3903 = ~n3899 ^ n4145;
  assign n3901 = ~n4876 | ~n3932;
  assign n3900 = ~n4142 | ~n5025;
  assign n3902 = n3901 & n3900;
  assign n3904 = ~n3903 | ~n3902;
  assign n4234 = ~n3905 | ~n3904;
  assign n3907 = ~n4928 | ~n4142;
  assign n3906 = n4902 | n4324;
  assign n3908 = ~n3907 | ~n3906;
  assign n3911 = ~n3908 ^ n4145;
  assign n3910 = ~n4928 | ~n4084;
  assign n3909 = ~n4142 | ~n4880;
  assign n3912 = ~n3910 | ~n3909;
  assign n4885 = ~n3911 ^ n3912;
  assign n3913 = ~n3911;
  assign n3914 = n3913 | n3912;
  assign n3926 = ~n4932;
  assign n3916 = ~n4879 | ~n4142;
  assign n3915 = n4925 | n4324;
  assign n3917 = ~n3916 | ~n3915;
  assign n3920 = ~n3917 ^ n4145;
  assign n3919 = ~n4879 | ~n4084;
  assign n3918 = ~n4142 | ~n4912;
  assign n3921 = n3919 & n3918;
  assign n3927 = n3920 | n3921;
  assign n3923 = ~n3920;
  assign n3922 = ~n3921;
  assign n3924 = n3923 | n3922;
  assign n4931 = ~n3927 | ~n3924;
  assign n3925 = ~n4931;
  assign n3928 = ~n3926 | ~n3925;
  assign n5081 = ~n3928 | ~n3927;
  assign n3930 = ~n6019 | ~n4142;
  assign n3929 = n6020 | n4324;
  assign n3931 = ~n3930 | ~n3929;
  assign n3936 = ~n3931 ^ n4145;
  assign n3935 = ~n6019 | ~n4084;
  assign n3934 = ~n4142 | ~n3933;
  assign n3937 = n3935 & n3934;
  assign n3941 = n3936 | n3937;
  assign n3939 = ~n3936;
  assign n3938 = ~n3937;
  assign n3940 = n3939 | n3938;
  assign n5080 = n3941 & n3940;
  assign n3942 = ~n5081 | ~n5080;
  assign n3949 = ~n3942 | ~n3941;
  assign n3944 = ~n5152 | ~n4142;
  assign n3943 = n5103 | n4324;
  assign n3945 = ~n3944 | ~n3943;
  assign n3948 = ~n3945 ^ n4367;
  assign n5095 = ~n3949 ^ n3948;
  assign n3947 = ~n5152 | ~n4084;
  assign n3946 = ~n4142 | ~n5045;
  assign n5094 = ~n3947 | ~n3946;
  assign n3950 = n3949 | n3948;
  assign n3953 = ~n5194 | ~n4142;
  assign n3952 = n5155 | n4324;
  assign n3954 = ~n3953 | ~n3952;
  assign n3957 = ~n3954 ^ n4145;
  assign n3956 = ~n5194 | ~n4084;
  assign n3955 = ~n4142 | ~n5119;
  assign n3958 = n3956 & n3955;
  assign n3962 = n3957 | n3958;
  assign n3960 = ~n3957;
  assign n3959 = ~n3958;
  assign n3961 = n3960 | n3959;
  assign n5146 = ~n3962 | ~n3961;
  assign n3964 = ~n5328 | ~n4142;
  assign n3963 = n5186 | n4324;
  assign n3965 = ~n3964 | ~n3963;
  assign n3968 = ~n3965 ^ n4145;
  assign n3967 = ~n5328 | ~n4084;
  assign n3966 = ~n4142 | ~n5277;
  assign n3969 = n3967 & n3966;
  assign n3973 = n3968 | n3969;
  assign n3971 = ~n3968;
  assign n3970 = ~n3969;
  assign n3972 = n3971 | n3970;
  assign n5274 = n3973 & n3972;
  assign n3974 = ~n5275 | ~n5274;
  assign n5332 = ~n3974 | ~n3973;
  assign n3976 = ~n5271 | ~n4142;
  assign n3975 = n5340 | n4324;
  assign n3977 = ~n3976 | ~n3975;
  assign n3980 = ~n3977 ^ n4145;
  assign n3979 = ~n5271 | ~n4084;
  assign n3978 = ~n4142 | ~n5237;
  assign n3981 = n3979 & n3978;
  assign n3985 = n3980 | n3981;
  assign n3983 = ~n3980;
  assign n3982 = ~n3981;
  assign n3984 = n3983 | n3982;
  assign n5331 = n3985 & n3984;
  assign n5335 = ~n5332 | ~n5331;
  assign n3987 = ~n5487 | ~n4142;
  assign n3986 = n5407 | n4324;
  assign n3988 = ~n3987 | ~n3986;
  assign n3992 = ~n3988 ^ n4367;
  assign n3990 = ~n5487 | ~n3932;
  assign n3989 = ~n4142 | ~n6024;
  assign n3991 = ~n3990 | ~n3989;
  assign n5404 = ~n3992 ^ n3991;
  assign n3993 = n3992 | n3991;
  assign n3995 = ~n5441 | ~n4142;
  assign n3994 = n5483 | n4324;
  assign n3996 = ~n3995 | ~n3994;
  assign n3999 = ~n3996 ^ n4145;
  assign n3998 = ~n5441 | ~n3932;
  assign n3997 = ~n4142 | ~n5361;
  assign n4000 = n3998 & n3997;
  assign n4002 = ~n3999;
  assign n4001 = ~n4000;
  assign n4003 = n4002 | n4001;
  assign n5491 = ~n4004 | ~n4003;
  assign n4007 = ~n5604 | ~n4142;
  assign n4006 = n5525 | n4324;
  assign n4008 = ~n4007 | ~n4006;
  assign n4011 = ~n4008 ^ n4367;
  assign n4010 = ~n5604 | ~n3932;
  assign n4009 = ~n4142 | ~n5446;
  assign n4012 = ~n4010 | ~n4009;
  assign n5533 = n4011 | n4012;
  assign n4015 = ~n5536 | ~n5533;
  assign n4014 = ~n4011;
  assign n4013 = ~n4012;
  assign n4018 = ~n5460 | ~n4142;
  assign n4017 = n4016 | n4324;
  assign n4019 = ~n4018 | ~n4017;
  assign n4027 = ~n4019 ^ n4145;
  assign n4021 = ~n5460 | ~n3932;
  assign n4020 = ~n4142 | ~n5594;
  assign n4028 = n4021 & n4020;
  assign n5597 = n4027 | n4028;
  assign n4023 = ~n5676 | ~n4142;
  assign n4022 = n5471 | n4324;
  assign n4024 = ~n4023 | ~n4022;
  assign n4036 = ~n4024 ^ n4145;
  assign n4026 = ~n5676 | ~n3932;
  assign n4025 = ~n4142 | ~n5465;
  assign n4037 = ~n4026 | ~n4025;
  assign n4403 = ~n4036 ^ n4037;
  assign n4030 = ~n4027;
  assign n4029 = ~n4028;
  assign n5598 = n4030 | n4029;
  assign n4044 = n4403 & n5598;
  assign n4033 = n5738 | n3196;
  assign n4032 = n4031 | n4324;
  assign n4034 = ~n4033 | ~n4032;
  assign n4043 = ~n4034 ^ n4367;
  assign n4035 = n4044 & n4043;
  assign n4039 = ~n4043;
  assign n4038 = ~n4036;
  assign n4041 = ~n4038 | ~n4037;
  assign n4040 = n4039 | n4041;
  assign n4042 = ~n4041;
  assign n4045 = ~n4043 & ~n4042;
  assign n4047 = n5738 | n4094;
  assign n4046 = ~n4369 | ~n5666;
  assign n5669 = ~n4047 | ~n4046;
  assign n5742 = ~n5673 | ~n3193;
  assign n4049 = ~n5943 | ~n4369;
  assign n4048 = n5744 | n4324;
  assign n4050 = ~n4049 | ~n4048;
  assign n4053 = ~n4050 ^ n4367;
  assign n4052 = ~n5943 | ~n4084;
  assign n4051 = ~n4369 | ~n5647;
  assign n4054 = ~n4052 | ~n4051;
  assign n4056 = ~n4053;
  assign n4055 = ~n4054;
  assign n4058 = ~n5817 | ~n4369;
  assign n4371 = ~n4324;
  assign n4057 = ~n4371 | ~n5701;
  assign n4059 = ~n4058 | ~n4057;
  assign n4062 = ~n4059 ^ n4145;
  assign n4061 = ~n5817 | ~n4084;
  assign n4060 = ~n4369 | ~n5701;
  assign n4063 = n4061 & n4060;
  assign n4065 = ~n4062;
  assign n4064 = ~n4063;
  assign n4066 = n4065 | n4064;
  assign n5947 = n4067 & n4066;
  assign n4069 = ~n5768 | ~n4369;
  assign n4068 = n5831 | n4324;
  assign n4070 = ~n4069 | ~n4068;
  assign n4073 = ~n4070 ^ n4145;
  assign n4072 = ~n5768 | ~n4084;
  assign n4071 = ~n4142 | ~n5864;
  assign n4074 = n4072 & n4071;
  assign n4076 = ~n4073;
  assign n4075 = ~n4074;
  assign n4077 = n4076 | n4075;
  assign n4079 = ~n5869 | ~n5870;
  assign n4419 = ~n4079 | ~n4078;
  assign n4082 = ~n5865 | ~n4142;
  assign n4081 = n4324 | n4080;
  assign n4083 = ~n4082 | ~n4081;
  assign n4088 = ~n4083 ^ n4367;
  assign n4086 = ~n5865 | ~n4084;
  assign n4085 = ~n4142 | ~n5763;
  assign n4087 = ~n4086 | ~n4085;
  assign n4420 = ~n4088 ^ n4087;
  assign n4092 = ~n6358 | ~n4369;
  assign n4091 = n4324 | n5780;
  assign n4093 = ~n4092 | ~n4091;
  assign n4130 = ~n4093 ^ n4367;
  assign n4096 = ~n6358 | ~n4084;
  assign n4095 = ~n4369 | ~n6247;
  assign n4129 = ~n4096 | ~n4095;
  assign n6347 = ~n4130 ^ n4129;
  assign n4098 = ~n6246 | ~n4369;
  assign n4097 = n6369 | n4324;
  assign n4099 = ~n4098 | ~n4097;
  assign n4126 = ~n4099 ^ n4145;
  assign n4101 = ~n6246 | ~n3932;
  assign n4100 = ~n4142 | ~n5924;
  assign n4127 = ~n4101 | ~n4100;
  assign n6350 = ~n4126 ^ n4127;
  assign n4131 = ~n6350;
  assign n6353 = n6347 | n4131;
  assign n4103 = ~n6365 | ~n4369;
  assign n4102 = n4324 | n4449;
  assign n4104 = ~n4103 | ~n4102;
  assign n4107 = ~n4104 ^ n4367;
  assign n4106 = ~n6365 | ~n3932;
  assign n4193 = ~n4449;
  assign n4105 = ~n4142 | ~n4193;
  assign n4108 = ~n4106 | ~n4105;
  assign n4133 = ~n4107 | ~n4108;
  assign n4110 = ~n4107;
  assign n4109 = ~n4108;
  assign n4111 = ~n4110 | ~n4109;
  assign n4196 = n6353 | n3237;
  assign n4113 = ~n6260 | ~n4369;
  assign n4112 = n4203 | n4324;
  assign n4114 = ~n4113 | ~n4112;
  assign n4135 = ~n4114 ^ n4145;
  assign n4116 = ~n6260 | ~n4084;
  assign n4115 = ~n4369 | ~n5963;
  assign n4136 = ~n4116 | ~n4115;
  assign n6459 = n4196 | n3201;
  assign n4118 = ~n6299 | ~n4369;
  assign n4117 = n6476 | n4324;
  assign n4119 = ~n4118 | ~n4117;
  assign n4123 = ~n4119 ^ n4145;
  assign n4122 = ~n6299 | ~n4084;
  assign n4121 = ~n4142 | ~n4120;
  assign n4124 = ~n4122 | ~n4121;
  assign n6463 = ~n4123 ^ n4124;
  assign n4140 = ~n6463;
  assign n4156 = n6459 | n4140;
  assign n4125 = ~n4123;
  assign n4141 = ~n4125 | ~n4124;
  assign n4128 = ~n4126;
  assign n4132 = n4128 & n4127;
  assign n6348 = ~n4130 | ~n4129;
  assign n6354 = ~n4131 & ~n6348;
  assign n4183 = ~n4132 & ~n6354;
  assign n4134 = n3237 | n4183;
  assign n4197 = n4134 & n4133;
  assign n4139 = n3201 | n4197;
  assign n4137 = ~n4135;
  assign n4138 = ~n4137 | ~n4136;
  assign n6461 = n4139 & n4138;
  assign n6467 = n4140 | n6461;
  assign n4158 = n4141 & n6467;
  assign n4144 = ~n6385 | ~n4142;
  assign n4143 = n6300 | n4324;
  assign n4146 = ~n4144 | ~n4143;
  assign n4247 = ~n4146 ^ n4145;
  assign n4148 = ~n6385 | ~n4084;
  assign n4147 = ~n4369 | ~n6288;
  assign n4248 = ~n4148 | ~n4147;
  assign n4155 = ~n4247 ^ n4248;
  assign n4150 = ~n4284 | ~n4282;
  assign n4174 = ~n4151 & ~n4150;
  assign n4170 = ~n4174 | ~n4505;
  assign n4172 = ~n4152 & ~n4169;
  assign n4153 = ~n6559 | ~n4172;
  assign n4159 = ~n4155;
  assign n4334 = n4156 | n4159;
  assign n4162 = ~n4553;
  assign n6219 = n4505 & n4162;
  assign n4165 = n4174 & n6219;
  assign n4166 = ~n4165;
  assign n6366 = ~n4166 & ~n4703;
  assign n4171 = n4170 | n6559;
  assign n4173 = ~n4172 & ~n6219;
  assign n4178 = ~n4174 & ~n4173;
  assign n4177 = ~n4176 | ~n4175;
  assign n6486 = ~n4237 & ~n4495;
  assign n4249 = ~n4247;
  assign n4338 = ~n4249 | ~n4248;
  assign n4252 = ~n6296 | ~n4369;
  assign n4251 = n4324 | n6375;
  assign n4253 = ~n4252 | ~n4251;
  assign n4257 = ~n4253 ^ n4367;
  assign n4255 = ~n6296 | ~n4084;
  assign n4254 = ~n4142 | ~n6388;
  assign n4256 = ~n4255 | ~n4254;
  assign n4342 = ~n4257 & ~n4256;
  assign n4336 = n4257 & n4256;
  assign n4379 = ~n6563;
  assign n4326 = ~n6563 | ~n4369;
  assign n4325 = n4324 | n4347;
  assign n4327 = ~n4326 | ~n4325;
  assign n4332 = ~n4327 ^ n4367;
  assign n4330 = ~n6563 | ~n4084;
  assign n4329 = ~n4142 | ~n4328;
  assign n4331 = ~n4330 | ~n4329;
  assign n4333 = ~n4332 & ~n4331;
  assign n4362 = n4332 & n4331;
  assign n4335 = ~n6460;
  assign n4344 = ~n4335 | ~n3197;
  assign n4337 = ~n4336;
  assign n4340 = n4338 & n4337;
  assign n4341 = n4340 & n4339;
  assign n4364 = ~n4361 | ~n4360;
  assign n4363 = ~n4362;
  assign n4377 = ~n4364 | ~n4363;
  assign n4366 = ~n5265 | ~n4084;
  assign n4365 = ~n4369 | ~n4370;
  assign n4368 = ~n4366 | ~n4365;
  assign n4375 = ~n4368 ^ n4367;
  assign n4373 = ~n5265 | ~n4369;
  assign n4372 = ~n4371 | ~n4370;
  assign n4374 = ~n4373 | ~n4372;
  assign n4376 = ~n4375 ^ n4374;
  assign n4378 = ~n4377 ^ n4376;
  assign n4389 = ~n4378 | ~n3178;
  assign n4381 = ~n6472 & ~n4379;
  assign n4380 = ~n6477 & ~n6568;
  assign n4383 = ~n4381 & ~n4380;
  assign n4382 = ~n6366 | ~n6556;
  assign n4387 = ~n4383 | ~n4382;
  assign n4385 = ~n6545 | ~n6486;
  assign n4384 = ~REG3_REG_28__SCAN_IN | ~U3149;
  assign n4386 = ~n4385 | ~n4384;
  assign n4388 = ~n4387 & ~n4386;
  assign U3217_Lock = ~n4389 | ~n4388;
  assign input_0 = keyinput_0 ^ DATAI_28_;
  assign input_1 = keyinput_1 ^ DATAI_27_;
  assign AND_1 = input_0 & input_1;
  assign input_2 = keyinput_2 ^ DATAI_26_;
  assign AND_2 = input_2 & AND_1;
  assign input_3 = ~keyinput_3 ^ DATAI_25_;
  assign AND_3 = input_3 & AND_2;
  assign input_4 = keyinput_4 ^ DATAI_24_;
  assign OR_4 = input_4 | AND_3;
  assign input_5 = keyinput_5 ^ DATAI_23_;
  assign AND_5 = input_5 & OR_4;
  assign input_6 = ~keyinput_6 ^ DATAI_22_;
  assign AND_6 = input_6 & AND_5;
  assign input_7 = keyinput_7 ^ DATAI_21_;
  assign OR_7 = input_7 | AND_6;
  assign input_8 = ~keyinput_8 ^ DATAI_20_;
  assign OR_8 = input_8 | OR_7;
  assign input_9 = keyinput_9 ^ DATAI_19_;
  assign OR_9 = input_9 | OR_8;
  assign input_10 = keyinput_10 ^ DATAI_18_;
  assign OR_10 = input_10 | OR_9;
  assign input_11 = ~keyinput_11 ^ DATAI_17_;
  assign AND_11 = input_11 & OR_10;
  assign input_12 = keyinput_12 ^ DATAI_16_;
  assign OR_12 = input_12 | AND_11;
  assign input_13 = ~keyinput_13 ^ DATAI_15_;
  assign OR_13 = input_13 | OR_12;
  assign input_14 = keyinput_14 ^ DATAI_14_;
  assign OR_14 = input_14 | OR_13;
  assign input_15 = keyinput_15 ^ DATAI_13_;
  assign AND_15 = input_15 & OR_14;
  assign input_16 = ~keyinput_16 ^ DATAI_12_;
  assign OR_16 = input_16 | AND_15;
  assign input_17 = ~keyinput_17 ^ DATAI_11_;
  assign AND_17 = input_17 & OR_16;
  assign input_18 = ~keyinput_18 ^ DATAI_10_;
  assign AND_18 = input_18 & AND_17;
  assign input_19 = keyinput_19 ^ DATAI_9_;
  assign AND_19 = input_19 & AND_18;
  assign input_20 = ~keyinput_20 ^ DATAI_8_;
  assign AND_20 = input_20 & AND_19;
  assign input_21 = ~keyinput_21 ^ DATAI_7_;
  assign AND_21 = input_21 & AND_20;
  assign input_22 = keyinput_22 ^ DATAI_6_;
  assign OR_22 = input_22 | AND_21;
  assign input_23 = ~keyinput_23 ^ DATAI_5_;
  assign OR_23 = input_23 | OR_22;
  assign input_24 = keyinput_24 ^ DATAI_4_;
  assign AND_24 = input_24 & OR_23;
  assign input_25 = keyinput_25 ^ DATAI_3_;
  assign OR_25 = input_25 | AND_24;
  assign input_26 = keyinput_26 ^ DATAI_2_;
  assign AND_26 = input_26 & OR_25;
  assign input_27 = keyinput_27 ^ DATAI_1_;
  assign AND_27 = input_27 & AND_26;
  assign input_28 = ~keyinput_28 ^ DATAI_0_;
  assign AND_28 = input_28 & AND_27;
  assign input_29 = ~keyinput_29 ^ STATE_REG_SCAN_IN;
  assign OR_29 = input_29 | AND_28;
  assign input_30 = keyinput_30 ^ REG3_REG_7__SCAN_IN;
  assign AND_30 = input_30 & OR_29;
  assign input_31 = keyinput_31 ^ REG3_REG_27__SCAN_IN;
  assign OR_31 = input_31 | AND_30;
  assign input_32 = keyinput_32 ^ REG3_REG_14__SCAN_IN;
  assign AND_32 = input_32 & OR_31;
  assign input_33 = ~keyinput_33 ^ REG3_REG_23__SCAN_IN;
  assign AND_33 = input_33 & AND_32;
  assign input_34 = ~keyinput_34 ^ REG3_REG_10__SCAN_IN;
  assign OR_34 = input_34 | AND_33;
  assign input_35 = ~keyinput_35 ^ REG3_REG_3__SCAN_IN;
  assign OR_35 = input_35 | OR_34;
  assign input_36 = ~keyinput_36 ^ REG3_REG_19__SCAN_IN;
  assign AND_36 = input_36 & OR_35;
  assign input_37 = keyinput_37 ^ REG3_REG_28__SCAN_IN;
  assign AND_37 = input_37 & AND_36;
  assign input_38 = ~keyinput_38 ^ REG3_REG_8__SCAN_IN;
  assign OR_38 = input_38 | AND_37;
  assign input_39 = keyinput_39 ^ REG3_REG_1__SCAN_IN;
  assign AND_39 = input_39 & OR_38;
  assign input_40 = ~keyinput_40 ^ REG3_REG_21__SCAN_IN;
  assign AND_40 = input_40 & AND_39;
  assign input_41 = ~keyinput_41 ^ REG3_REG_12__SCAN_IN;
  assign OR_41 = input_41 | AND_40;
  assign input_42 = ~keyinput_42 ^ REG3_REG_25__SCAN_IN;
  assign OR_42 = input_42 | OR_41;
  assign input_43 = ~keyinput_43 ^ REG3_REG_16__SCAN_IN;
  assign AND_43 = input_43 & OR_42;
  assign input_44 = keyinput_44 ^ REG3_REG_5__SCAN_IN;
  assign AND_44 = input_44 & AND_43;
  assign input_45 = keyinput_45 ^ REG3_REG_17__SCAN_IN;
  assign OR_45 = input_45 | AND_44;
  assign input_46 = ~keyinput_46 ^ REG3_REG_24__SCAN_IN;
  assign OR_46 = input_46 | OR_45;
  assign input_47 = keyinput_47 ^ REG3_REG_4__SCAN_IN;
  assign OR_47 = input_47 | OR_46;
  assign input_48 = ~keyinput_48 ^ REG3_REG_9__SCAN_IN;
  assign AND_48 = input_48 & OR_47;
  assign input_49 = ~keyinput_49 ^ REG3_REG_0__SCAN_IN;
  assign OR_49 = input_49 | AND_48;
  assign input_50 = ~keyinput_50 ^ REG3_REG_20__SCAN_IN;
  assign AND_50 = input_50 & OR_49;
  assign input_51 = ~keyinput_51 ^ REG3_REG_13__SCAN_IN;
  assign OR_51 = input_51 | AND_50;
  assign input_52 = ~keyinput_52 ^ IR_REG_0__SCAN_IN;
  assign OR_52 = input_52 | OR_51;
  assign input_53 = keyinput_53 ^ IR_REG_1__SCAN_IN;
  assign OR_53 = input_53 | OR_52;
  assign input_54 = keyinput_54 ^ IR_REG_2__SCAN_IN;
  assign OR_54 = input_54 | OR_53;
  assign input_55 = ~keyinput_55 ^ IR_REG_3__SCAN_IN;
  assign AND_55 = input_55 & OR_54;
  assign input_56 = ~keyinput_56 ^ IR_REG_4__SCAN_IN;
  assign OR_56 = input_56 | AND_55;
  assign input_57 = ~keyinput_57 ^ IR_REG_5__SCAN_IN;
  assign AND_57 = input_57 & OR_56;
  assign input_58 = ~keyinput_58 ^ IR_REG_6__SCAN_IN;
  assign AND_58 = input_58 & AND_57;
  assign input_59 = ~keyinput_59 ^ IR_REG_7__SCAN_IN;
  assign OR_59 = input_59 | AND_58;
  assign input_60 = keyinput_60 ^ IR_REG_8__SCAN_IN;
  assign OR_60 = input_60 | OR_59;
  assign input_61 = ~keyinput_61 ^ IR_REG_9__SCAN_IN;
  assign OR_61 = input_61 | OR_60;
  assign input_62 = keyinput_62 ^ IR_REG_10__SCAN_IN;
  assign AND_62 = input_62 & OR_61;
  assign input_63 = keyinput_63 ^ IR_REG_11__SCAN_IN;
  assign OR_63 = input_63 | AND_62;
  assign input_64 = ~keyinput_64 ^ IR_REG_12__SCAN_IN;
  assign OR_64 = input_64 | OR_63;
  assign input_65 = ~keyinput_65 ^ IR_REG_13__SCAN_IN;
  assign OR_65 = input_65 | OR_64;
  assign input_66 = ~keyinput_66 ^ IR_REG_14__SCAN_IN;
  assign OR_66 = input_66 | OR_65;
  assign input_67 = ~keyinput_67 ^ IR_REG_15__SCAN_IN;
  assign OR_67 = input_67 | OR_66;
  assign input_68 = keyinput_68 ^ IR_REG_16__SCAN_IN;
  assign OR_68 = input_68 | OR_67;
  assign input_69 = keyinput_69 ^ IR_REG_17__SCAN_IN;
  assign AND_69 = input_69 & OR_68;
  assign input_70 = keyinput_70 ^ IR_REG_18__SCAN_IN;
  assign OR_70 = input_70 | AND_69;
  assign input_71 = keyinput_71 ^ IR_REG_19__SCAN_IN;
  assign OR_71 = input_71 | OR_70;
  assign input_72 = keyinput_72 ^ IR_REG_20__SCAN_IN;
  assign AND_72 = input_72 & OR_71;
  assign input_73 = ~keyinput_73 ^ IR_REG_21__SCAN_IN;
  assign OR_73 = input_73 | AND_72;
  assign input_74 = ~keyinput_74 ^ IR_REG_22__SCAN_IN;
  assign OR_74 = input_74 | OR_73;
  assign input_75 = keyinput_75 ^ IR_REG_23__SCAN_IN;
  assign AND_75 = input_75 & OR_74;
  assign input_76 = ~keyinput_76 ^ IR_REG_24__SCAN_IN;
  assign OR_76 = input_76 | AND_75;
  assign input_77 = keyinput_77 ^ IR_REG_25__SCAN_IN;
  assign OR_77 = input_77 | OR_76;
  assign input_78 = keyinput_78 ^ IR_REG_26__SCAN_IN;
  assign OR_78 = input_78 | OR_77;
  assign input_79 = keyinput_79 ^ IR_REG_27__SCAN_IN;
  assign OR_79 = input_79 | OR_78;
  assign input_80 = keyinput_80 ^ DATAI_28_;
  assign input_81 = keyinput_81 ^ DATAI_27_;
  assign AND_81 = input_80 & input_81;
  assign input_82 = keyinput_82 ^ DATAI_26_;
  assign AND_82 = input_82 & AND_81;
  assign input_83 = keyinput_83 ^ DATAI_25_;
  assign AND_83 = input_83 & AND_82;
  assign input_84 = keyinput_84 ^ DATAI_24_;
  assign OR_84 = input_84 | AND_83;
  assign input_85 = ~keyinput_85 ^ DATAI_23_;
  assign AND_85 = input_85 & OR_84;
  assign input_86 = keyinput_86 ^ DATAI_22_;
  assign AND_86 = input_86 & AND_85;
  assign input_87 = ~keyinput_87 ^ DATAI_21_;
  assign OR_87 = input_87 | AND_86;
  assign input_88 = ~keyinput_88 ^ DATAI_20_;
  assign OR_88 = input_88 | OR_87;
  assign input_89 = ~keyinput_89 ^ DATAI_19_;
  assign OR_89 = input_89 | OR_88;
  assign input_90 = ~keyinput_90 ^ DATAI_18_;
  assign OR_90 = input_90 | OR_89;
  assign input_91 = keyinput_91 ^ DATAI_17_;
  assign AND_91 = input_91 & OR_90;
  assign input_92 = ~keyinput_92 ^ DATAI_16_;
  assign OR_92 = input_92 | AND_91;
  assign input_93 = keyinput_93 ^ DATAI_15_;
  assign OR_93 = input_93 | OR_92;
  assign input_94 = ~keyinput_94 ^ DATAI_14_;
  assign OR_94 = input_94 | OR_93;
  assign input_95 = keyinput_95 ^ DATAI_13_;
  assign AND_95 = input_95 & OR_94;
  assign input_96 = keyinput_96 ^ DATAI_12_;
  assign OR_96 = input_96 | AND_95;
  assign input_97 = ~keyinput_97 ^ DATAI_11_;
  assign AND_97 = input_97 & OR_96;
  assign input_98 = keyinput_98 ^ DATAI_10_;
  assign AND_98 = input_98 & AND_97;
  assign input_99 = keyinput_99 ^ DATAI_9_;
  assign AND_99 = input_99 & AND_98;
  assign input_100 = ~keyinput_100 ^ DATAI_8_;
  assign AND_100 = input_100 & AND_99;
  assign input_101 = ~keyinput_101 ^ DATAI_7_;
  assign AND_101 = input_101 & AND_100;
  assign input_102 = ~keyinput_102 ^ DATAI_6_;
  assign OR_102 = input_102 | AND_101;
  assign input_103 = ~keyinput_103 ^ DATAI_5_;
  assign OR_103 = input_103 | OR_102;
  assign input_104 = keyinput_104 ^ DATAI_4_;
  assign AND_104 = input_104 & OR_103;
  assign input_105 = keyinput_105 ^ DATAI_3_;
  assign OR_105 = input_105 | AND_104;
  assign input_106 = keyinput_106 ^ DATAI_2_;
  assign AND_106 = input_106 & OR_105;
  assign input_107 = ~keyinput_107 ^ DATAI_1_;
  assign AND_107 = input_107 & AND_106;
  assign input_108 = ~keyinput_108 ^ DATAI_0_;
  assign AND_108 = input_108 & AND_107;
  assign input_109 = ~keyinput_109 ^ STATE_REG_SCAN_IN;
  assign OR_109 = input_109 | AND_108;
  assign input_110 = ~keyinput_110 ^ REG3_REG_7__SCAN_IN;
  assign AND_110 = input_110 & OR_109;
  assign input_111 = keyinput_111 ^ REG3_REG_27__SCAN_IN;
  assign OR_111 = input_111 | AND_110;
  assign input_112 = keyinput_112 ^ REG3_REG_14__SCAN_IN;
  assign AND_112 = input_112 & OR_111;
  assign input_113 = keyinput_113 ^ REG3_REG_23__SCAN_IN;
  assign AND_113 = input_113 & AND_112;
  assign input_114 = ~keyinput_114 ^ REG3_REG_10__SCAN_IN;
  assign OR_114 = input_114 | AND_113;
  assign input_115 = keyinput_115 ^ REG3_REG_3__SCAN_IN;
  assign OR_115 = input_115 | OR_114;
  assign input_116 = keyinput_116 ^ REG3_REG_19__SCAN_IN;
  assign AND_116 = input_116 & OR_115;
  assign input_117 = ~keyinput_117 ^ REG3_REG_28__SCAN_IN;
  assign AND_117 = input_117 & AND_116;
  assign input_118 = keyinput_118 ^ REG3_REG_8__SCAN_IN;
  assign OR_118 = input_118 | AND_117;
  assign input_119 = ~keyinput_119 ^ REG3_REG_1__SCAN_IN;
  assign AND_119 = input_119 & OR_118;
  assign input_120 = keyinput_120 ^ REG3_REG_21__SCAN_IN;
  assign AND_120 = input_120 & AND_119;
  assign input_121 = keyinput_121 ^ REG3_REG_12__SCAN_IN;
  assign OR_121 = input_121 | AND_120;
  assign input_122 = ~keyinput_122 ^ REG3_REG_25__SCAN_IN;
  assign OR_122 = input_122 | OR_121;
  assign input_123 = ~keyinput_123 ^ REG3_REG_16__SCAN_IN;
  assign AND_123 = input_123 & OR_122;
  assign input_124 = ~keyinput_124 ^ REG3_REG_5__SCAN_IN;
  assign AND_124 = input_124 & AND_123;
  assign input_125 = keyinput_125 ^ REG3_REG_17__SCAN_IN;
  assign OR_125 = input_125 | AND_124;
  assign input_126 = keyinput_126 ^ REG3_REG_24__SCAN_IN;
  assign OR_126 = input_126 | OR_125;
  assign input_127 = keyinput_127 ^ REG3_REG_4__SCAN_IN;
  assign OR_127 = input_127 | OR_126;
  assign input_128 = ~keyinput_128 ^ REG3_REG_9__SCAN_IN;
  assign AND_128 = input_128 & OR_127;
  assign input_129 = keyinput_129 ^ REG3_REG_0__SCAN_IN;
  assign OR_129 = input_129 | AND_128;
  assign input_130 = ~keyinput_130 ^ REG3_REG_20__SCAN_IN;
  assign AND_130 = input_130 & OR_129;
  assign input_131 = keyinput_131 ^ REG3_REG_13__SCAN_IN;
  assign OR_131 = input_131 | AND_130;
  assign input_132 = ~keyinput_132 ^ IR_REG_0__SCAN_IN;
  assign OR_132 = input_132 | OR_131;
  assign input_133 = keyinput_133 ^ IR_REG_1__SCAN_IN;
  assign OR_133 = input_133 | OR_132;
  assign input_134 = ~keyinput_134 ^ IR_REG_2__SCAN_IN;
  assign OR_134 = input_134 | OR_133;
  assign input_135 = ~keyinput_135 ^ IR_REG_3__SCAN_IN;
  assign AND_135 = input_135 & OR_134;
  assign input_136 = ~keyinput_136 ^ IR_REG_4__SCAN_IN;
  assign OR_136 = input_136 | AND_135;
  assign input_137 = keyinput_137 ^ IR_REG_5__SCAN_IN;
  assign AND_137 = input_137 & OR_136;
  assign input_138 = keyinput_138 ^ IR_REG_6__SCAN_IN;
  assign AND_138 = input_138 & AND_137;
  assign input_139 = ~keyinput_139 ^ IR_REG_7__SCAN_IN;
  assign OR_139 = input_139 | AND_138;
  assign input_140 = keyinput_140 ^ IR_REG_8__SCAN_IN;
  assign OR_140 = input_140 | OR_139;
  assign input_141 = keyinput_141 ^ IR_REG_9__SCAN_IN;
  assign OR_141 = input_141 | OR_140;
  assign input_142 = ~keyinput_142 ^ IR_REG_10__SCAN_IN;
  assign AND_142 = input_142 & OR_141;
  assign input_143 = keyinput_143 ^ IR_REG_11__SCAN_IN;
  assign OR_143 = input_143 | AND_142;
  assign input_144 = ~keyinput_144 ^ IR_REG_12__SCAN_IN;
  assign OR_144 = input_144 | OR_143;
  assign input_145 = ~keyinput_145 ^ IR_REG_13__SCAN_IN;
  assign OR_145 = input_145 | OR_144;
  assign input_146 = ~keyinput_146 ^ IR_REG_14__SCAN_IN;
  assign OR_146 = input_146 | OR_145;
  assign input_147 = keyinput_147 ^ IR_REG_15__SCAN_IN;
  assign OR_147 = input_147 | OR_146;
  assign input_148 = keyinput_148 ^ IR_REG_16__SCAN_IN;
  assign OR_148 = input_148 | OR_147;
  assign input_149 = keyinput_149 ^ IR_REG_17__SCAN_IN;
  assign AND_149 = input_149 & OR_148;
  assign input_150 = ~keyinput_150 ^ IR_REG_18__SCAN_IN;
  assign OR_150 = input_150 | AND_149;
  assign input_151 = ~keyinput_151 ^ IR_REG_19__SCAN_IN;
  assign OR_151 = input_151 | OR_150;
  assign input_152 = ~keyinput_152 ^ IR_REG_20__SCAN_IN;
  assign AND_152 = input_152 & OR_151;
  assign input_153 = ~keyinput_153 ^ IR_REG_21__SCAN_IN;
  assign OR_153 = input_153 | AND_152;
  assign input_154 = ~keyinput_154 ^ IR_REG_22__SCAN_IN;
  assign OR_154 = input_154 | OR_153;
  assign input_155 = keyinput_155 ^ IR_REG_23__SCAN_IN;
  assign AND_155 = input_155 & OR_154;
  assign input_156 = keyinput_156 ^ IR_REG_24__SCAN_IN;
  assign OR_156 = input_156 | AND_155;
  assign input_157 = ~keyinput_157 ^ IR_REG_25__SCAN_IN;
  assign OR_157 = input_157 | OR_156;
  assign input_158 = ~keyinput_158 ^ IR_REG_26__SCAN_IN;
  assign OR_158 = input_158 | OR_157;
  assign input_159 = keyinput_159 ^ IR_REG_27__SCAN_IN;
  assign OR_159 = input_159 | OR_158;
  assign OR_159_INV = ~OR_159;
  assign CASOP = OR_79 & OR_159_INV;
  assign U3217 = U3217_Lock ^ CASOP;
endmodule


