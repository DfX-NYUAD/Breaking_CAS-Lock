// Benchmark "c3540" written by ABC on Thu Mar  5 01:06:55 2020

module c3540 ( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire G432, G442, G447, G456, G460, G463, G467, G476, G479, G483, G492,
    G501, G504, G513, G517, G526, G530, G540, G587, G704, G707, G714, G717,
    G724, G731, G732, G736, G741, G758, G776, G780, G788, G791, G798, G799,
    G802, G826, G828, G831, G833, G836, G839, G842, G845, G848, G851, G890,
    G898, G907, G1032, G1035, G1048, G1049, G1050, G1051, G1540, G1699,
    G1826, G1827, G1828, G2051, G2478, G2865, G2868, G2931, G2934, G2939,
    G2942, G2947, G2950, G2957, G2960, G3007, G3079, G3087, G3095, G3103,
    G3419, G588, G759, G1541, G1772, G1829, G1834, G2052, G625, G545, G546,
    G547, G548, G549, G550, G551, G552, G2937, G2938, G2945, G2946, G621,
    G626, G635, G636, G3085, G3101, G657, G675, G721, G784, G794, G807,
    G816, G823, G860, G861, G864, G893, G896, G897, G3093, G905, G906,
    G3109, G973, G980, G987, G994, G1001, G1008, G1015, G1022, G1038,
    G1043, G1054, G1057, G1512, G1681, G1717, G1724, G1731, G1738, G1745,
    G1752, G1759, G1766, G1773, G1790, G1808, G2278, G2481, G3425, G2871,
    G2874, G2953, G2954, G2963, G2964, G3010, G3013, G3017, G3020, G3027,
    G3030, G3037, G3040, G3082, G3090, G3098, G3106, G352, G553, G554,
    G555, G556, G560, G561, G650, G956, G974, G975, G976, G981, G982, G988,
    G989, G990, G995, G996, G997, G1002, G1003, G1004, G1009, G1010, G1016,
    G1017, G1018, G1023, G1024, G1025, G1720, G1727, G1734, G1741, G1748,
    G1755, G1762, G1769, G1791, G1809, G1851, G1901, G1952, G2002, G2057,
    G2109, G2162, G2214, G2955, G2956, G2965, G2966, G354, G557, G562,
    G586, G630, G634, G639, G642, G3086, G644, G646, G3102, G654, G660,
    G678, G804, G806, G855, G867, G903, G3094, G912, G3110, G915, G927,
    G941, G977, G978, G984, G985, G991, G992, G998, G999, G1005, G1006,
    G1012, G1013, G1019, G1020, G1026, G1027, G1060, G1063, G1066, G1069,
    G1527, G1530, G1542, G1563, G1572, G1581, G1585, G1589, G1593, G1597,
    G1601, G1605, G1716, G1718, G1723, G1725, G1730, G1732, G1737, G1739,
    G1744, G1746, G1751, G1753, G1758, G1760, G1765, G1767, G1852, G1856,
    G1870, G1902, G1906, G1920, G1953, G1957, G1971, G2003, G2007, G2021,
    G2058, G2062, G2076, G2110, G2114, G2128, G2163, G2167, G2181, G2215,
    G2219, G2233, G2285, G2288, G2289, G2293, G2298, G2302, G2877, G2983,
    G2986, G3014, G3015, G3023, G3024, G3033, G3034, G3043, G3044, G643,
    G647, G680, G904, G913, G920, G979, G993, G1000, G1007, G1021, G1028,
    G1719, G1721, G1726, G1728, G1733, G1735, G1740, G1742, G1747, G1749,
    G1754, G1756, G1761, G1763, G1768, G1770, G1794, G1799, G1812, G1817,
    G1859, G1909, G1960, G2010, G2065, G2117, G2170, G2222, G2678, G2697,
    G2716, G2733, G2751, G2768, G2785, G2802, G3016, G3025, G3026, G3035,
    G3036, G3045, G3046, G2989, G2990, G610, G613, G616, G640, G648, G655,
    G665, G668, G671, G683, G685, G688, G694, G696, G699, G870, G887, G901,
    G910, G914, G916, G942, G943, G1072, G1084, G1096, G1108, G1120, G1132,
    G1144, G1156, G1533, G1534, G1535, G1545, G1554, G1610, G1619, G1628,
    G1637, G1646, G1655, G1664, G1673, G1722, G1729, G1736, G1743, G1750,
    G1757, G1764, G1771, G1853, G1954, G2004, G2059, G2164, G2216, G2485,
    G2900, G2903, G2967, G2970, G2975, G2978, G3047, G3050, G3055, G3058,
    G574, G575, G617, G641, G649, G662, G672, G690, G691, G701, G702, G902,
    G911, G917, G923, G1538, G1871, G1872, G1873, G1921, G1922, G1923,
    G1972, G1973, G1974, G2022, G2023, G2024, G2077, G2078, G2079, G2129,
    G2130, G2131, G2182, G2183, G2184, G2234, G2235, G2236, G2973, G2974,
    G2981, G2982, G576, G3053, G3054, G3061, G3062, G645, G926, G928, G947,
    G983, G1011, G1075, G1087, G1099, G1111, G1123, G1135, G1147, G1159,
    G1168, G1177, G1186, G1195, G1204, G1213, G1222, G1231, G1609, G1611,
    G1618, G1620, G1627, G1629, G1636, G1638, G1645, G1647, G1654, G1656,
    G1663, G1665, G1672, G1674, G1862, G1866, G1874, G1924, G1963, G1967,
    G1975, G2013, G2017, G2025, G2068, G2072, G2080, G2132, G2173, G2177,
    G2185, G2225, G2229, G2237, G2488, G2679, G2680, G2698, G2699, G2717,
    G2718, G2734, G2735, G2752, G2753, G2769, G2770, G2786, G2787, G2803,
    G2804, G359, G1029, G565, G566, G569, G570, G589, G590, G595, G596,
    G929, G938, G944, G986, G1014, G1616, G1625, G1634, G1643, G360, G567,
    G571, G579, G591, G597, G614, G1240, G1241, G1242, G1243, G1244, G1245,
    G1246, G1247, G1257, G1258, G1259, G1260, G1261, G1262, G1263, G1264,
    G1274, G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1291, G1292,
    G1293, G1294, G1295, G1296, G1297, G1298, G1308, G1309, G1310, G1311,
    G1312, G1313, G1314, G1315, G1325, G1326, G1327, G1328, G1329, G1330,
    G1331, G1332, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349,
    G1359, G1360, G1361, G1362, G1363, G1364, G1365, G1366, G1376, G1377,
    G1378, G1379, G1380, G1381, G1382, G1383, G1393, G1394, G1395, G1396,
    G1397, G1398, G1399, G1400, G1410, G1411, G1412, G1413, G1414, G1415,
    G1416, G1417, G1427, G1428, G1429, G1430, G1431, G1432, G1433, G1434,
    G1444, G1445, G1446, G1447, G1448, G1449, G1450, G1451, G1461, G1462,
    G1463, G1464, G1465, G1466, G1467, G1468, G1478, G1479, G1480, G1481,
    G1482, G1483, G1484, G1485, G1495, G1496, G1497, G1498, G1499, G1500,
    G1501, G1502, G1877, G1880, G1891, G1903, G1927, G1930, G1978, G1981,
    G1992, G2028, G2031, G2042, G2085, G2088, G2099, G2111, G2137, G2140,
    G2190, G2193, G2204, G2242, G2245, G2256, G2320, G2341, G2354, G2367,
    G2383, G2391, G2474, G2475, G2476, G2477, G2482, G568, G618, G1248,
    G1249, G1250, G1251, G1252, G1253, G1254, G1255, G1265, G1266, G1267,
    G1268, G1269, G1270, G1271, G1272, G1282, G1283, G1284, G1285, G1286,
    G1287, G1288, G1289, G1299, G1300, G1301, G1302, G1303, G1304, G1305,
    G1306, G1316, G1317, G1318, G1319, G1320, G1321, G1322, G1323, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1350, G1351, G1352,
    G1353, G1354, G1355, G1356, G1357, G1367, G1368, G1369, G1370, G1371,
    G1372, G1373, G1374, G1384, G1385, G1386, G1387, G1388, G1389, G1390,
    G1391, G1401, G1402, G1403, G1404, G1405, G1406, G1407, G1408, G1418,
    G1419, G1420, G1421, G1422, G1423, G1424, G1425, G1435, G1436, G1437,
    G1438, G1439, G1440, G1441, G1442, G1452, G1453, G1454, G1455, G1456,
    G1457, G1458, G1459, G1469, G1470, G1471, G1472, G1473, G1474, G1475,
    G1476, G1486, G1487, G1488, G1489, G1490, G1491, G1492, G1493, G1503,
    G1504, G1505, G1506, G1507, G1508, G1509, G1510, G2483, G600, G661,
    G669, G679, G1256, G1273, G1290, G1307, G1324, G1341, G1358, G1375,
    G1392, G1409, G1426, G1443, G1460, G1477, G1494, G1511, G1652, G1883,
    G1886, G1889, G1890, G1912, G1916, G1984, G1987, G1990, G1991, G2034,
    G2037, G2040, G2041, G2091, G2094, G2097, G2098, G2120, G2124, G2196,
    G2199, G2202, G2203, G2248, G2251, G2254, G2255, G2484, G2991, G2994,
    G2999, G3002, G3063, G3071, G3124, G3134, G3158, G3166, G3174, G3182,
    G3190, G3200, G3224, G3232, G3240, G3248, G663, G673, G681, G1536,
    G1537, G1582, G1583, G1586, G1587, G1590, G1591, G1594, G1595, G1598,
    G1599, G1602, G1603, G1606, G1607, G1894, G1997, G2047, G2102, G2209,
    G2261, G2489, G3005, G3006, G3077, G3069, G2997, G2998, G689, G700,
    G1539, G1584, G1588, G1592, G1596, G1600, G1604, G1608, G1661, G1892,
    G1893, G1933, G1936, G1939, G1940, G1941, G1993, G1996, G2043, G2046,
    G2100, G2101, G2143, G2146, G2149, G2150, G2151, G2205, G2208, G2257,
    G2260, G3138, G2328, G3162, G3170, G3178, G3186, G3204, G2375, G3236,
    G3244, G3252, G3228, G3066, G3074, G3128, G3194, G619, G620, G582,
    G583, G692, G703, G1612, G1621, G1630, G1639, G1648, G1657, G1666,
    G1675, G1895, G1946, G1998, G2048, G2103, G2156, G2210, G2262, G2271,
    G2311, G356, G357, G603, G3078, G606, G3070, G1670, G1679, G1942,
    G1945, G2152, G2155, G2445, G2448, G2455, G2458, G3142, G3150, G3208,
    G3216, G604, G607, G1947, G2157, G2317, G2338, G2351, G2364, G2380,
    G2388, G605, G608, G2272, G2312, G3146, G3154, G3220, G3212, G2444,
    G2451, G2454, G2461, G2530, G3323, G349, G350, G2265, G2273, G2274,
    G2309, G2313, G2314, G2325, G2372, G2523, G2533, G3121, G3131, G3155,
    G3163, G3171, G3179, G3187, G3197, G3221, G3229, G3237, G3245, G2275,
    G2315, G3329, G2324, G2350, G2363, G2371, G2387, G2400, G2268, G3137,
    G3161, G2345, G3169, G3177, G2358, G3185, G3203, G3235, G3243, G2395,
    G3251, G3227, G2432, G2490, G3127, G3130, G3139, G3147, G3193, G3196,
    G3205, G3213, G2307, G2308, G2323, G2349, G2362, G2370, G2386, G2399,
    G2344, G2357, G2394, G2431, G2464, G2491, G3129, G3195, G368, G1615,
    G2337, G1633, G1642, G1651, G2379, G1669, G1678, G3145, G2332, G3153,
    G2346, G2359, G3219, G2396, G3211, G2425, G2433, G3272, G3308, G1613,
    G2336, G1631, G1640, G1649, G2378, G1667, G1676, G2331, G2424, G2467,
    G2495, G3295, G3374, G1614, G1624, G1632, G1641, G1650, G1660, G1668,
    G1677, G2333, G2406, G2409, G2415, G2419, G2426, G2439, G2518, G3276,
    G3312, G2612, G3326, G1617, G1622, G1635, G1644, G1653, G1658, G1671,
    G1680, G2500, G2505, G2519, G3378, G2642, G2645, G3301, G1623, G1659,
    G2401, G2501, G2511, G2512, G2513, G2514, G2517, G2531, G2532, G2534,
    G2535, G2607, G3330, G2643, G2687, G2725, G2742, G2760, G2794, G2811,
    G3280, G3290, G3298, G3316, G3406, G3414, G3422, G1626, G1662, G2567,
    G2589, G2608, G2654, G3253, G3277, G3287, G3305, G3313, G3350, G932,
    G2508, G2524, G2525, G2526, G3294, G2609, G3410, G3418, G2624, G3426,
    G2629, G2647, G2706, G2777, G3264, G3284, G3302, G3303, G3320, G3398,
    G2657, G398, G933, G2527, G3259, G3354, G3293, G2563, G3311, G2585,
    G2625, G3283, G3286, G3304, G3319, G3322, G3358, G3366, G3382, G3390,
    G397, G2544, G2562, G2584, G3402, G2626, G2632, G2634, G2650, G3268,
    G3256, G3285, G3321, G3371, G3403, G3411, G362, G1030, G2564, G3362,
    G3370, G2586, G3386, G3394, G2633, G3261, G3269, G3347, G3395, G363,
    G2536, G3260, G3377, G2580, G3409, G2616, G3417, G2622, G2635, G2805,
    G2808, G3334, G3342, G3454, G2537, G3275, G2540, G3353, G2557, G2579,
    G3401, G2602, G2615, G2621, G3267, G3112, G3355, G3363, G3379, G3387,
    G2538, G2539, G3338, G3346, G2556, G2581, G2601, G2617, G2623, G2638,
    G3458, G2814, G2816, G3111, G2541, G2558, G3361, G2571, G3369, G2577,
    G3385, G2593, G3393, G2598, G2603, G3113, G3116, G3451, G395, G2570,
    G2576, G2592, G2597, G2736, G2739, G2788, G3438, G3446, G3459, G3119,
    G3120, G2572, G2578, G2594, G2599, G2677, G3457, G2700, G2771, G3331,
    G3339, G3427, G3443, G954, G955, G2600, G3442, G3450, G2676, G2745,
    G2748, G3465, G3435, G950, G3337, G2548, G3345, G2553, G2661, G2662,
    G3433, G3449, G2672, G2674, G2719, G2754, G3430, G383, G951, G2547,
    G2552, G2663, G2670, G3441, G2671, G2675, G3491, G3499, G2549, G2554,
    G2664, G3434, G2669, G2673, G2757, G2791, G365, G1031, G2555, G2665,
    G2667, G2774, G3497, G3505, G366, G2658, G2659, G2666, G2668, G2681,
    G2763, G2765, G2797, G2799, G2660, G2703, G2722, G2780, G2782, G386,
    G392, G2684, G3462, G3470, G389, G2709, G2713, G2728, G2730, G2922,
    G3467, G2690, G2694, G2821, G3466, G3474, G380, G2822, G3473, G2827,
    G2839, G2883, G3507, G2823, G2826, G2880, G2925, G2928, G3510, G2828,
    G3494, G3502, G3513, G3544, G3552, G406, G2929, G3475, G3483, G3514,
    G3515, G3541, G3549, G2930, G2842, G3498, G2852, G3506, G3548, G3556,
    G3478, G3486, G3516, G408, G3481, G3489, G2843, G2853, G3547, G2887,
    G2896, G3555, G3520, G2831, G3482, G2836, G3490, G2844, G2848, G2886,
    G2895, G2832, G2837, G2849, G3524, G2888, G2891, G2833, G2838, G2892,
    G3517, G2906, G2908, G2913, G3523, G2855, G2907, G2909, G3525, G3533,
    G2854, G2910, G3560, G3568, G2856, G3539, G3531, G3572, G3564, G3557,
    G3565, G3528, G3536, G2921, G2917, G3571, G3563, G2863, G2859, G2920,
    G2916, G3540, G3532, G2864, G2860, G403, G404, G400, G401;
  assign G432 = G50;
  assign G442 = ~G50;
  assign G447 = G58;
  assign G456 = ~G58;
  assign G460 = G68;
  assign G463 = ~G68;
  assign G467 = G68;
  assign G476 = G77;
  assign G479 = ~G77;
  assign G483 = G77;
  assign G492 = G87;
  assign G501 = ~G87;
  assign G504 = G97;
  assign G513 = ~G97;
  assign G517 = G107;
  assign G526 = ~G107;
  assign G530 = G116;
  assign G540 = ~G116;
  assign G587 = G257 | G264;
  assign G704 = ~G1;
  assign G707 = G1;
  assign G714 = ~G1;
  assign G717 = G13;
  assign G724 = ~G13;
  assign G731 = G13 & G20;
  assign G732 = ~G20;
  assign G736 = G20;
  assign G741 = ~G20;
  assign G758 = ~G33;
  assign G776 = G33;
  assign G780 = ~G33;
  assign G788 = G33 & G41;
  assign G791 = ~G41;
  assign G798 = G41 | G45;
  assign G799 = G45;
  assign G802 = ~G45;
  assign G826 = ~G50;
  assign G828 = G58;
  assign G831 = ~G58;
  assign G833 = G68;
  assign G836 = ~G68;
  assign G839 = G87;
  assign G842 = ~G87;
  assign G845 = G97;
  assign G848 = ~G97;
  assign G851 = ~G107;
  assign G890 = G1;
  assign G898 = G68;
  assign G907 = G107;
  assign G1032 = ~G20;
  assign G1035 = G190;
  assign G1048 = ~G200;
  assign G1049 = G20 & G200;
  assign G1050 = ~G20 | ~G200;
  assign G1051 = G20 & G179;
  assign G1540 = ~G20;
  assign G1699 = G1698 | G33;
  assign G1826 = ~G1 | ~G13;
  assign G1827 = ~G33 | ~G1 | ~G20;
  assign G1828 = ~G20;
  assign G2051 = ~G33;
  assign G2478 = G179;
  assign G2865 = ~G213;
  assign G2868 = G343;
  assign G2931 = G226;
  assign G2934 = G232;
  assign G2939 = G238;
  assign G2942 = G244;
  assign G2947 = G250;
  assign G2950 = G257;
  assign G2957 = G264;
  assign G2960 = G270;
  assign G3007 = G50;
  assign G3079 = G58;
  assign G3087 = G58;
  assign G3095 = G97;
  assign G3103 = G97;
  assign G3419 = G330;
  assign G588 = G250 & G587;
  assign G759 = G758 | G20;
  assign G1541 = G1540 | G169;
  assign G1772 = ~G731;
  assign G1829 = G1828 | G1;
  assign G1834 = G1826 & G1827;
  assign G2052 = G2051 | G1;
  assign G625 = G836 & G826 & G831;
  assign G545 = ~G226 | ~G432;
  assign G546 = ~G232 | ~G447;
  assign G547 = ~G238 | ~G467;
  assign G548 = ~G244 | ~G483;
  assign G549 = ~G250 | ~G492;
  assign G550 = ~G257 | ~G504;
  assign G551 = ~G264 | ~G517;
  assign G552 = ~G270 | ~G530;
  assign G2937 = ~G2931;
  assign G2938 = ~G2934;
  assign G2945 = ~G2939;
  assign G2946 = ~G2942;
  assign G621 = ~G456 | ~G463;
  assign G626 = ~G513 | ~G526;
  assign G635 = ~G460 | ~G476;
  assign G636 = G442;
  assign G3085 = ~G3079;
  assign G3101 = ~G3095;
  assign G657 = G802;
  assign G675 = G802;
  assign G721 = G717;
  assign G784 = G780;
  assign G794 = G791;
  assign G807 = G714 & G798;
  assign G816 = G791 & G714 & G799;
  assign G823 = G704 & G799;
  assign G860 = G736 & G707 & G724;
  assign G861 = ~G736 | ~G707 | ~G724;
  assign G864 = ~G707 | ~G724;
  assign G893 = G890;
  assign G896 = ~G45 | ~G717 | ~G732;
  assign G897 = ~G836 | ~G826 | ~G831;
  assign G3093 = ~G3087;
  assign G905 = G851 & G842 & G848;
  assign G906 = ~G851 | ~G842 | ~G848;
  assign G3109 = ~G3103;
  assign G973 = ~G741;
  assign G980 = ~G741;
  assign G987 = ~G741;
  assign G994 = ~G741;
  assign G1001 = ~G741;
  assign G1008 = ~G741;
  assign G1015 = ~G741;
  assign G1022 = ~G741;
  assign G1038 = G1032 | G1035;
  assign G1043 = ~G1032 & ~G1035;
  assign G1054 = G1051;
  assign G1057 = ~G1051;
  assign G1512 = G776;
  assign G1681 = G780;
  assign G1717 = ~G1699;
  assign G1724 = ~G1699;
  assign G1731 = ~G1699;
  assign G1738 = ~G1699;
  assign G1745 = ~G1699;
  assign G1752 = ~G1699;
  assign G1759 = ~G1699;
  assign G1766 = ~G1699;
  assign G1773 = G1 | G1772;
  assign G1790 = ~G788;
  assign G1808 = ~G788;
  assign G2278 = G732 & G704 & G717;
  assign G2481 = ~G2478;
  assign G3425 = ~G3419;
  assign G2871 = G2865 | G2868;
  assign G2874 = ~G2865 & ~G2868;
  assign G2953 = ~G2947;
  assign G2954 = ~G2950;
  assign G2963 = ~G2957;
  assign G2964 = ~G2960;
  assign G3010 = G456;
  assign G3013 = ~G3007;
  assign G3017 = G463;
  assign G3020 = G479;
  assign G3027 = G501;
  assign G3030 = G513;
  assign G3037 = G526;
  assign G3040 = G540;
  assign G3082 = G898;
  assign G3090 = G898;
  assign G3098 = G907;
  assign G3106 = G907;
  assign G352 = ~G479 | ~G625;
  assign G553 = G548 & G547 & G545 & G546;
  assign G554 = G552 & G551 & G549 & G550;
  assign G555 = ~G2934 | ~G2937;
  assign G556 = ~G2931 | ~G2938;
  assign G560 = ~G2942 | ~G2945;
  assign G561 = ~G2939 | ~G2946;
  assign G650 = G432 & G621;
  assign G956 = G890 & G896;
  assign G974 = ~G759;
  assign G975 = G741 & G759;
  assign G976 = G897 & G973;
  assign G981 = ~G759;
  assign G982 = G741 & G759;
  assign G988 = ~G759;
  assign G989 = G741 & G759;
  assign G990 = G836 & G987;
  assign G995 = ~G759;
  assign G996 = G741 & G759;
  assign G997 = G77 & G994;
  assign G1002 = ~G759;
  assign G1003 = G741 & G759;
  assign G1004 = G906 & G1001;
  assign G1009 = ~G759;
  assign G1010 = G741 & G759;
  assign G1016 = ~G759;
  assign G1017 = G741 & G759;
  assign G1018 = G851 & G1015;
  assign G1023 = ~G759;
  assign G1024 = G741 & G759;
  assign G1025 = G116 & G1022;
  assign G1720 = G222 & G1717;
  assign G1727 = G223 & G1724;
  assign G1734 = G226 & G1731;
  assign G1741 = G232 & G1738;
  assign G1748 = G238 & G1745;
  assign G1755 = G244 & G1752;
  assign G1762 = G250 & G1759;
  assign G1769 = G257 & G1766;
  assign G1791 = G1790 & G1 & G13;
  assign G1809 = G1808 & G1 & G13;
  assign G1851 = ~G1834;
  assign G1901 = ~G1834;
  assign G1952 = ~G1834;
  assign G2002 = ~G1834;
  assign G2057 = ~G1834;
  assign G2109 = ~G1834;
  assign G2162 = ~G1834;
  assign G2214 = ~G1834;
  assign G2955 = ~G2950 | ~G2953;
  assign G2956 = ~G2947 | ~G2954;
  assign G2965 = ~G2960 | ~G2963;
  assign G2966 = ~G2957 | ~G2964;
  assign G353 = ~G352;
  assign G354 = G87 & G626;
  assign G557 = ~G555 | ~G556;
  assign G562 = ~G560 | ~G561;
  assign G586 = ~G553 | ~G554;
  assign G630 = G540 & G905;
  assign G634 = ~G540 | ~G905;
  assign G639 = ~G636;
  assign G642 = ~G3082 | ~G3085;
  assign G3086 = ~G3082;
  assign G644 = G460 & G636;
  assign G646 = ~G3098 | ~G3101;
  assign G3102 = ~G3098;
  assign G654 = ~G87 | ~G626;
  assign G660 = ~G657;
  assign G678 = ~G675;
  assign G804 = ~G860 | ~G776;
  assign G806 = ~G860 | ~G780;
  assign G855 = ~G736 | ~G707 | ~G721;
  assign G867 = ~G794 | ~G736 | ~G707 | ~G724;
  assign G903 = ~G3090 | ~G3093;
  assign G3094 = ~G3090;
  assign G912 = ~G3106 | ~G3109;
  assign G3110 = ~G3106;
  assign G915 = ~G861;
  assign G927 = ~G893;
  assign G941 = ~G864;
  assign G977 = G828 & G974;
  assign G978 = G150 & G975;
  assign G984 = G833 & G981;
  assign G985 = G159 & G982;
  assign G991 = G77 & G988;
  assign G992 = G50 & G989;
  assign G998 = G839 & G995;
  assign G999 = G828 & G996;
  assign G1005 = G845 & G1002;
  assign G1006 = G833 & G1003;
  assign G1012 = G107 & G1009;
  assign G1013 = G77 & G1010;
  assign G1019 = G116 & G1016;
  assign G1020 = G839 & G1017;
  assign G1026 = G283 & G1023;
  assign G1027 = G845 & G1024;
  assign G1060 = G200 & G1054;
  assign G1063 = G1048 & G1054;
  assign G1066 = G1049 & G1057;
  assign G1069 = G1050 & G1057;
  assign G1527 = ~G784 | ~G794;
  assign G1530 = ~G776 | ~G794;
  assign G1542 = ~G1541 | ~G707 | ~G721;
  assign G1563 = ~G784 | ~G724 | ~G732;
  assign G1572 = ~G724 | ~G784;
  assign G1581 = ~G1512;
  assign G1585 = ~G1512;
  assign G1589 = ~G1512;
  assign G1593 = ~G1512;
  assign G1597 = ~G1512;
  assign G1601 = ~G1512;
  assign G1605 = ~G1512;
  assign G1716 = ~G1681;
  assign G1718 = G1681 & G1699;
  assign G1723 = ~G1681;
  assign G1725 = G1681 & G1699;
  assign G1730 = ~G1681;
  assign G1732 = G1681 & G1699;
  assign G1737 = ~G1681;
  assign G1739 = G1681 & G1699;
  assign G1744 = ~G1681;
  assign G1746 = G1681 & G1699;
  assign G1751 = ~G1681;
  assign G1753 = G1681 & G1699;
  assign G1758 = ~G1681;
  assign G1760 = G1681 & G1699;
  assign G1765 = ~G1681;
  assign G1767 = G1681 & G1699;
  assign G1852 = G1834 & G1773;
  assign G1856 = ~G50 & ~G1773;
  assign G1870 = ~G807;
  assign G1902 = G1834 & G1773;
  assign G1906 = ~G58 & ~G1773;
  assign G1920 = ~G807;
  assign G1953 = G1834 & G1773;
  assign G1957 = ~G68 & ~G1773;
  assign G1971 = ~G807;
  assign G2003 = G1834 & G1773;
  assign G2007 = ~G77 & ~G1773;
  assign G2021 = ~G807;
  assign G2058 = G1834 & G1773;
  assign G2062 = ~G87 & ~G1773;
  assign G2076 = ~G823;
  assign G2110 = G1834 & G1773;
  assign G2114 = ~G97 & ~G1773;
  assign G2128 = ~G816;
  assign G2163 = G1834 & G1773;
  assign G2167 = ~G107 & ~G1773;
  assign G2181 = ~G816;
  assign G2215 = G1834 & G1773;
  assign G2219 = ~G116 & ~G1773;
  assign G2233 = ~G816;
  assign G2285 = G2278 & G213;
  assign G2288 = ~G2278 | ~G213;
  assign G2289 = G343 & G2278 & G213;
  assign G2293 = ~G343 | ~G2278 | ~G213;
  assign G2298 = G343 & G2278 & G213;
  assign G2302 = ~G343 | ~G2278 | ~G213;
  assign G2877 = G2874;
  assign G2983 = ~G2955 | ~G2956;
  assign G2986 = ~G2965 | ~G2966;
  assign G3014 = ~G3010;
  assign G3015 = ~G3010 | ~G3013;
  assign G3023 = ~G3017;
  assign G3024 = ~G3020;
  assign G3033 = ~G3027;
  assign G3034 = ~G3030;
  assign G3043 = ~G3037;
  assign G3044 = ~G3040;
  assign G355 = ~G354;
  assign G643 = ~G3079 | ~G3086;
  assign G647 = ~G3095 | ~G3102;
  assign G680 = G650 & G675;
  assign G904 = ~G3087 | ~G3094;
  assign G913 = ~G3103 | ~G3110;
  assign G920 = G588 & G915;
  assign G979 = G978 | G976 | G977;
  assign G993 = G992 | G990 | G991;
  assign G1000 = G999 | G997 | G998;
  assign G1007 = G1006 | G1004 | G1005;
  assign G1021 = G1020 | G1018 | G1019;
  assign G1028 = G1027 | G1025 | G1026;
  assign G1719 = G77 & G1716;
  assign G1721 = G223 & G1718;
  assign G1726 = G87 & G1723;
  assign G1728 = G226 & G1725;
  assign G1733 = G97 & G1730;
  assign G1735 = G232 & G1732;
  assign G1740 = G107 & G1737;
  assign G1742 = G238 & G1739;
  assign G1747 = G116 & G1744;
  assign G1749 = G244 & G1746;
  assign G1754 = G283 & G1751;
  assign G1756 = G250 & G1753;
  assign G1761 = G294 & G1758;
  assign G1763 = G257 & G1760;
  assign G1768 = G303 & G1765;
  assign G1770 = G264 & G1767;
  assign G1794 = G1791;
  assign G1799 = ~G1791;
  assign G1812 = G1809;
  assign G1817 = ~G1809;
  assign G1859 = G1852 & G50 & G1829;
  assign G1909 = G1902 & G58 & G1829;
  assign G1960 = G1953 & G68 & G1829;
  assign G2010 = G2003 & G77 & G1829;
  assign G2065 = G2058 & G87 & G2052;
  assign G2117 = G2110 & G97 & G2052;
  assign G2170 = G2163 & G107 & G2052;
  assign G2222 = G2215 & G116 & G2052;
  assign G2678 = ~G956;
  assign G2697 = ~G956;
  assign G2716 = ~G956;
  assign G2733 = ~G956;
  assign G2751 = ~G956;
  assign G2768 = ~G956;
  assign G2785 = ~G956;
  assign G2802 = ~G956;
  assign G3016 = ~G3007 | ~G3014;
  assign G3025 = ~G3020 | ~G3023;
  assign G3026 = ~G3017 | ~G3024;
  assign G3035 = ~G3030 | ~G3033;
  assign G3036 = ~G3027 | ~G3034;
  assign G3045 = ~G3040 | ~G3043;
  assign G3046 = ~G3037 | ~G3044;
  assign G2989 = ~G2983;
  assign G2990 = ~G2986;
  assign G610 = ~G804;
  assign G613 = G804 & G806;
  assign G616 = ~G806;
  assign G640 = ~G642 | ~G643;
  assign G648 = ~G646 | ~G647;
  assign G655 = G58 & G442 & G630 & G635;
  assign G665 = ~G804;
  assign G668 = G804 & G806;
  assign G671 = ~G806;
  assign G683 = ~G804;
  assign G685 = ~G806;
  assign G688 = G804 & G806;
  assign G694 = ~G804;
  assign G696 = ~G806;
  assign G699 = G804 & G806;
  assign G870 = G867;
  assign G887 = G867;
  assign G901 = ~G903 | ~G904;
  assign G910 = ~G912 | ~G913;
  assign G914 = ~G855;
  assign G916 = G855 & G861;
  assign G942 = ~G855;
  assign G943 = G864 & G855;
  assign G1072 = ~G1043 | ~G1069;
  assign G1084 = ~G1043 | ~G1066;
  assign G1096 = ~G1038 | ~G1069;
  assign G1108 = ~G1038 | ~G1066;
  assign G1120 = ~G1043 | ~G1063;
  assign G1132 = ~G1043 | ~G1060;
  assign G1144 = ~G1038 | ~G1063;
  assign G1156 = ~G1038 | ~G1060;
  assign G1533 = ~G1527;
  assign G1534 = ~G1530;
  assign G1535 = G1527 & G1530;
  assign G1545 = G1542;
  assign G1554 = G1542;
  assign G1610 = ~G1572;
  assign G1619 = ~G1572;
  assign G1628 = ~G1572;
  assign G1637 = ~G1572;
  assign G1646 = ~G1563;
  assign G1655 = ~G1563;
  assign G1664 = ~G1563;
  assign G1673 = ~G1563;
  assign G1722 = G1721 | G1719 | G1720;
  assign G1729 = G1728 | G1726 | G1727;
  assign G1736 = G1735 | G1733 | G1734;
  assign G1743 = G1742 | G1740 | G1741;
  assign G1750 = G1749 | G1747 | G1748;
  assign G1757 = G1756 | G1754 | G1755;
  assign G1764 = G1763 | G1761 | G1762;
  assign G1771 = G1770 | G1768 | G1769;
  assign G1853 = G979 & G1851;
  assign G1954 = G993 & G1952;
  assign G2004 = G1000 & G2002;
  assign G2059 = G1007 & G2057;
  assign G2164 = G1021 & G2162;
  assign G2216 = G1028 & G2214;
  assign G2485 = G2293;
  assign G2900 = G2877 & G2897;
  assign G2903 = ~G2877 | ~G2897;
  assign G2967 = G557;
  assign G2970 = G562;
  assign G2975 = G557;
  assign G2978 = G562;
  assign G3047 = ~G3015 | ~G3016;
  assign G3050 = ~G3025 | ~G3026;
  assign G3055 = ~G3035 | ~G3036;
  assign G3058 = ~G3045 | ~G3046;
  assign G574 = ~G2986 | ~G2989;
  assign G575 = ~G2983 | ~G2990;
  assign G617 = G501 & G613;
  assign G641 = G639 & G640 & G476;
  assign G649 = G530 & G648;
  assign G662 = G655 & G657;
  assign G672 = G513 & G668;
  assign G690 = G654 & G685;
  assign G691 = G540 & G688;
  assign G701 = G634 & G696;
  assign G702 = G526 & G699;
  assign G902 = ~G901;
  assign G911 = ~G910;
  assign G917 = G650 & G914;
  assign G923 = G586 & G916;
  assign G1538 = G442 & G1535;
  assign G1871 = G1870 & G1817 & G226;
  assign G1872 = G807 & G1817 & G274;
  assign G1873 = G1812 & G1722;
  assign G1921 = G1920 & G1817 & G232;
  assign G1922 = G807 & G1817 & G274;
  assign G1923 = G1812 & G1729;
  assign G1972 = G1971 & G1817 & G238;
  assign G1973 = G807 & G1817 & G274;
  assign G1974 = G1812 & G1736;
  assign G2022 = G2021 & G1817 & G244;
  assign G2023 = G807 & G1817 & G274;
  assign G2024 = G1812 & G1743;
  assign G2077 = G2076 & G1799 & G250;
  assign G2078 = G823 & G1799 & G274;
  assign G2079 = G1794 & G1750;
  assign G2129 = G2128 & G1799 & G257;
  assign G2130 = G816 & G1799 & G274;
  assign G2131 = G1794 & G1757;
  assign G2182 = G2181 & G1799 & G264;
  assign G2183 = G816 & G1799 & G274;
  assign G2184 = G1794 & G1764;
  assign G2234 = G2233 & G1799 & G270;
  assign G2235 = G816 & G1799 & G274;
  assign G2236 = G1794 & G1771;
  assign G2973 = ~G2967;
  assign G2974 = ~G2970;
  assign G2981 = ~G2975;
  assign G2982 = ~G2978;
  assign G576 = ~G574 | ~G575;
  assign G3053 = ~G3047;
  assign G3054 = ~G3050;
  assign G3061 = ~G3055;
  assign G3062 = ~G3058;
  assign G645 = G641 | G644;
  assign G926 = ~G887;
  assign G928 = G887 & G893;
  assign G947 = G649 & G942;
  assign G983 = G902 & G980;
  assign G1011 = G911 & G1008;
  assign G1075 = G1072;
  assign G1087 = G1084;
  assign G1099 = G1096;
  assign G1111 = G1108;
  assign G1123 = G1120;
  assign G1135 = G1132;
  assign G1147 = G1144;
  assign G1159 = G1156;
  assign G1168 = G1072;
  assign G1177 = G1084;
  assign G1186 = G1096;
  assign G1195 = G1108;
  assign G1204 = G1120;
  assign G1213 = G1132;
  assign G1222 = G1144;
  assign G1231 = G1156;
  assign G1609 = ~G1545;
  assign G1611 = G1545 & G1572;
  assign G1618 = ~G1545;
  assign G1620 = G1545 & G1572;
  assign G1627 = ~G1545;
  assign G1629 = G1545 & G1572;
  assign G1636 = ~G1545;
  assign G1638 = G1545 & G1572;
  assign G1645 = ~G1554;
  assign G1647 = G1554 & G1563;
  assign G1654 = ~G1554;
  assign G1656 = G1554 & G1563;
  assign G1663 = ~G1554;
  assign G1665 = G1554 & G1563;
  assign G1672 = ~G1554;
  assign G1674 = G1554 & G1563;
  assign G1862 = G1859 | G1853 | G1856;
  assign G1866 = ~G1859 & ~G1853 & ~G1856;
  assign G1874 = G1873 | G1871 | G1872;
  assign G1924 = G1923 | G1921 | G1922;
  assign G1963 = G1960 | G1954 | G1957;
  assign G1967 = ~G1960 & ~G1954 & ~G1957;
  assign G1975 = G1974 | G1972 | G1973;
  assign G2013 = G2010 | G2004 | G2007;
  assign G2017 = ~G2010 & ~G2004 & ~G2007;
  assign G2025 = G2024 | G2022 | G2023;
  assign G2068 = G2065 | G2059 | G2062;
  assign G2072 = ~G2065 & ~G2059 & ~G2062;
  assign G2080 = G2079 | G2077 | G2078;
  assign G2132 = G2131 | G2129 | G2130;
  assign G2173 = G2170 | G2164 | G2167;
  assign G2177 = ~G2170 & ~G2164 & ~G2167;
  assign G2185 = G2184 | G2182 | G2183;
  assign G2225 = G2222 | G2216 | G2219;
  assign G2229 = ~G2222 & ~G2216 & ~G2219;
  assign G2237 = G2236 | G2234 | G2235;
  assign G2488 = ~G2485;
  assign G2679 = ~G870;
  assign G2680 = G956 & G870;
  assign G2698 = ~G870;
  assign G2699 = G956 & G870;
  assign G2717 = ~G870;
  assign G2718 = G956 & G870;
  assign G2734 = ~G870;
  assign G2735 = G956 & G870;
  assign G2752 = ~G870;
  assign G2753 = G956 & G870;
  assign G2769 = ~G870;
  assign G2770 = G956 & G870;
  assign G2786 = ~G870;
  assign G2787 = G956 & G870;
  assign G2803 = ~G870;
  assign G2804 = G956 & G870;
  assign G359 = G923 | G917 | G920;
  assign G1029 = ~G923 & ~G917 & ~G920;
  assign G565 = ~G2970 | ~G2973;
  assign G566 = ~G2967 | ~G2974;
  assign G569 = ~G2978 | ~G2981;
  assign G570 = ~G2975 | ~G2982;
  assign G589 = ~G3050 | ~G3053;
  assign G590 = ~G3047 | ~G3054;
  assign G595 = ~G3058 | ~G3061;
  assign G596 = ~G3055 | ~G3062;
  assign G929 = G650 & G926;
  assign G938 = G630 & G928;
  assign G944 = G645 & G941;
  assign G986 = G985 | G983 | G984;
  assign G1014 = G1013 | G1011 | G1012;
  assign G1616 = G442 & G1611;
  assign G1625 = G456 & G1620;
  assign G1634 = G463 & G1629;
  assign G1643 = G479 & G1638;
  assign G360 = ~G1029;
  assign G567 = ~G565 | ~G566;
  assign G571 = ~G569 | ~G570;
  assign G579 = G576;
  assign G591 = ~G589 | ~G590;
  assign G597 = ~G595 | ~G596;
  assign G614 = G576 & G610;
  assign G1240 = ~G1075;
  assign G1241 = ~G1087;
  assign G1242 = ~G1099;
  assign G1243 = ~G1111;
  assign G1244 = ~G1123;
  assign G1245 = ~G1135;
  assign G1246 = ~G1147;
  assign G1247 = ~G1159;
  assign G1257 = ~G1075;
  assign G1258 = ~G1087;
  assign G1259 = ~G1099;
  assign G1260 = ~G1111;
  assign G1261 = ~G1123;
  assign G1262 = ~G1135;
  assign G1263 = ~G1147;
  assign G1264 = ~G1159;
  assign G1274 = ~G1075;
  assign G1275 = ~G1087;
  assign G1276 = ~G1099;
  assign G1277 = ~G1111;
  assign G1278 = ~G1123;
  assign G1279 = ~G1135;
  assign G1280 = ~G1147;
  assign G1281 = ~G1159;
  assign G1291 = ~G1075;
  assign G1292 = ~G1087;
  assign G1293 = ~G1099;
  assign G1294 = ~G1111;
  assign G1295 = ~G1123;
  assign G1296 = ~G1135;
  assign G1297 = ~G1147;
  assign G1298 = ~G1159;
  assign G1308 = ~G1075;
  assign G1309 = ~G1087;
  assign G1310 = ~G1099;
  assign G1311 = ~G1111;
  assign G1312 = ~G1123;
  assign G1313 = ~G1135;
  assign G1314 = ~G1147;
  assign G1315 = ~G1159;
  assign G1325 = ~G1075;
  assign G1326 = ~G1087;
  assign G1327 = ~G1099;
  assign G1328 = ~G1111;
  assign G1329 = ~G1123;
  assign G1330 = ~G1135;
  assign G1331 = ~G1147;
  assign G1332 = ~G1159;
  assign G1342 = ~G1075;
  assign G1343 = ~G1087;
  assign G1344 = ~G1099;
  assign G1345 = ~G1111;
  assign G1346 = ~G1123;
  assign G1347 = ~G1135;
  assign G1348 = ~G1147;
  assign G1349 = ~G1159;
  assign G1359 = ~G1075;
  assign G1360 = ~G1087;
  assign G1361 = ~G1099;
  assign G1362 = ~G1111;
  assign G1363 = ~G1123;
  assign G1364 = ~G1135;
  assign G1365 = ~G1147;
  assign G1366 = ~G1159;
  assign G1376 = ~G1168;
  assign G1377 = ~G1177;
  assign G1378 = ~G1186;
  assign G1379 = ~G1195;
  assign G1380 = ~G1204;
  assign G1381 = ~G1213;
  assign G1382 = ~G1222;
  assign G1383 = ~G1231;
  assign G1393 = ~G1168;
  assign G1394 = ~G1177;
  assign G1395 = ~G1186;
  assign G1396 = ~G1195;
  assign G1397 = ~G1204;
  assign G1398 = ~G1213;
  assign G1399 = ~G1222;
  assign G1400 = ~G1231;
  assign G1410 = ~G1168;
  assign G1411 = ~G1177;
  assign G1412 = ~G1186;
  assign G1413 = ~G1195;
  assign G1414 = ~G1204;
  assign G1415 = ~G1213;
  assign G1416 = ~G1222;
  assign G1417 = ~G1231;
  assign G1427 = ~G1168;
  assign G1428 = ~G1177;
  assign G1429 = ~G1186;
  assign G1430 = ~G1195;
  assign G1431 = ~G1204;
  assign G1432 = ~G1213;
  assign G1433 = ~G1222;
  assign G1434 = ~G1231;
  assign G1444 = ~G1168;
  assign G1445 = ~G1177;
  assign G1446 = ~G1186;
  assign G1447 = ~G1195;
  assign G1448 = ~G1204;
  assign G1449 = ~G1213;
  assign G1450 = ~G1222;
  assign G1451 = ~G1231;
  assign G1461 = ~G1168;
  assign G1462 = ~G1177;
  assign G1463 = ~G1186;
  assign G1464 = ~G1195;
  assign G1465 = ~G1204;
  assign G1466 = ~G1213;
  assign G1467 = ~G1222;
  assign G1468 = ~G1231;
  assign G1478 = ~G1168;
  assign G1479 = ~G1177;
  assign G1480 = ~G1186;
  assign G1481 = ~G1195;
  assign G1482 = ~G1204;
  assign G1483 = ~G1213;
  assign G1484 = ~G1222;
  assign G1485 = ~G1231;
  assign G1495 = ~G1168;
  assign G1496 = ~G1177;
  assign G1497 = ~G1186;
  assign G1498 = ~G1195;
  assign G1499 = ~G1204;
  assign G1500 = ~G1213;
  assign G1501 = ~G1222;
  assign G1502 = ~G1231;
  assign G1877 = G1874;
  assign G1880 = ~G1874;
  assign G1891 = ~G1866;
  assign G1903 = G986 & G1901;
  assign G1927 = G1924;
  assign G1930 = ~G1924;
  assign G1978 = G1975;
  assign G1981 = ~G1975;
  assign G1992 = ~G1967;
  assign G2028 = G2025;
  assign G2031 = ~G2025;
  assign G2042 = ~G2017;
  assign G2085 = G2080;
  assign G2088 = ~G2080;
  assign G2099 = ~G2072;
  assign G2111 = G1014 & G2109;
  assign G2137 = G2132;
  assign G2140 = ~G2132;
  assign G2190 = G2185;
  assign G2193 = ~G2185;
  assign G2204 = ~G2177;
  assign G2242 = G2237;
  assign G2245 = ~G2237;
  assign G2256 = ~G2229;
  assign G2320 = G2285 & G1862;
  assign G2341 = G2289 & G1963;
  assign G2354 = G2289 & G2013;
  assign G2367 = G2289 & G2068;
  assign G2383 = G2298 & G2173;
  assign G2391 = G2298 & G2225;
  assign G2474 = ~G2080;
  assign G2475 = ~G2132;
  assign G2476 = ~G2185;
  assign G2477 = ~G2237;
  assign G2482 = G2481 & G2237 & G2185 & G2080 & G2132;
  assign G361 = ~G359 | ~G360;
  assign G568 = ~G567;
  assign G618 = G617 | G614 | G616;
  assign G1248 = G124 & G1240;
  assign G1249 = G159 & G1241;
  assign G1250 = G150 & G1242;
  assign G1251 = G143 & G1243;
  assign G1252 = G137 & G1244;
  assign G1253 = G132 & G1245;
  assign G1254 = G128 & G1246;
  assign G1255 = G125 & G1247;
  assign G1265 = G125 & G1257;
  assign G1266 = G432 & G1258;
  assign G1267 = G159 & G1259;
  assign G1268 = G150 & G1260;
  assign G1269 = G143 & G1261;
  assign G1270 = G137 & G1262;
  assign G1271 = G132 & G1263;
  assign G1272 = G128 & G1264;
  assign G1282 = G128 & G1274;
  assign G1283 = G447 & G1275;
  assign G1284 = G432 & G1276;
  assign G1285 = G159 & G1277;
  assign G1286 = G150 & G1278;
  assign G1287 = G143 & G1279;
  assign G1288 = G137 & G1280;
  assign G1289 = G132 & G1281;
  assign G1299 = G132 & G1291;
  assign G1300 = G467 & G1292;
  assign G1301 = G447 & G1293;
  assign G1302 = G432 & G1294;
  assign G1303 = G159 & G1295;
  assign G1304 = G150 & G1296;
  assign G1305 = G143 & G1297;
  assign G1306 = G137 & G1298;
  assign G1316 = G137 & G1308;
  assign G1317 = G483 & G1309;
  assign G1318 = G467 & G1310;
  assign G1319 = G447 & G1311;
  assign G1320 = G432 & G1312;
  assign G1321 = G159 & G1313;
  assign G1322 = G150 & G1314;
  assign G1323 = G143 & G1315;
  assign G1333 = G143 & G1325;
  assign G1334 = G492 & G1326;
  assign G1335 = G483 & G1327;
  assign G1336 = G467 & G1328;
  assign G1337 = G447 & G1329;
  assign G1338 = G432 & G1330;
  assign G1339 = G159 & G1331;
  assign G1340 = G150 & G1332;
  assign G1350 = G150 & G1342;
  assign G1351 = G504 & G1343;
  assign G1352 = G492 & G1344;
  assign G1353 = G483 & G1345;
  assign G1354 = G467 & G1346;
  assign G1355 = G447 & G1347;
  assign G1356 = G432 & G1348;
  assign G1357 = G159 & G1349;
  assign G1367 = G159 & G1359;
  assign G1368 = G517 & G1360;
  assign G1369 = G504 & G1361;
  assign G1370 = G492 & G1362;
  assign G1371 = G483 & G1363;
  assign G1372 = G467 & G1364;
  assign G1373 = G447 & G1365;
  assign G1374 = G432 & G1366;
  assign G1384 = G283 & G1376;
  assign G1385 = G447 & G1377;
  assign G1386 = G467 & G1378;
  assign G1387 = G483 & G1379;
  assign G1388 = G492 & G1380;
  assign G1389 = G504 & G1381;
  assign G1390 = G517 & G1382;
  assign G1391 = G530 & G1383;
  assign G1401 = G294 & G1393;
  assign G1402 = G467 & G1394;
  assign G1403 = G483 & G1395;
  assign G1404 = G492 & G1396;
  assign G1405 = G504 & G1397;
  assign G1406 = G517 & G1398;
  assign G1407 = G530 & G1399;
  assign G1408 = G283 & G1400;
  assign G1418 = G303 & G1410;
  assign G1419 = G483 & G1411;
  assign G1420 = G492 & G1412;
  assign G1421 = G504 & G1413;
  assign G1422 = G517 & G1414;
  assign G1423 = G530 & G1415;
  assign G1424 = G283 & G1416;
  assign G1425 = G294 & G1417;
  assign G1435 = G311 & G1427;
  assign G1436 = G492 & G1428;
  assign G1437 = G504 & G1429;
  assign G1438 = G517 & G1430;
  assign G1439 = G530 & G1431;
  assign G1440 = G283 & G1432;
  assign G1441 = G294 & G1433;
  assign G1442 = G303 & G1434;
  assign G1452 = G317 & G1444;
  assign G1453 = G504 & G1445;
  assign G1454 = G517 & G1446;
  assign G1455 = G530 & G1447;
  assign G1456 = G283 & G1448;
  assign G1457 = G294 & G1449;
  assign G1458 = G303 & G1450;
  assign G1459 = G311 & G1451;
  assign G1469 = G322 & G1461;
  assign G1470 = G517 & G1462;
  assign G1471 = G530 & G1463;
  assign G1472 = G283 & G1464;
  assign G1473 = G294 & G1465;
  assign G1474 = G303 & G1466;
  assign G1475 = G311 & G1467;
  assign G1476 = G317 & G1468;
  assign G1486 = G326 & G1478;
  assign G1487 = G530 & G1479;
  assign G1488 = G283 & G1480;
  assign G1489 = G294 & G1481;
  assign G1490 = G303 & G1482;
  assign G1491 = G311 & G1483;
  assign G1492 = G317 & G1484;
  assign G1493 = G322 & G1485;
  assign G1503 = G329 & G1495;
  assign G1504 = G283 & G1496;
  assign G1505 = G294 & G1497;
  assign G1506 = G303 & G1498;
  assign G1507 = G311 & G1499;
  assign G1508 = G317 & G1500;
  assign G1509 = G322 & G1501;
  assign G1510 = G326 & G1502;
  assign G2483 = G2478 & G2477 & G2476 & G2474 & G2475;
  assign G600 = G597;
  assign G661 = G568 & G660;
  assign G669 = G597 & G665;
  assign G679 = G591 & G678;
  assign G1256 = ~G1255 & ~G1254 & ~G1253 & ~G1252 & ~G1251 & ~G1250 & ~G1248 & ~G1249;
  assign G1273 = ~G1272 & ~G1271 & ~G1270 & ~G1269 & ~G1268 & ~G1267 & ~G1265 & ~G1266;
  assign G1290 = ~G1289 & ~G1288 & ~G1287 & ~G1286 & ~G1285 & ~G1284 & ~G1282 & ~G1283;
  assign G1307 = ~G1306 & ~G1305 & ~G1304 & ~G1303 & ~G1302 & ~G1301 & ~G1299 & ~G1300;
  assign G1324 = ~G1323 & ~G1322 & ~G1321 & ~G1320 & ~G1319 & ~G1318 & ~G1316 & ~G1317;
  assign G1341 = ~G1340 & ~G1339 & ~G1338 & ~G1337 & ~G1336 & ~G1335 & ~G1333 & ~G1334;
  assign G1358 = ~G1357 & ~G1356 & ~G1355 & ~G1354 & ~G1353 & ~G1352 & ~G1350 & ~G1351;
  assign G1375 = ~G1374 & ~G1373 & ~G1372 & ~G1371 & ~G1370 & ~G1369 & ~G1367 & ~G1368;
  assign G1392 = ~G1391 & ~G1390 & ~G1389 & ~G1388 & ~G1387 & ~G1386 & ~G1384 & ~G1385;
  assign G1409 = ~G1408 & ~G1407 & ~G1406 & ~G1405 & ~G1404 & ~G1403 & ~G1401 & ~G1402;
  assign G1426 = ~G1425 & ~G1424 & ~G1423 & ~G1422 & ~G1421 & ~G1420 & ~G1418 & ~G1419;
  assign G1443 = ~G1442 & ~G1441 & ~G1440 & ~G1439 & ~G1438 & ~G1437 & ~G1435 & ~G1436;
  assign G1460 = ~G1459 & ~G1458 & ~G1457 & ~G1456 & ~G1455 & ~G1454 & ~G1452 & ~G1453;
  assign G1477 = ~G1476 & ~G1475 & ~G1474 & ~G1473 & ~G1472 & ~G1471 & ~G1469 & ~G1470;
  assign G1494 = ~G1493 & ~G1492 & ~G1491 & ~G1490 & ~G1489 & ~G1488 & ~G1486 & ~G1487;
  assign G1511 = ~G1510 & ~G1509 & ~G1508 & ~G1507 & ~G1506 & ~G1505 & ~G1503 & ~G1504;
  assign G1652 = G618 & G1647;
  assign G1883 = G1877 & G169 & G1862;
  assign G1886 = G1880 & G179 & G1862;
  assign G1889 = G1880 & G190 & G1866;
  assign G1890 = G1877 & G200 & G1866;
  assign G1912 = G1909 | G1903 | G1906;
  assign G1916 = ~G1909 & ~G1903 & ~G1906;
  assign G1984 = G1978 & G169 & G1963;
  assign G1987 = G1981 & G179 & G1963;
  assign G1990 = G1981 & G190 & G1967;
  assign G1991 = G1978 & G200 & G1967;
  assign G2034 = G2028 & G169 & G2013;
  assign G2037 = G2031 & G179 & G2013;
  assign G2040 = G2031 & G190 & G2017;
  assign G2041 = G2028 & G200 & G2017;
  assign G2091 = G2085 & G169 & G2068;
  assign G2094 = G2088 & G179 & G2068;
  assign G2097 = G2088 & G190 & G2072;
  assign G2098 = G2085 & G200 & G2072;
  assign G2120 = G2117 | G2111 | G2114;
  assign G2124 = ~G2117 & ~G2111 & ~G2114;
  assign G2196 = G2190 & G169 & G2173;
  assign G2199 = G2193 & G179 & G2173;
  assign G2202 = G2193 & G190 & G2177;
  assign G2203 = G2190 & G200 & G2177;
  assign G2248 = G2242 & G169 & G2225;
  assign G2251 = G2245 & G179 & G2225;
  assign G2254 = G2245 & G190 & G2229;
  assign G2255 = G2242 & G200 & G2229;
  assign G2484 = G2482 | G2483;
  assign G2991 = G571;
  assign G2994 = G579;
  assign G2999 = G571;
  assign G3002 = G579;
  assign G3063 = G591;
  assign G3071 = G591;
  assign G3124 = G2320;
  assign G3134 = G2320;
  assign G3158 = G2341;
  assign G3166 = G2341;
  assign G3174 = G2354;
  assign G3182 = G2354;
  assign G3190 = G2367;
  assign G3200 = G2367;
  assign G3224 = G2383;
  assign G3232 = G2383;
  assign G3240 = G2391;
  assign G3248 = G2391;
  assign G663 = ~G661 & ~G662;
  assign G673 = G672 | G669 | G671;
  assign G681 = ~G679 & ~G680;
  assign G1536 = G1256 & G1533;
  assign G1537 = G1392 & G1534;
  assign G1582 = G1273 & G1581;
  assign G1583 = G1409 & G1512;
  assign G1586 = G1290 & G1585;
  assign G1587 = G1426 & G1512;
  assign G1590 = G1307 & G1589;
  assign G1591 = G1443 & G1512;
  assign G1594 = G1324 & G1593;
  assign G1595 = G1460 & G1512;
  assign G1598 = G1341 & G1597;
  assign G1599 = G1477 & G1512;
  assign G1602 = G1358 & G1601;
  assign G1603 = G1494 & G1512;
  assign G1606 = G1375 & G1605;
  assign G1607 = G1511 & G1512;
  assign G1894 = G1891 | G1889 | G1890;
  assign G1997 = G1992 | G1990 | G1991;
  assign G2047 = G2042 | G2040 | G2041;
  assign G2102 = G2099 | G2097 | G2098;
  assign G2209 = G2204 | G2202 | G2203;
  assign G2261 = G2256 | G2254 | G2255;
  assign G2489 = G2484 & G2488;
  assign G3005 = ~G2999;
  assign G3006 = ~G3002;
  assign G3077 = ~G3071;
  assign G3069 = ~G3063;
  assign G2997 = ~G2991;
  assign G2998 = ~G2994;
  assign G689 = G681 & G683;
  assign G700 = G663 & G694;
  assign G1539 = G1538 | G1536 | G1537;
  assign G1584 = G1582 | G1583;
  assign G1588 = G1586 | G1587;
  assign G1592 = G1590 | G1591;
  assign G1596 = G1594 | G1595;
  assign G1600 = G1598 | G1599;
  assign G1604 = G1602 | G1603;
  assign G1608 = G1606 | G1607;
  assign G1661 = G673 & G1656;
  assign G1892 = G1883 | G1886;
  assign G1893 = ~G1883 & ~G1886;
  assign G1933 = G1927 & G169 & G1912;
  assign G1936 = G1930 & G179 & G1912;
  assign G1939 = G1930 & G190 & G1916;
  assign G1940 = G1927 & G200 & G1916;
  assign G1941 = ~G1916;
  assign G1993 = G1984 | G1987;
  assign G1996 = ~G1984 & ~G1987;
  assign G2043 = G2034 | G2037;
  assign G2046 = ~G2034 & ~G2037;
  assign G2100 = G2091 | G2094;
  assign G2101 = ~G2091 & ~G2094;
  assign G2143 = G2137 & G169 & G2120;
  assign G2146 = G2140 & G179 & G2120;
  assign G2149 = G2140 & G190 & G2124;
  assign G2150 = G2137 & G200 & G2124;
  assign G2151 = ~G2124;
  assign G2205 = G2196 | G2199;
  assign G2208 = ~G2196 & ~G2199;
  assign G2257 = G2248 | G2251;
  assign G2260 = ~G2248 & ~G2251;
  assign G3138 = ~G3134;
  assign G2328 = G2285 & G1912;
  assign G3162 = ~G3158;
  assign G3170 = ~G3166;
  assign G3178 = ~G3174;
  assign G3186 = ~G3182;
  assign G3204 = ~G3200;
  assign G2375 = G2298 & G2120;
  assign G3236 = ~G3232;
  assign G3244 = ~G3240;
  assign G3252 = ~G3248;
  assign G3228 = ~G3224;
  assign G3066 = G600;
  assign G3074 = G600;
  assign G3128 = ~G3124;
  assign G3194 = ~G3190;
  assign G619 = ~G2994 | ~G2997;
  assign G620 = ~G2991 | ~G2998;
  assign G582 = ~G3002 | ~G3005;
  assign G583 = ~G2999 | ~G3006;
  assign G692 = G691 | G689 | G690;
  assign G703 = G702 | G700 | G701;
  assign G1612 = G1539 & G1609;
  assign G1621 = G1584 & G1618;
  assign G1630 = G1588 & G1627;
  assign G1639 = G1592 & G1636;
  assign G1648 = G1596 & G1645;
  assign G1657 = G1600 & G1654;
  assign G1666 = G1604 & G1663;
  assign G1675 = G1608 & G1672;
  assign G1895 = G1893 & G1894;
  assign G1946 = G1941 | G1939 | G1940;
  assign G1998 = G1996 & G1997;
  assign G2048 = G2046 & G2047;
  assign G2103 = G2101 & G2102;
  assign G2156 = G2151 | G2149 | G2150;
  assign G2210 = G2208 & G2209;
  assign G2262 = G2260 & G2261;
  assign G2271 = ~G1892;
  assign G2311 = ~G2100;
  assign G356 = ~G619 | ~G620;
  assign G357 = ~G582 | ~G583;
  assign G603 = ~G3074 | ~G3077;
  assign G3078 = ~G3074;
  assign G606 = ~G3066 | ~G3069;
  assign G3070 = ~G3066;
  assign G1670 = G703 & G1665;
  assign G1679 = G692 & G1674;
  assign G1942 = G1933 | G1936;
  assign G1945 = ~G1933 & ~G1936;
  assign G2152 = G2143 | G2146;
  assign G2155 = ~G2143 & ~G2146;
  assign G2445 = G1993 & G2293;
  assign G2448 = G2043 & G2293;
  assign G2455 = G2205 & G2302;
  assign G2458 = G2257 & G2302;
  assign G3142 = G2328;
  assign G3150 = G2328;
  assign G3208 = G2375;
  assign G3216 = G2375;
  assign G358 = ~G356 | ~G357;
  assign G604 = ~G3071 | ~G3078;
  assign G607 = ~G3063 | ~G3070;
  assign G1947 = G1945 & G1946;
  assign G2157 = G2155 & G2156;
  assign G2317 = G1895;
  assign G2338 = G1998;
  assign G2351 = G2048;
  assign G2364 = G2103;
  assign G2380 = G2210;
  assign G2388 = G2262;
  assign G605 = ~G603 | ~G604;
  assign G608 = ~G606 | ~G607;
  assign G2272 = ~G1895 | ~G1942;
  assign G2312 = ~G2103 | ~G2152;
  assign G3146 = ~G3142;
  assign G3154 = ~G3150;
  assign G3220 = ~G3216;
  assign G3212 = ~G3208;
  assign G2444 = G1942 & G2288;
  assign G2451 = G2448;
  assign G2454 = G2152 & G2293;
  assign G2461 = G2458;
  assign G2530 = ~G2445;
  assign G3323 = G2458;
  assign G349 = ~G605;
  assign G350 = ~G608;
  assign G2265 = G2048 & G1998 & G1895 & G1947;
  assign G2273 = ~G1993 | ~G1895 | ~G1947;
  assign G2274 = ~G1895 | ~G1998 | ~G2043 | ~G1947;
  assign G2309 = G2262 & G2210 & G2103 & G2157;
  assign G2313 = ~G2205 | ~G2103 | ~G2157;
  assign G2314 = ~G2103 | ~G2210 | ~G2257 | ~G2157;
  assign G2325 = G1947;
  assign G2372 = G2157;
  assign G2523 = ~G2444;
  assign G2533 = ~G2454;
  assign G3121 = G2317;
  assign G3131 = G2317;
  assign G3155 = G2338;
  assign G3163 = G2338;
  assign G3171 = G2351;
  assign G3179 = G2351;
  assign G3187 = G2364;
  assign G3197 = G2364;
  assign G3221 = G2380;
  assign G3229 = G2380;
  assign G3237 = G2388;
  assign G3245 = G2388;
  assign G351 = ~G349 | ~G350;
  assign G2275 = ~G2274 | ~G2273 | ~G2271 | ~G2272;
  assign G2315 = ~G2314 | ~G2313 | ~G2311 | ~G2312;
  assign G3329 = ~G3323;
  assign G372 = G2309 & G2265;
  assign G2324 = ~G3131 | ~G3138;
  assign G2350 = ~G3163 | ~G3170;
  assign G2363 = ~G3179 | ~G3186;
  assign G2371 = ~G3197 | ~G3204;
  assign G2387 = ~G3229 | ~G3236;
  assign G2400 = ~G3245 | ~G3252;
  assign G2268 = G2265;
  assign G3137 = ~G3131;
  assign G3161 = ~G3155;
  assign G2345 = ~G3155 | ~G3162;
  assign G3169 = ~G3163;
  assign G3177 = ~G3171;
  assign G2358 = ~G3171 | ~G3178;
  assign G3185 = ~G3179;
  assign G3203 = ~G3197;
  assign G3235 = ~G3229;
  assign G3243 = ~G3237;
  assign G2395 = ~G3237 | ~G3244;
  assign G3251 = ~G3245;
  assign G3227 = ~G3221;
  assign G2432 = ~G3221 | ~G3228;
  assign G2490 = G2309 & G2485;
  assign G3127 = ~G3121;
  assign G3130 = ~G3121 | ~G3128;
  assign G3139 = G2325;
  assign G3147 = G2325;
  assign G3193 = ~G3187;
  assign G3196 = ~G3187 | ~G3194;
  assign G3205 = G2372;
  assign G3213 = G2372;
  assign G2307 = ~G2265 | ~G2315;
  assign G2308 = ~G2275;
  assign G2323 = ~G3134 | ~G3137;
  assign G2349 = ~G3166 | ~G3169;
  assign G2362 = ~G3182 | ~G3185;
  assign G2370 = ~G3200 | ~G3203;
  assign G2386 = ~G3232 | ~G3235;
  assign G2399 = ~G3248 | ~G3251;
  assign G2344 = ~G3158 | ~G3161;
  assign G2357 = ~G3174 | ~G3177;
  assign G2394 = ~G3240 | ~G3243;
  assign G2431 = ~G3224 | ~G3227;
  assign G2464 = G2315 & G2302;
  assign G2491 = G2489 | G2490;
  assign G3129 = ~G3124 | ~G3127;
  assign G3195 = ~G3190 | ~G3193;
  assign G368 = G2307 & G2308;
  assign G1615 = ~G2323 | ~G2324;
  assign G2337 = ~G3147 | ~G3154;
  assign G1633 = ~G2349 | ~G2350;
  assign G1642 = ~G2362 | ~G2363;
  assign G1651 = ~G2370 | ~G2371;
  assign G2379 = ~G3213 | ~G3220;
  assign G1669 = ~G2386 | ~G2387;
  assign G1678 = ~G2399 | ~G2400;
  assign G3145 = ~G3139;
  assign G2332 = ~G3139 | ~G3146;
  assign G3153 = ~G3147;
  assign G2346 = ~G2344 | ~G2345;
  assign G2359 = ~G2357 | ~G2358;
  assign G3219 = ~G3213;
  assign G2396 = ~G2394 | ~G2395;
  assign G3211 = ~G3205;
  assign G2425 = ~G3205 | ~G3212;
  assign G2433 = ~G2431 | ~G2432;
  assign G3272 = ~G3129 | ~G3130;
  assign G3308 = ~G3195 | ~G3196;
  assign G369 = ~G368;
  assign G1613 = ~G1615;
  assign G2336 = ~G3150 | ~G3153;
  assign G1631 = ~G1633;
  assign G1640 = ~G1642;
  assign G1649 = ~G1651;
  assign G2378 = ~G3216 | ~G3219;
  assign G1667 = ~G1669;
  assign G1676 = ~G1678;
  assign G2331 = ~G3142 | ~G3145;
  assign G2424 = ~G3208 | ~G3211;
  assign G2467 = G2464;
  assign G2495 = G2491;
  assign G3295 = G2464;
  assign G3374 = G330 & G2491;
  assign G1614 = G1613 & G1610;
  assign G1624 = ~G2336 | ~G2337;
  assign G1632 = G1631 & G1628;
  assign G1641 = G1640 & G1637;
  assign G1650 = G1649 & G1646;
  assign G1660 = ~G2378 | ~G2379;
  assign G1668 = G1667 & G1664;
  assign G1677 = G1676 & G1673;
  assign G2333 = ~G2331 | ~G2332;
  assign G2406 = G2346;
  assign G2409 = G2346;
  assign G2415 = G2359;
  assign G2419 = G2359;
  assign G2426 = ~G2424 | ~G2425;
  assign G2439 = G2396;
  assign G2518 = G2433 & G2461;
  assign G3276 = ~G3272;
  assign G3312 = ~G3308;
  assign G2612 = G330 & G2396;
  assign G3326 = G2433;
  assign G1617 = ~G1616 & ~G1612 & ~G1614;
  assign G1622 = ~G1624;
  assign G1635 = ~G1634 & ~G1630 & ~G1632;
  assign G1644 = ~G1643 & ~G1639 & ~G1641;
  assign G1653 = ~G1652 & ~G1648 & ~G1650;
  assign G1658 = ~G1660;
  assign G1671 = ~G1670 & ~G1666 & ~G1668;
  assign G1680 = ~G1679 & ~G1675 & ~G1677;
  assign G2500 = G2467 & G2268;
  assign G2505 = G2495 & G2268;
  assign G2519 = G2455 | G2518;
  assign G3378 = ~G3374;
  assign G2642 = ~G2467;
  assign G2645 = G2467;
  assign G3301 = ~G3295;
  assign G1623 = G1622 & G1619;
  assign G1659 = G1658 & G1655;
  assign G2401 = G2333;
  assign G2501 = G2275 | G2500;
  assign G2511 = G2409 & G2495 & G2419;
  assign G2512 = G2495 & G2415;
  assign G2513 = G2426 & G2439 & G2433;
  assign G2514 = G2439 & G2433;
  assign G2517 = G2467 & G2415;
  assign G2531 = ~G2409 | ~G2451;
  assign G2532 = ~G2467 | ~G2409 | ~G2419;
  assign G2534 = ~G2426 | ~G2455;
  assign G2535 = ~G2461 | ~G2426 | ~G2433;
  assign G2607 = ~G3326 | ~G3329;
  assign G3330 = ~G3326;
  assign G2643 = G2642 & G330 & G2491;
  assign G2687 = G1617 & G2680;
  assign G2725 = G1635 & G2718;
  assign G2742 = G1644 & G2735;
  assign G2760 = G1653 & G2753;
  assign G2794 = G1671 & G2787;
  assign G2811 = G1680 & G2804;
  assign G3280 = G2333;
  assign G3290 = G2409;
  assign G3298 = G2415;
  assign G3316 = G2426;
  assign G3406 = G2612;
  assign G3414 = G2612;
  assign G3422 = G2439 & G2439;
  assign G1626 = ~G1625 & ~G1621 & ~G1623;
  assign G1662 = ~G1661 & ~G1657 & ~G1659;
  assign G2567 = G330 & G2512;
  assign G2589 = G330 & G2513;
  assign G2608 = ~G3323 | ~G3330;
  assign G2654 = G2519;
  assign G3253 = G2505;
  assign G3277 = ~G2532 | ~G2530 | ~G2531;
  assign G3287 = G2448 | G2517;
  assign G3305 = ~G2535 | ~G2533 | ~G2534;
  assign G3313 = G2519;
  assign G3350 = G330 & G2511;
  assign G932 = G2643 | G2645;
  assign G2508 = G2419 & G2409 & G2495 & G2401;
  assign G2524 = ~G2401 | ~G2445;
  assign G2525 = ~G2451 | ~G2401 | ~G2406;
  assign G2526 = ~G2467 | ~G2419 | ~G2401 | ~G2406;
  assign G3294 = ~G3290;
  assign G2609 = ~G2607 | ~G2608;
  assign G3410 = ~G3406;
  assign G3418 = ~G3414;
  assign G2624 = ~G3422 | ~G3425;
  assign G3426 = ~G3422;
  assign G2629 = G2501;
  assign G2647 = ~G2643 & ~G2645;
  assign G2706 = G1626 & G2699;
  assign G2777 = G1662 & G2770;
  assign G3264 = G2501;
  assign G3284 = ~G3280;
  assign G3302 = ~G3298;
  assign G3303 = ~G3298 | ~G3301;
  assign G3320 = ~G3316;
  assign G3398 = G330 & G2514;
  assign G2657 = ~G2654;
  assign G398 = G2519 & G2654;
  assign G933 = G932 & G927;
  assign G2527 = ~G2526 | ~G2525 | ~G2523 | ~G2524;
  assign G3259 = ~G3253;
  assign G3354 = ~G3350;
  assign G3293 = ~G3287;
  assign G2563 = ~G3287 | ~G3294;
  assign G3311 = ~G3305;
  assign G2585 = ~G3305 | ~G3312;
  assign G2625 = ~G3419 | ~G3426;
  assign G3283 = ~G3277;
  assign G3286 = ~G3277 | ~G3284;
  assign G3304 = ~G3295 | ~G3302;
  assign G3319 = ~G3313;
  assign G3322 = ~G3313 | ~G3320;
  assign G3358 = G2567;
  assign G3366 = G2567;
  assign G3382 = G2589;
  assign G3390 = G2589;
  assign G397 = G2657 & G330 & G2514;
  assign G2544 = G330 & G2508;
  assign G2562 = ~G3290 | ~G3293;
  assign G2584 = ~G3308 | ~G3311;
  assign G3402 = ~G3398;
  assign G2626 = ~G2624 | ~G2625;
  assign G2632 = ~G2629;
  assign G2634 = G2501 & G2629;
  assign G2650 = G2647;
  assign G3268 = ~G3264;
  assign G3256 = G2508;
  assign G3285 = ~G3280 | ~G3283;
  assign G3321 = ~G3316 | ~G3319;
  assign G3371 = ~G3303 | ~G3304;
  assign G3403 = G2609;
  assign G3411 = G2609;
  assign G362 = G938 | G929 | G933;
  assign G1030 = ~G938 & ~G929 & ~G933;
  assign G399 = G397 | G398;
  assign G2564 = ~G2562 | ~G2563;
  assign G3362 = ~G3358;
  assign G3370 = ~G3366;
  assign G2586 = ~G2584 | ~G2585;
  assign G3386 = ~G3382;
  assign G3394 = ~G3390;
  assign G2633 = G2632 & G330 & G2505;
  assign G3261 = G2527;
  assign G3269 = G2527;
  assign G3347 = ~G3285 | ~G3286;
  assign G3395 = ~G3321 | ~G3322;
  assign G363 = ~G1030;
  assign G2536 = ~G3256 | ~G3259;
  assign G3260 = ~G3256;
  assign G3377 = ~G3371;
  assign G2580 = ~G3371 | ~G3378;
  assign G3409 = ~G3403;
  assign G2616 = ~G3403 | ~G3410;
  assign G3417 = ~G3411;
  assign G2622 = ~G3411 | ~G3418;
  assign G2635 = ~G2633 & ~G2634;
  assign G2805 = G2626 & G2802;
  assign G2808 = G2626 & G2803;
  assign G3334 = G2544;
  assign G3342 = G2544;
  assign G3454 = G2650;
  assign G364 = G362 & G363;
  assign G2537 = ~G3253 | ~G3260;
  assign G3275 = ~G3269;
  assign G2540 = ~G3269 | ~G3276;
  assign G3353 = ~G3347;
  assign G2557 = ~G3347 | ~G3354;
  assign G2579 = ~G3374 | ~G3377;
  assign G3401 = ~G3395;
  assign G2602 = ~G3395 | ~G3402;
  assign G2615 = ~G3406 | ~G3409;
  assign G2621 = ~G3414 | ~G3417;
  assign G3267 = ~G3261;
  assign G3112 = ~G3261 | ~G3268;
  assign G3355 = G2564;
  assign G3363 = G2564;
  assign G3379 = G2586;
  assign G3387 = G2586;
  assign G2538 = ~G2536 | ~G2537;
  assign G2539 = ~G3272 | ~G3275;
  assign G3338 = ~G3334;
  assign G3346 = ~G3342;
  assign G2556 = ~G3350 | ~G3353;
  assign G2581 = ~G2579 | ~G2580;
  assign G2601 = ~G3398 | ~G3401;
  assign G2617 = ~G2615 | ~G2616;
  assign G2623 = ~G2621 | ~G2622;
  assign G2638 = G2635;
  assign G3458 = ~G3454;
  assign G2814 = G2811 | G2805 | G2808;
  assign G2816 = ~G2811 & ~G2805 & ~G2808;
  assign G3111 = ~G3264 | ~G3267;
  assign G2541 = ~G2539 | ~G2540;
  assign G2558 = ~G2556 | ~G2557;
  assign G3361 = ~G3355;
  assign G2571 = ~G3355 | ~G3362;
  assign G3369 = ~G3363;
  assign G2577 = ~G3363 | ~G3370;
  assign G3385 = ~G3379;
  assign G2593 = ~G3379 | ~G3386;
  assign G3393 = ~G3387;
  assign G2598 = ~G3387 | ~G3394;
  assign G2603 = ~G2601 | ~G2602;
  assign G3113 = ~G3111 | ~G3112;
  assign G3116 = G330 & G2538;
  assign G3451 = ~G2623;
  assign G395 = ~G2816;
  assign G2570 = ~G3358 | ~G3361;
  assign G2576 = ~G3366 | ~G3369;
  assign G2592 = ~G3382 | ~G3385;
  assign G2597 = ~G3390 | ~G3393;
  assign G2736 = G2581 & G2733;
  assign G2739 = G2581 & G2734;
  assign G2788 = G2617 & G2785;
  assign G3438 = G2638;
  assign G3446 = G2617 & G2647;
  assign G3459 = G2814;
  assign G396 = G2814 & G395;
  assign G3119 = ~G3113;
  assign G3120 = ~G3116;
  assign G2572 = ~G2570 | ~G2571;
  assign G2578 = ~G2576 | ~G2577;
  assign G2594 = ~G2592 | ~G2593;
  assign G2599 = ~G2597 | ~G2598;
  assign G2677 = ~G3451 | ~G3458;
  assign G3457 = ~G3451;
  assign G2700 = G2558 & G2697;
  assign G2771 = G2603 & G2768;
  assign G3331 = G2541;
  assign G3339 = G2541;
  assign G3427 = G2558;
  assign G3443 = G2603;
  assign G954 = ~G3116 | ~G3119;
  assign G955 = ~G3113 | ~G3120;
  assign G2600 = ~G2599;
  assign G3442 = ~G3438;
  assign G3450 = ~G3446;
  assign G2676 = ~G3454 | ~G3457;
  assign G2745 = G2742 | G2736 | G2739;
  assign G2748 = ~G2742 & ~G2736 & ~G2739;
  assign G3465 = ~G3459;
  assign G3435 = ~G2578;
  assign G950 = ~G954 | ~G955;
  assign G3337 = ~G3331;
  assign G2548 = ~G3331 | ~G3338;
  assign G3345 = ~G3339;
  assign G2553 = ~G3339 | ~G3346;
  assign G2661 = ~G2600 & ~G2650;
  assign G2662 = G2650 & G2594 & G2617 & G2603;
  assign G3433 = ~G3427;
  assign G3449 = ~G3443;
  assign G2672 = ~G3443 | ~G3450;
  assign G2674 = ~G2676 | ~G2677;
  assign G2719 = G2572 & G2716;
  assign G2754 = G2594 & G2751;
  assign G3430 = G2572 & G2635;
  assign G383 = ~G2748;
  assign G951 = G950 & G943;
  assign G2547 = ~G3334 | ~G3337;
  assign G2552 = ~G3342 | ~G3345;
  assign G2663 = G2661 | G2662;
  assign G2670 = ~G3435 | ~G3442;
  assign G3441 = ~G3435;
  assign G2671 = ~G3446 | ~G3449;
  assign G2675 = ~G2674;
  assign G3491 = G2745;
  assign G3499 = G2745;
  assign G384 = G2745 & G383;
  assign G2549 = ~G2547 | ~G2548;
  assign G2554 = ~G2552 | ~G2553;
  assign G2664 = ~G3430 | ~G3433;
  assign G3434 = ~G3430;
  assign G2669 = ~G3438 | ~G3441;
  assign G2673 = ~G2671 | ~G2672;
  assign G2757 = G2663 & G2752;
  assign G2791 = G2675 & G2786;
  assign G365 = G951 | G944 | G947;
  assign G1031 = ~G951 & ~G944 & ~G947;
  assign G2555 = ~G2554;
  assign G2665 = ~G3427 | ~G3434;
  assign G2667 = ~G2669 | ~G2670;
  assign G2774 = G2673 & G2769;
  assign G3497 = ~G3491;
  assign G3505 = ~G3499;
  assign G366 = ~G1031;
  assign G2658 = ~G2555 & ~G2638;
  assign G2659 = G2638 & G2549 & G2572 & G2558;
  assign G2666 = ~G2664 | ~G2665;
  assign G2668 = ~G2667;
  assign G2681 = G2549 & G2678;
  assign G2763 = G2760 | G2754 | G2757;
  assign G2765 = ~G2760 & ~G2754 & ~G2757;
  assign G2797 = G2794 | G2788 | G2791;
  assign G2799 = ~G2794 & ~G2788 & ~G2791;
  assign G367 = G365 & G366;
  assign G2660 = G2658 | G2659;
  assign G2703 = G2666 & G2698;
  assign G2722 = G2668 & G2717;
  assign G2780 = G2777 | G2771 | G2774;
  assign G2782 = ~G2777 & ~G2771 & ~G2774;
  assign G386 = ~G2765;
  assign G392 = ~G2799;
  assign G2684 = G2660 & G2679;
  assign G3462 = G2797;
  assign G3470 = G2763;
  assign G387 = G2763 & G386;
  assign G389 = ~G2782;
  assign G393 = G2797 & G392;
  assign G2709 = G2706 | G2700 | G2703;
  assign G2713 = ~G2706 & ~G2700 & ~G2703;
  assign G2728 = G2725 | G2719 | G2722;
  assign G2730 = ~G2725 & ~G2719 & ~G2722;
  assign G2922 = G2765 & G2782 & G2816 & G2799;
  assign G3467 = G2780;
  assign G390 = G2780 & G389;
  assign G2690 = G2687 | G2681 | G2684;
  assign G2694 = ~G2687 & ~G2681 & ~G2684;
  assign G2821 = ~G3462 | ~G3465;
  assign G3466 = ~G3462;
  assign G3474 = ~G3470;
  assign G378 = G2709 & G2709;
  assign G380 = ~G2730;
  assign G2822 = ~G3459 | ~G3466;
  assign G3473 = ~G3467;
  assign G2827 = ~G3467 | ~G3474;
  assign G2839 = G2728;
  assign G2883 = G2709 & G2871;
  assign G3507 = G2709;
  assign G375 = G2690 & G2690;
  assign G381 = G2728 & G380;
  assign G2823 = ~G2821 | ~G2822;
  assign G2826 = ~G3470 | ~G3473;
  assign G2880 = G2871 & G2690;
  assign G2925 = G2694 & G2713 & G2748 & G2730;
  assign G2928 = G2874 & G2713 & G2694;
  assign G3510 = G2690;
  assign G2828 = ~G2826 | ~G2827;
  assign G3494 = G2839;
  assign G3502 = G2839;
  assign G3513 = ~G3507;
  assign G3544 = G2883;
  assign G3552 = G2883;
  assign G406 = G2922 & G2925;
  assign G2929 = G2922 & G2925;
  assign G3475 = G2823;
  assign G3483 = G2823;
  assign G3514 = ~G3510;
  assign G3515 = ~G3510 | ~G3513;
  assign G3541 = G2880;
  assign G3549 = G2880;
  assign G407 = ~G406;
  assign G2930 = ~G2928 & ~G2929;
  assign G2842 = ~G3494 | ~G3497;
  assign G3498 = ~G3494;
  assign G2852 = ~G3502 | ~G3505;
  assign G3506 = ~G3502;
  assign G3548 = ~G3544;
  assign G3556 = ~G3552;
  assign G3478 = G2828;
  assign G3486 = G2828;
  assign G3516 = ~G3507 | ~G3514;
  assign G408 = G213 & G2930;
  assign G3481 = ~G3475;
  assign G3489 = ~G3483;
  assign G2843 = ~G3491 | ~G3498;
  assign G2853 = ~G3499 | ~G3506;
  assign G3547 = ~G3541;
  assign G2887 = ~G3541 | ~G3548;
  assign G2896 = ~G3549 | ~G3556;
  assign G3555 = ~G3549;
  assign G3520 = ~G3515 | ~G3516;
  assign G409 = ~G408;
  assign G2831 = ~G3478 | ~G3481;
  assign G3482 = ~G3478;
  assign G2836 = ~G3486 | ~G3489;
  assign G3490 = ~G3486;
  assign G2844 = ~G2842 | ~G2843;
  assign G2848 = ~G2852 | ~G2853;
  assign G2886 = ~G3544 | ~G3547;
  assign G2895 = ~G3552 | ~G3555;
  assign G2832 = ~G3475 | ~G3482;
  assign G2837 = ~G3483 | ~G3490;
  assign G2849 = ~G2848;
  assign G3524 = ~G3520;
  assign G2888 = ~G2886 | ~G2887;
  assign G2891 = ~G2895 | ~G2896;
  assign G2833 = ~G2831 | ~G2832;
  assign G2838 = ~G2836 | ~G2837;
  assign G2892 = ~G2891;
  assign G3517 = G2844;
  assign G2906 = G2900 & G2844 & G2888;
  assign G2908 = G2903 & G2849 & G2888;
  assign G2913 = ~G2838;
  assign G3523 = ~G3517;
  assign G2855 = ~G3517 | ~G3524;
  assign G2907 = G2903 & G2844 & G2892;
  assign G2909 = G2900 & G2849 & G2892;
  assign G3525 = G2833;
  assign G3533 = G2833;
  assign G2854 = ~G3520 | ~G3523;
  assign G2910 = G2909 | G2908 | G2906 | G2907;
  assign G3560 = G2913;
  assign G3568 = G2913;
  assign G2856 = ~G2854 | ~G2855;
  assign G3539 = ~G3533;
  assign G3531 = ~G3525;
  assign G3572 = ~G3568;
  assign G3564 = ~G3560;
  assign G3557 = G2910;
  assign G3565 = G2910;
  assign G3528 = G2856;
  assign G3536 = G2856;
  assign G2921 = ~G3557 | ~G3564;
  assign G2917 = ~G3565 | ~G3572;
  assign G3571 = ~G3565;
  assign G3563 = ~G3557;
  assign G2863 = ~G3528 | ~G3531;
  assign G2859 = ~G3536 | ~G3539;
  assign G2920 = ~G3560 | ~G3563;
  assign G2916 = ~G3568 | ~G3571;
  assign G3540 = ~G3536;
  assign G3532 = ~G3528;
  assign G2864 = ~G3525 | ~G3532;
  assign G2860 = ~G3533 | ~G3540;
  assign G403 = ~G2920 | ~G2921;
  assign G404 = ~G2916 | ~G2917;
  assign G400 = ~G2863 | ~G2864;
  assign G401 = ~G2859 | ~G2860;
  assign G405 = G403 & G404;
  assign G402 = ~G400 | ~G401;
endmodule


