// Benchmark "c880" written by ABC on Thu Mar  5 01:08:09 2020

module c880 ( 
    G1GAT, G8GAT, G13GAT, G17GAT, G26GAT, G29GAT, G36GAT, G42GAT, G51GAT,
    G55GAT, G59GAT, G68GAT, G72GAT, G73GAT, G74GAT, G75GAT, G80GAT, G85GAT,
    G86GAT, G87GAT, G88GAT, G89GAT, G90GAT, G91GAT, G96GAT, G101GAT,
    G106GAT, G111GAT, G116GAT, G121GAT, G126GAT, G130GAT, G135GAT, G138GAT,
    G143GAT, G146GAT, G149GAT, G152GAT, G153GAT, G156GAT, G159GAT, G165GAT,
    G171GAT, G177GAT, G183GAT, G189GAT, G195GAT, G201GAT, G207GAT, G210GAT,
    G219GAT, G228GAT, G237GAT, G246GAT, G255GAT, G259GAT, G260GAT, G261GAT,
    G267GAT, G268GAT,
    G388GAT, G389GAT, G390GAT, G391GAT, G418GAT, G419GAT, G420GAT, G421GAT,
    G422GAT, G423GAT, G446GAT, G447GAT, G448GAT, G449GAT, G450GAT, G767GAT,
    G768GAT, G850GAT, G863GAT, G864GAT, G865GAT, G866GAT, G874GAT, G878GAT,
    G879GAT, G880GAT  );
  input  G1GAT, G8GAT, G13GAT, G17GAT, G26GAT, G29GAT, G36GAT, G42GAT,
    G51GAT, G55GAT, G59GAT, G68GAT, G72GAT, G73GAT, G74GAT, G75GAT, G80GAT,
    G85GAT, G86GAT, G87GAT, G88GAT, G89GAT, G90GAT, G91GAT, G96GAT,
    G101GAT, G106GAT, G111GAT, G116GAT, G121GAT, G126GAT, G130GAT, G135GAT,
    G138GAT, G143GAT, G146GAT, G149GAT, G152GAT, G153GAT, G156GAT, G159GAT,
    G165GAT, G171GAT, G177GAT, G183GAT, G189GAT, G195GAT, G201GAT, G207GAT,
    G210GAT, G219GAT, G228GAT, G237GAT, G246GAT, G255GAT, G259GAT, G260GAT,
    G261GAT, G267GAT, G268GAT;
  output G388GAT, G389GAT, G390GAT, G391GAT, G418GAT, G419GAT, G420GAT,
    G421GAT, G422GAT, G423GAT, G446GAT, G447GAT, G448GAT, G449GAT, G450GAT,
    G767GAT, G768GAT, G850GAT, G863GAT, G864GAT, G865GAT, G866GAT, G874GAT,
    G878GAT, G879GAT, G880GAT;
  wire G269GAT, G270GAT, G273GAT, G276GAT, G279GAT, G280GAT, G284GAT,
    G285GAT, G286GAT, G287GAT, G290GAT, G291GAT, G292GAT, G293GAT, G294GAT,
    G295GAT, G296GAT, G297GAT, G298GAT, G301GAT, G302GAT, G303GAT, G304GAT,
    G305GAT, G306GAT, G307GAT, G308GAT, G309GAT, G310GAT, G316GAT, G317GAT,
    G318GAT, G319GAT, G322GAT, G323GAT, G324GAT, G325GAT, G326GAT, G327GAT,
    G328GAT, G329GAT, G330GAT, G331GAT, G332GAT, G333GAT, G334GAT, G335GAT,
    G336GAT, G337GAT, G338GAT, G339GAT, G340GAT, G341GAT, G342GAT, G343GAT,
    G344GAT, G345GAT, G346GAT, G347GAT, G348GAT, G349GAT, G350GAT, G351GAT,
    G352GAT, G353GAT, G354GAT, G355GAT, G356GAT, G357GAT, G360GAT, G363GAT,
    G366GAT, G369GAT, G375GAT, G376GAT, G379GAT, G382GAT, G385GAT, G392GAT,
    G393GAT, G399GAT, G400GAT, G401GAT, G402GAT, G403GAT, G404GAT, G405GAT,
    G406GAT, G407GAT, G408GAT, G409GAT, G410GAT, G411GAT, G412GAT, G413GAT,
    G414GAT, G415GAT, G416GAT, G417GAT, G424GAT, G425GAT, G426GAT, G427GAT,
    G432GAT, G437GAT, G442GAT, G443GAT, G444GAT, G445GAT, G451GAT, G460GAT,
    G463GAT, G466GAT, G475GAT, G476GAT, G477GAT, G478GAT, G479GAT, G480GAT,
    G481GAT, G482GAT, G483GAT, G488GAT, G489GAT, G490GAT, G491GAT, G492GAT,
    G495GAT, G498GAT, G499GAT, G500GAT, G501GAT, G502GAT, G503GAT, G504GAT,
    G505GAT, G506GAT, G507GAT, G508GAT, G509GAT, G510GAT, G511GAT, G512GAT,
    G513GAT, G514GAT, G515GAT, G516GAT, G517GAT, G518GAT, G519GAT, G520GAT,
    G521GAT, G522GAT, G523GAT, G524GAT, G525GAT, G526GAT, G527GAT, G528GAT,
    G529GAT, G530GAT, G533GAT, G536GAT, G537GAT, G538GAT, G539GAT, G540GAT,
    G541GAT, G542GAT, G543GAT, G544GAT, G547GAT, G550GAT, G551GAT, G552GAT,
    G553GAT, G557GAT, G561GAT, G565GAT, G569GAT, G573GAT, G577GAT, G581GAT,
    G585GAT, G586GAT, G587GAT, G588GAT, G589GAT, G590GAT, G593GAT, G596GAT,
    G597GAT, G600GAT, G605GAT, G606GAT, G609GAT, G615GAT, G616GAT, G619GAT,
    G624GAT, G625GAT, G628GAT, G631GAT, G632GAT, G635GAT, G640GAT, G641GAT,
    G644GAT, G650GAT, G651GAT, G654GAT, G659GAT, G660GAT, G661GAT, G662GAT,
    G665GAT, G669GAT, G670GAT, G673GAT, G677GAT, G678GAT, G682GAT, G686GAT,
    G687GAT, G692GAT, G696GAT, G697GAT, G700GAT, G704GAT, G705GAT, G708GAT,
    G712GAT, G713GAT, G717GAT, G721GAT, G722GAT, G727GAT, G731GAT, G732GAT,
    G733GAT, G734GAT, G735GAT, G736GAT, G737GAT, G738GAT, G739GAT, G740GAT,
    G741GAT, G742GAT, G743GAT, G744GAT, G745GAT, G746GAT, G747GAT, G748GAT,
    G749GAT, G750GAT, G751GAT, G752GAT, G753GAT, G754GAT, G755GAT, G756GAT,
    G757GAT, G758GAT, G759GAT, G760GAT, G761GAT, G762GAT, G763GAT, G764GAT,
    G765GAT, G766GAT, G769GAT, G770GAT, G771GAT, G772GAT, G773GAT, G777GAT,
    G778GAT, G781GAT, G782GAT, G785GAT, G786GAT, G787GAT, G788GAT, G789GAT,
    G790GAT, G791GAT, G792GAT, G793GAT, G794GAT, G795GAT, G796GAT, G802GAT,
    G803GAT, G804GAT, G805GAT, G806GAT, G807GAT, G808GAT, G809GAT, G810GAT,
    G811GAT, G812GAT, G813GAT, G814GAT, G815GAT, G819GAT, G822GAT, G825GAT,
    G826GAT, G827GAT, G828GAT, G829GAT, G830GAT, G831GAT, G832GAT, G833GAT,
    G834GAT, G835GAT, G836GAT, G837GAT, G838GAT, G839GAT, G840GAT, G841GAT,
    G842GAT, G843GAT, G844GAT, G845GAT, G846GAT, G847GAT, G848GAT, G849GAT,
    G851GAT, G852GAT, G853GAT, G854GAT, G855GAT, G856GAT, G857GAT, G858GAT,
    G859GAT, G860GAT, G861GAT, G862GAT, G867GAT, G868GAT, G869GAT, G870GAT,
    G871GAT, G872GAT, G873GAT, G875GAT, G876GAT, G877GAT;
  assign G269GAT = ~G17GAT | ~G13GAT | ~G1GAT | ~G8GAT;
  assign G270GAT = ~G17GAT | ~G13GAT | ~G1GAT | ~G26GAT;
  assign G273GAT = G42GAT & G29GAT & G36GAT;
  assign G276GAT = G51GAT & G1GAT & G26GAT;
  assign G279GAT = ~G17GAT | ~G51GAT | ~G1GAT | ~G8GAT;
  assign G280GAT = ~G55GAT | ~G13GAT | ~G1GAT | ~G8GAT;
  assign G284GAT = ~G72GAT | ~G68GAT | ~G59GAT | ~G42GAT;
  assign G285GAT = ~G29GAT | ~G68GAT;
  assign G286GAT = ~G74GAT | ~G59GAT | ~G68GAT;
  assign G287GAT = G80GAT & G29GAT & G75GAT;
  assign G290GAT = G42GAT & G29GAT & G75GAT;
  assign G291GAT = G80GAT & G29GAT & G36GAT;
  assign G292GAT = G42GAT & G29GAT & G36GAT;
  assign G293GAT = G80GAT & G59GAT & G75GAT;
  assign G294GAT = G42GAT & G59GAT & G75GAT;
  assign G295GAT = G80GAT & G59GAT & G36GAT;
  assign G296GAT = G42GAT & G59GAT & G36GAT;
  assign G297GAT = G85GAT & G86GAT;
  assign G298GAT = G87GAT | G88GAT;
  assign G301GAT = ~G91GAT | ~G96GAT;
  assign G302GAT = G91GAT | G96GAT;
  assign G303GAT = ~G101GAT | ~G106GAT;
  assign G304GAT = G101GAT | G106GAT;
  assign G305GAT = ~G111GAT | ~G116GAT;
  assign G306GAT = G111GAT | G116GAT;
  assign G307GAT = ~G121GAT | ~G126GAT;
  assign G308GAT = G121GAT | G126GAT;
  assign G309GAT = G8GAT & G138GAT;
  assign G310GAT = ~G268GAT;
  assign G316GAT = G51GAT & G138GAT;
  assign G317GAT = G17GAT & G138GAT;
  assign G318GAT = G152GAT & G138GAT;
  assign G319GAT = ~G59GAT | ~G156GAT;
  assign G322GAT = ~G17GAT & ~G42GAT;
  assign G323GAT = G17GAT & G42GAT;
  assign G324GAT = ~G159GAT | ~G165GAT;
  assign G325GAT = G159GAT | G165GAT;
  assign G326GAT = ~G171GAT | ~G177GAT;
  assign G327GAT = G171GAT | G177GAT;
  assign G328GAT = ~G183GAT | ~G189GAT;
  assign G329GAT = G183GAT | G189GAT;
  assign G330GAT = ~G195GAT | ~G201GAT;
  assign G331GAT = G195GAT | G201GAT;
  assign G332GAT = G210GAT & G91GAT;
  assign G333GAT = G210GAT & G96GAT;
  assign G334GAT = G210GAT & G101GAT;
  assign G335GAT = G210GAT & G106GAT;
  assign G336GAT = G210GAT & G111GAT;
  assign G337GAT = G255GAT & G259GAT;
  assign G338GAT = G210GAT & G116GAT;
  assign G339GAT = G255GAT & G260GAT;
  assign G340GAT = G210GAT & G121GAT;
  assign G341GAT = G255GAT & G267GAT;
  assign G342GAT = ~G269GAT;
  assign G343GAT = ~G273GAT;
  assign G344GAT = G270GAT | G273GAT;
  assign G345GAT = ~G276GAT;
  assign G346GAT = ~G276GAT;
  assign G347GAT = ~G279GAT;
  assign G348GAT = ~G280GAT & ~G284GAT;
  assign G349GAT = G280GAT | G285GAT;
  assign G350GAT = G280GAT | G286GAT;
  assign G351GAT = ~G293GAT;
  assign G352GAT = ~G294GAT;
  assign G353GAT = ~G295GAT;
  assign G354GAT = ~G296GAT;
  assign G355GAT = ~G89GAT | ~G298GAT;
  assign G356GAT = G90GAT & G298GAT;
  assign G357GAT = ~G301GAT | ~G302GAT;
  assign G360GAT = ~G303GAT | ~G304GAT;
  assign G363GAT = ~G305GAT | ~G306GAT;
  assign G366GAT = ~G307GAT | ~G308GAT;
  assign G369GAT = ~G310GAT;
  assign G375GAT = ~G322GAT & ~G323GAT;
  assign G376GAT = ~G324GAT | ~G325GAT;
  assign G379GAT = ~G326GAT | ~G327GAT;
  assign G382GAT = ~G328GAT | ~G329GAT;
  assign G385GAT = ~G330GAT | ~G331GAT;
  assign G388GAT = G290GAT;
  assign G389GAT = G291GAT;
  assign G390GAT = G292GAT;
  assign G391GAT = G297GAT;
  assign G392GAT = G270GAT | G343GAT;
  assign G393GAT = ~G345GAT;
  assign G399GAT = ~G346GAT;
  assign G400GAT = G348GAT & G73GAT;
  assign G401GAT = ~G349GAT;
  assign G402GAT = ~G350GAT;
  assign G403GAT = ~G355GAT;
  assign G404GAT = ~G357GAT;
  assign G405GAT = ~G360GAT;
  assign G406GAT = G357GAT & G360GAT;
  assign G407GAT = ~G363GAT;
  assign G408GAT = ~G366GAT;
  assign G409GAT = G363GAT & G366GAT;
  assign G410GAT = ~G347GAT | ~G352GAT;
  assign G411GAT = ~G376GAT;
  assign G412GAT = ~G379GAT;
  assign G413GAT = G376GAT & G379GAT;
  assign G414GAT = ~G382GAT;
  assign G415GAT = ~G385GAT;
  assign G416GAT = G382GAT & G385GAT;
  assign G417GAT = G210GAT & G369GAT;
  assign G418GAT = G342GAT;
  assign G419GAT = G344GAT;
  assign G420GAT = G351GAT;
  assign G421GAT = G353GAT;
  assign G422GAT = G354GAT;
  assign G423GAT = G356GAT;
  assign G424GAT = ~G400GAT;
  assign G425GAT = G404GAT & G405GAT;
  assign G426GAT = G407GAT & G408GAT;
  assign G427GAT = G55GAT & G319GAT & G393GAT;
  assign G432GAT = G287GAT & G393GAT & G17GAT;
  assign G437GAT = ~G55GAT | ~G393GAT | ~G287GAT;
  assign G442GAT = ~G393GAT | ~G156GAT | ~G375GAT | ~G59GAT;
  assign G443GAT = ~G17GAT | ~G393GAT | ~G319GAT;
  assign G444GAT = G411GAT & G412GAT;
  assign G445GAT = G414GAT & G415GAT;
  assign G446GAT = G392GAT;
  assign G447GAT = G399GAT;
  assign G448GAT = G401GAT;
  assign G449GAT = G402GAT;
  assign G450GAT = G403GAT;
  assign G451GAT = ~G424GAT;
  assign G460GAT = ~G406GAT & ~G425GAT;
  assign G463GAT = ~G409GAT & ~G426GAT;
  assign G466GAT = ~G442GAT | ~G410GAT;
  assign G475GAT = G143GAT & G427GAT;
  assign G476GAT = G310GAT & G432GAT;
  assign G477GAT = G146GAT & G427GAT;
  assign G478GAT = G310GAT & G432GAT;
  assign G479GAT = G149GAT & G427GAT;
  assign G480GAT = G310GAT & G432GAT;
  assign G481GAT = G153GAT & G427GAT;
  assign G482GAT = G310GAT & G432GAT;
  assign G483GAT = ~G443GAT | ~G1GAT;
  assign G488GAT = G369GAT | G437GAT;
  assign G489GAT = G369GAT | G437GAT;
  assign G490GAT = G369GAT | G437GAT;
  assign G491GAT = G369GAT | G437GAT;
  assign G492GAT = ~G413GAT & ~G444GAT;
  assign G495GAT = ~G416GAT & ~G445GAT;
  assign G498GAT = ~G130GAT | ~G460GAT;
  assign G499GAT = G130GAT | G460GAT;
  assign G500GAT = ~G463GAT | ~G135GAT;
  assign G501GAT = G463GAT | G135GAT;
  assign G502GAT = G91GAT & G466GAT;
  assign G503GAT = ~G475GAT & ~G476GAT;
  assign G504GAT = G96GAT & G466GAT;
  assign G505GAT = ~G477GAT & ~G478GAT;
  assign G506GAT = G101GAT & G466GAT;
  assign G507GAT = ~G479GAT & ~G480GAT;
  assign G508GAT = G106GAT & G466GAT;
  assign G509GAT = ~G481GAT & ~G482GAT;
  assign G510GAT = G143GAT & G483GAT;
  assign G511GAT = G111GAT & G466GAT;
  assign G512GAT = G146GAT & G483GAT;
  assign G513GAT = G116GAT & G466GAT;
  assign G514GAT = G149GAT & G483GAT;
  assign G515GAT = G121GAT & G466GAT;
  assign G516GAT = G153GAT & G483GAT;
  assign G517GAT = G126GAT & G466GAT;
  assign G518GAT = ~G130GAT | ~G492GAT;
  assign G519GAT = G130GAT | G492GAT;
  assign G520GAT = ~G495GAT | ~G207GAT;
  assign G521GAT = G495GAT | G207GAT;
  assign G522GAT = G451GAT & G159GAT;
  assign G523GAT = G451GAT & G165GAT;
  assign G524GAT = G451GAT & G171GAT;
  assign G525GAT = G451GAT & G177GAT;
  assign G526GAT = G451GAT & G183GAT;
  assign G527GAT = ~G451GAT | ~G189GAT;
  assign G528GAT = ~G451GAT | ~G195GAT;
  assign G529GAT = ~G451GAT | ~G201GAT;
  assign G530GAT = ~G498GAT | ~G499GAT;
  assign G533GAT = ~G500GAT | ~G501GAT;
  assign G536GAT = ~G309GAT & ~G502GAT;
  assign G537GAT = ~G316GAT & ~G504GAT;
  assign G538GAT = ~G317GAT & ~G506GAT;
  assign G539GAT = ~G318GAT & ~G508GAT;
  assign G540GAT = ~G510GAT & ~G511GAT;
  assign G541GAT = ~G512GAT & ~G513GAT;
  assign G542GAT = ~G514GAT & ~G515GAT;
  assign G543GAT = ~G516GAT & ~G517GAT;
  assign G544GAT = ~G518GAT | ~G519GAT;
  assign G547GAT = ~G520GAT | ~G521GAT;
  assign G550GAT = ~G530GAT;
  assign G551GAT = ~G533GAT;
  assign G552GAT = G530GAT & G533GAT;
  assign G553GAT = ~G536GAT | ~G503GAT;
  assign G557GAT = ~G537GAT | ~G505GAT;
  assign G561GAT = ~G538GAT | ~G507GAT;
  assign G565GAT = ~G539GAT | ~G509GAT;
  assign G569GAT = ~G488GAT | ~G540GAT;
  assign G573GAT = ~G489GAT | ~G541GAT;
  assign G577GAT = ~G490GAT | ~G542GAT;
  assign G581GAT = ~G491GAT | ~G543GAT;
  assign G585GAT = ~G544GAT;
  assign G586GAT = ~G547GAT;
  assign G587GAT = G544GAT & G547GAT;
  assign G588GAT = G550GAT & G551GAT;
  assign G589GAT = G585GAT & G586GAT;
  assign G590GAT = ~G553GAT | ~G159GAT;
  assign G593GAT = G553GAT | G159GAT;
  assign G596GAT = G246GAT & G553GAT;
  assign G597GAT = ~G557GAT | ~G165GAT;
  assign G600GAT = G557GAT | G165GAT;
  assign G605GAT = G246GAT & G557GAT;
  assign G606GAT = ~G561GAT | ~G171GAT;
  assign G609GAT = G561GAT | G171GAT;
  assign G615GAT = G246GAT & G561GAT;
  assign G616GAT = ~G565GAT | ~G177GAT;
  assign G619GAT = G565GAT | G177GAT;
  assign G624GAT = G246GAT & G565GAT;
  assign G625GAT = ~G569GAT | ~G183GAT;
  assign G628GAT = G569GAT | G183GAT;
  assign G631GAT = G246GAT & G569GAT;
  assign G632GAT = ~G573GAT | ~G189GAT;
  assign G635GAT = G573GAT | G189GAT;
  assign G640GAT = G246GAT & G573GAT;
  assign G641GAT = ~G577GAT | ~G195GAT;
  assign G644GAT = G577GAT | G195GAT;
  assign G650GAT = G246GAT & G577GAT;
  assign G651GAT = ~G581GAT | ~G201GAT;
  assign G654GAT = G581GAT | G201GAT;
  assign G659GAT = G246GAT & G581GAT;
  assign G660GAT = ~G552GAT & ~G588GAT;
  assign G661GAT = ~G587GAT & ~G589GAT;
  assign G662GAT = ~G590GAT;
  assign G665GAT = G593GAT & G590GAT;
  assign G669GAT = ~G596GAT & ~G522GAT;
  assign G670GAT = ~G597GAT;
  assign G673GAT = G600GAT & G597GAT;
  assign G677GAT = ~G605GAT & ~G523GAT;
  assign G678GAT = ~G606GAT;
  assign G682GAT = G609GAT & G606GAT;
  assign G686GAT = ~G615GAT & ~G524GAT;
  assign G687GAT = ~G616GAT;
  assign G692GAT = G619GAT & G616GAT;
  assign G696GAT = ~G624GAT & ~G525GAT;
  assign G697GAT = ~G625GAT;
  assign G700GAT = G628GAT & G625GAT;
  assign G704GAT = ~G631GAT & ~G526GAT;
  assign G705GAT = ~G632GAT;
  assign G708GAT = G635GAT & G632GAT;
  assign G712GAT = ~G337GAT & ~G640GAT;
  assign G713GAT = ~G641GAT;
  assign G717GAT = G644GAT & G641GAT;
  assign G721GAT = ~G339GAT & ~G650GAT;
  assign G722GAT = ~G651GAT;
  assign G727GAT = G654GAT & G651GAT;
  assign G731GAT = ~G341GAT & ~G659GAT;
  assign G732GAT = ~G654GAT | ~G261GAT;
  assign G733GAT = ~G261GAT | ~G644GAT | ~G654GAT;
  assign G734GAT = ~G261GAT | ~G654GAT | ~G635GAT | ~G644GAT;
  assign G735GAT = ~G662GAT;
  assign G736GAT = G228GAT & G665GAT;
  assign G737GAT = G237GAT & G662GAT;
  assign G738GAT = ~G670GAT;
  assign G739GAT = G228GAT & G673GAT;
  assign G740GAT = G237GAT & G670GAT;
  assign G741GAT = ~G678GAT;
  assign G742GAT = G228GAT & G682GAT;
  assign G743GAT = G237GAT & G678GAT;
  assign G744GAT = ~G687GAT;
  assign G745GAT = G228GAT & G692GAT;
  assign G746GAT = G237GAT & G687GAT;
  assign G747GAT = ~G697GAT;
  assign G748GAT = G228GAT & G700GAT;
  assign G749GAT = G237GAT & G697GAT;
  assign G750GAT = ~G705GAT;
  assign G751GAT = G228GAT & G708GAT;
  assign G752GAT = G237GAT & G705GAT;
  assign G753GAT = ~G713GAT;
  assign G754GAT = G228GAT & G717GAT;
  assign G755GAT = G237GAT & G713GAT;
  assign G756GAT = ~G722GAT;
  assign G757GAT = ~G727GAT & ~G261GAT;
  assign G758GAT = G727GAT & G261GAT;
  assign G759GAT = G228GAT & G727GAT;
  assign G760GAT = G237GAT & G722GAT;
  assign G761GAT = ~G644GAT | ~G722GAT;
  assign G762GAT = ~G635GAT | ~G713GAT;
  assign G763GAT = ~G722GAT | ~G635GAT | ~G644GAT;
  assign G764GAT = ~G609GAT | ~G687GAT;
  assign G765GAT = ~G600GAT | ~G678GAT;
  assign G766GAT = ~G687GAT | ~G600GAT | ~G609GAT;
  assign G767GAT = G660GAT;
  assign G768GAT = G661GAT;
  assign G769GAT = ~G736GAT & ~G737GAT;
  assign G770GAT = ~G739GAT & ~G740GAT;
  assign G771GAT = ~G742GAT & ~G743GAT;
  assign G772GAT = ~G745GAT & ~G746GAT;
  assign G773GAT = ~G734GAT | ~G763GAT | ~G750GAT | ~G762GAT;
  assign G777GAT = ~G748GAT & ~G749GAT;
  assign G778GAT = ~G733GAT | ~G753GAT | ~G761GAT;
  assign G781GAT = ~G751GAT & ~G752GAT;
  assign G782GAT = ~G756GAT | ~G732GAT;
  assign G785GAT = ~G754GAT & ~G755GAT;
  assign G786GAT = ~G757GAT & ~G758GAT;
  assign G787GAT = ~G759GAT & ~G760GAT;
  assign G788GAT = ~G700GAT & ~G773GAT;
  assign G789GAT = G700GAT & G773GAT;
  assign G790GAT = ~G708GAT & ~G778GAT;
  assign G791GAT = G708GAT & G778GAT;
  assign G792GAT = ~G717GAT & ~G782GAT;
  assign G793GAT = G717GAT & G782GAT;
  assign G794GAT = G219GAT & G786GAT;
  assign G795GAT = ~G628GAT | ~G773GAT;
  assign G796GAT = ~G795GAT | ~G747GAT;
  assign G802GAT = ~G788GAT & ~G789GAT;
  assign G803GAT = ~G790GAT & ~G791GAT;
  assign G804GAT = ~G792GAT & ~G793GAT;
  assign G805GAT = ~G340GAT & ~G794GAT;
  assign G806GAT = ~G692GAT & ~G796GAT;
  assign G807GAT = G692GAT & G796GAT;
  assign G808GAT = G219GAT & G802GAT;
  assign G809GAT = G219GAT & G803GAT;
  assign G810GAT = G219GAT & G804GAT;
  assign G811GAT = ~G529GAT | ~G731GAT | ~G805GAT | ~G787GAT;
  assign G812GAT = ~G619GAT | ~G796GAT;
  assign G813GAT = ~G796GAT | ~G609GAT | ~G619GAT;
  assign G814GAT = ~G796GAT | ~G619GAT | ~G600GAT | ~G609GAT;
  assign G815GAT = ~G814GAT | ~G766GAT | ~G738GAT | ~G765GAT;
  assign G819GAT = ~G813GAT | ~G741GAT | ~G764GAT;
  assign G822GAT = ~G744GAT | ~G812GAT;
  assign G825GAT = ~G806GAT & ~G807GAT;
  assign G826GAT = ~G335GAT & ~G808GAT;
  assign G827GAT = ~G336GAT & ~G809GAT;
  assign G828GAT = ~G338GAT & ~G810GAT;
  assign G829GAT = ~G811GAT;
  assign G830GAT = ~G665GAT & ~G815GAT;
  assign G831GAT = G665GAT & G815GAT;
  assign G832GAT = ~G673GAT & ~G819GAT;
  assign G833GAT = G673GAT & G819GAT;
  assign G834GAT = ~G682GAT & ~G822GAT;
  assign G835GAT = G682GAT & G822GAT;
  assign G836GAT = G219GAT & G825GAT;
  assign G837GAT = ~G704GAT | ~G826GAT | ~G777GAT;
  assign G838GAT = ~G527GAT | ~G712GAT | ~G827GAT | ~G781GAT;
  assign G839GAT = ~G528GAT | ~G721GAT | ~G828GAT | ~G785GAT;
  assign G840GAT = ~G829GAT;
  assign G841GAT = ~G815GAT | ~G593GAT;
  assign G842GAT = ~G830GAT & ~G831GAT;
  assign G843GAT = ~G832GAT & ~G833GAT;
  assign G844GAT = ~G834GAT & ~G835GAT;
  assign G845GAT = ~G334GAT & ~G836GAT;
  assign G846GAT = ~G837GAT;
  assign G847GAT = ~G838GAT;
  assign G848GAT = ~G839GAT;
  assign G849GAT = G735GAT & G841GAT;
  assign G850GAT = G840GAT;
  assign G851GAT = G219GAT & G842GAT;
  assign G852GAT = G219GAT & G843GAT;
  assign G853GAT = G219GAT & G844GAT;
  assign G854GAT = ~G696GAT | ~G845GAT | ~G772GAT;
  assign G855GAT = ~G846GAT;
  assign G856GAT = ~G847GAT;
  assign G857GAT = ~G848GAT;
  assign G858GAT = ~G849GAT;
  assign G859GAT = ~G417GAT & ~G851GAT;
  assign G860GAT = ~G332GAT & ~G852GAT;
  assign G861GAT = ~G333GAT & ~G853GAT;
  assign G862GAT = ~G854GAT;
  assign G863GAT = G855GAT;
  assign G864GAT = G856GAT;
  assign G865GAT = G857GAT;
  assign G866GAT = G858GAT;
  assign G867GAT = ~G669GAT | ~G859GAT | ~G769GAT;
  assign G868GAT = ~G677GAT | ~G860GAT | ~G770GAT;
  assign G869GAT = ~G686GAT | ~G861GAT | ~G771GAT;
  assign G870GAT = ~G862GAT;
  assign G871GAT = ~G867GAT;
  assign G872GAT = ~G868GAT;
  assign G873GAT = ~G869GAT;
  assign G874GAT = G870GAT;
  assign G875GAT = ~G871GAT;
  assign G876GAT = ~G872GAT;
  assign G877GAT = ~G873GAT;
  assign G878GAT = G875GAT;
  assign G879GAT = G876GAT;
  assign G880GAT = G877GAT;
endmodule


