// Benchmark "c2670" written by ABC on Thu Mar  5 01:06:36 2020

module c2670 ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194,
    G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206,
    G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241,
    G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253,
    G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269,
    G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452, G483,
    G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384,
    G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066,
    G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106,
    G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179,
    G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193,
    G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205,
    G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240,
    G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252,
    G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268,
    G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452,
    G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348,
    G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996,
    G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105,
    G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474,
    G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire G546, G560, G1385, G157, G547, G258, G480, G486, G654, G655, G658,
    G772, G795, G865, G875, G882, G1251, G1254, G1261, G1284, G1344, G1351,
    G1394, G1418, G2433, G2434, G2441, G2442, G2449, G2450, G2478, G1631,
    G1655, G1710, G1721, G2682, G1955, G1959, G1964, G1969, G1974, G1979,
    G1984, G1989, G1994, G1999, G2001, G2012, G2070, G2076, G2082, G2088,
    G2094, G2099, G2103, G2457, G2458, G2461, G2464, G2471, G2479, G2482,
    G2487, G2490, G2495, G2498, G2505, G2508, G2675, G2683, G2686, G2691,
    G2694, G2699, G2702, G487, G1475, G1476, G1484, G1485, G1493, G1494,
    G2459, G2460, G216, G1253, G1256, G558, G748, G784, G807, G821, G825,
    G829, G833, G837, G881, G994, G1273, G1296, G1310, G1314, G1318, G1322,
    G1326, G1406, G1430, G1444, G1448, G1452, G1456, G1460, G1477, G1486,
    G1495, G2477, G1499, G2485, G2486, G2493, G2494, G1643, G1667, G1681,
    G1685, G1689, G1693, G1697, G1716, G1728, G2681, G1776, G2689, G2690,
    G2697, G2698, G1831, G1893, G2007, G2018, G2467, G2468, G2501, G2502,
    G2511, G2512, G2518, G2551, G2559, G2567, G2575, G2583, G2591, G2599,
    G2607, G2615, G2623, G2705, G2706, G2735, G2743, G2751, G2759, G2767,
    G2775, G550, G552, G894, G1498, G1507, G1508, G1516, G1517, G1775,
    G1784, G1785, G1793, G1794, G2469, G2470, G2503, G2504, G2513, G2514,
    G2707, G2708, G551, G553, G818, G819, G820, G822, G823, G824, G826,
    G827, G828, G830, G831, G832, G834, G835, G836, G1307, G1308, G1309,
    G1311, G1312, G1313, G1315, G1316, G1317, G1319, G1320, G1321, G1323,
    G1324, G1325, G1441, G1442, G1443, G1445, G1446, G1447, G1449, G1450,
    G1451, G1453, G1454, G1455, G1457, G1458, G1459, G1481, G1490, G1500,
    G1509, G1518, G1521, G1525, G2557, G2565, G2573, G2581, G2589, G2597,
    G2605, G2613, G2621, G2629, G1678, G1679, G1680, G1682, G1683, G1684,
    G1686, G1687, G1688, G1690, G1691, G1692, G1694, G1695, G1696, G1734,
    G1736, G1738, G1740, G1742, G1744, G1746, G1748, G1750, G1777, G1786,
    G1795, G2023, G2025, G2027, G2029, G2031, G2033, G2035, G2037, G2741,
    G2749, G2757, G2765, G2773, G2781, G2515, G2522, G2525, G2528, G2730,
    G554, G838, G841, G846, G854, G857, G1327, G1329, G1331, G1333, G1335,
    G1461, G1464, G1467, G1470, G1473, G1698, G1701, G1704, G1707, G2634,
    G1504, G1513, G1524, G1528, G1529, G1533, G1538, G1541, G1781, G1790,
    G1806, G1810, G2734, G2521, G2524, G2531, G2532, G144, G147, G152,
    G175, G187, G516, G852, G885, G887, G893, G1028, G1031, G1035, G1041,
    G1049, G1057, G1060, G1066, G1072, G1078, G1213, G1218, G1250, G1387,
    G1389, G1537, G1540, G1735, G1737, G1739, G1741, G1743, G1745, G1747,
    G1749, G1751, G2638, G2024, G2026, G2028, G2030, G2032, G2034, G2036,
    G2038, G2154, G2523, G2533, G2534, G2631, G2639, G2642, G2647, G2650,
    G2655, G2658, G2665, G2668, G1532, G1536, G1539, G1542, G1544, G1547,
    G2065, G1809, G1813, G1821, G1824, G2538, G2546, G2554, G2562, G2570,
    G2578, G2586, G2594, G2602, G2610, G2618, G2626, G2738, G2746, G2754,
    G2762, G2770, G2778, G456, G466, G562, G883, G889, G891, G1043, G1051,
    G1062, G1068, G1074, G1080, G1225, G1227, G1232, G1234, G1543, G1546,
    G2637, G1753, G2645, G2646, G2653, G2654, G1820, G1823, G2107, G2110,
    G2118, G2123, G2151, G2158, G2161, G2164, G2172, G2235, G2262, G2350,
    G2535, G2661, G2662, G2671, G2672, G468, G897, G898, G1228, G1235,
    G1545, G1548, G2542, G2550, G1561, G2558, G1565, G2566, G1569, G2574,
    G1573, G2582, G1577, G2590, G1581, G2598, G1585, G2606, G1589, G2614,
    G1593, G2622, G1597, G2630, G1752, G1761, G1762, G1770, G1771, G1822,
    G1825, G2039, G2742, G2043, G2750, G2047, G2758, G2051, G2766, G2055,
    G2774, G2059, G2782, G2663, G2664, G2673, G2674, G146, G462, G2113,
    G2114, G2122, G2129, G592, G2167, G2168, G2176, G2241, G2266, G743,
    G749, G886, G995, G1006, G1550, G2354, G2541, G1562, G1566, G1570,
    G1574, G1578, G1582, G1586, G1590, G1594, G1598, G1754, G1763, G1772,
    G2040, G2044, G2048, G2052, G2056, G2060, G2115, G2126, G2131, G2134,
    G2141, G2144, G2157, G2160, G2169, G2177, G2180, G2187, G2190, G2207,
    G2254, G2334, G2342, G2422, G2543, G2709, G2712, G2727, G569, G570,
    G599, G600, G896, G1549, G1243, G1245, G1257, G1258, G1563, G1567,
    G1571, G1575, G1579, G1583, G1587, G1591, G1595, G1599, G2041, G2045,
    G2049, G2053, G2057, G2061, G2159, G475, G490, G496, G502, G508, G765,
    G769, G571, G2121, G579, G587, G2130, G596, G601, G2175, G609, G2258,
    G1014, G1018, G717, G723, G729, G735, G753, G2338, G999, G1091, G2346,
    G2426, G1337, G2549, G1552, G1600, G1596, G1592, G1588, G1584, G1580,
    G1576, G1572, G1568, G1564, G2062, G2058, G2054, G2050, G2046, G2042,
    G1758, G1767, G1798, G1802, G2733, G1829, G2137, G2138, G2147, G2148,
    G2183, G2184, G2193, G2194, G2210, G2213, G2715, G2716, G1094, G1096,
    G578, G588, G608, G742, G1005, G1092, G1551, G1554, G1555, G1557,
    G1558, G1828, G1845, G1907, G2139, G2140, G2149, G2150, G2185, G2186,
    G2195, G2196, G2717, G2718, G154, G155, G763, G767, G531, G537, G575,
    G580, G589, G605, G610, G1012, G1016, G705, G711, G1093, G1355, G1553,
    G1556, G1559, G1601, G1801, G1805, G1815, G1818, G1830, G1836, G1850,
    G1898, G1912, G2197, G2200, G2214, G2215, G2217, G2220, G2722, G492,
    G498, G504, G510, G519, G525, G533, G539, G693, G699, G707, G713, G719,
    G725, G731, G737, G1560, G1814, G1817, G2216, G493, G499, G505, G511,
    G521, G527, G534, G540, G584, G613, G617, G621, G625, G676, G695, G701,
    G708, G714, G720, G726, G732, G738, G1087, G1108, G1361, G1369, G1373,
    G1377, G1607, G1615, G1619, G1623, G1816, G1819, G2726, G1842, G1858,
    G1863, G1866, G1868, G1870, G1872, G1874, G1876, G1904, G1920, G1925,
    G1928, G1930, G1932, G1934, G1936, G1938, G2203, G2204, G2223, G2224,
    G2238, G522, G528, G696, G702, G1881, G1883, G1885, G1887, G1889,
    G1891, G1943, G1945, G1947, G1949, G1951, G1953, G2205, G2206, G2225,
    G2226, G2719, G616, G620, G624, G628, G630, G633, G636, G639, G645,
    G2242, G675, G1107, G1368, G1371, G1375, G1614, G1617, G1621, G1856,
    G1861, G1918, G1923, G2230, G2246, G2270, G2278, G2286, G2294, G2302,
    G2310, G2358, G2366, G2374, G2382, G2390, G2398, G629, G632, G635,
    G638, G646, G677, G1827, G907, G915, G922, G924, G937, G946, G1109,
    G1125, G1133, G1140, G1142, G1155, G1164, G1378, G1380, G1382, G1624,
    G1626, G1628, G2725, G1859, G1864, G1921, G1926, G2267, G2275, G2283,
    G2291, G2299, G2307, G2318, G2326, G2355, G2363, G2371, G2379, G2387,
    G2395, G2406, G2414, G647, G631, G634, G637, G640, G2234, G2250, G679,
    G1826, G2274, G2282, G2290, G2298, G2306, G2314, G1110, G2362, G2370,
    G2378, G2386, G2394, G2402, G1877, G1879, G1939, G1941, G143, G671,
    G674, G686, G2273, G900, G2281, G909, G2289, G917, G2297, G926, G2305,
    G929, G2313, G939, G2322, G2330, G967, G1104, G1106, G2361, G1118,
    G2369, G1127, G2377, G1135, G2385, G1144, G2393, G1147, G2401, G1157,
    G2410, G2418, G1184, G2227, G2243, G2251, G2259, G2331, G2339, G2347,
    G2419, G687, G899, G908, G916, G925, G928, G938, G954, G961, G1117,
    G1126, G1134, G1143, G1146, G1156, G1172, G1179, G2315, G2323, G2403,
    G2411, G2233, G642, G2249, G649, G2257, G665, G684, G2265, G688, G901,
    G910, G918, G927, G930, G940, G2337, G963, G2345, G1099, G1115, G2353,
    G1119, G1128, G1136, G1145, G1148, G1158, G2425, G1181, G641, G648,
    G664, G683, G2321, G948, G2329, G956, G962, G1098, G1114, G2409, G1166,
    G2417, G1174, G1180, G643, G650, G666, G681, G690, G947, G955, G964,
    G968, G970, G971, G972, G978, G979, G1100, G1112, G1165, G1173, G1182,
    G1185, G1187, G1188, G1189, G1195, G1196, G644, G884, G949, G957, G969,
    G973, G1167, G1175, G1186, G1190, G680, G682, G895, G1025, G1111,
    G1113, G685, G976, G977, G980, G981, G1116, G1193, G1194, G1197, G1198,
    G982, G983, G988, G1027, G1199, G1200, G1205, G984, G1085, G1201, G987,
    G990, G1204, G1207, G989, G1206, G991, G1208, G1221, G1238, G1239,
    G1240, G1247, G471, G473, G1088, G1089;
  assign G350 = G452;
  assign G335 = G452;
  assign G409 = G452;
  assign G546 = G1 & G3;
  assign G560 = ~G559;
  assign G369 = G1083;
  assign G367 = G1083;
  assign G1385 = ~G1384;
  assign G411 = G2066;
  assign G337 = G2066;
  assign G384 = G2066;
  assign G157 = G2072 & G2078 & G2090 & G2084;
  assign G547 = ~G546;
  assign G218 = ~G44;
  assign G219 = ~G132;
  assign G220 = ~G82;
  assign G221 = ~G96;
  assign G235 = ~G69;
  assign G236 = ~G120;
  assign G237 = ~G57;
  assign G238 = ~G108;
  assign G258 = G661 & G2 & G15;
  assign G480 = G661;
  assign G486 = G37 & G37;
  assign G654 = G452;
  assign G655 = G8;
  assign G658 = G8;
  assign G772 = G543;
  assign G795 = G651;
  assign G865 = ~G860;
  assign G875 = ~G868;
  assign G882 = G11 & G868;
  assign G1251 = G44 & G96 & G132 & G82;
  assign G1254 = G69 & G108 & G120 & G57;
  assign G1261 = G543;
  assign G1284 = G651;
  assign G1344 = ~G1341;
  assign G1351 = ~G1348;
  assign G1394 = G2104;
  assign G1418 = G2105;
  assign G2433 = ~G2427;
  assign G2434 = ~G2430;
  assign G2441 = ~G2435;
  assign G2442 = ~G2438;
  assign G2449 = ~G2443;
  assign G2450 = ~G2446;
  assign G2478 = ~G2474;
  assign G1631 = G2104;
  assign G1655 = G2105;
  assign G1710 = G16;
  assign G1721 = G16;
  assign G2682 = ~G2678;
  assign G1955 = G7 & G661;
  assign G1959 = ~G1956;
  assign G1964 = ~G1961;
  assign G1969 = ~G1966;
  assign G1974 = ~G1971;
  assign G1979 = ~G1976;
  assign G1984 = ~G1981;
  assign G1989 = ~G1986;
  assign G1994 = ~G1991;
  assign G1999 = ~G1996;
  assign G2001 = G29;
  assign G2012 = G29;
  assign G2070 = ~G2067;
  assign G2076 = ~G2072;
  assign G2082 = ~G2078;
  assign G2088 = ~G2084;
  assign G2094 = ~G2090;
  assign G2099 = ~G2096;
  assign G2103 = ~G2100;
  assign G2457 = ~G2451;
  assign G2458 = ~G2454;
  assign G2461 = G1348;
  assign G2464 = G1341;
  assign G2471 = G1956;
  assign G2479 = G1966;
  assign G2482 = G1961;
  assign G2487 = G1976;
  assign G2490 = G1971;
  assign G2495 = G1986;
  assign G2498 = G1981;
  assign G2505 = G1996;
  assign G2508 = G1991;
  assign G2675 = G2067;
  assign G2683 = G2078;
  assign G2686 = G2072;
  assign G2691 = G2090;
  assign G2694 = G2084;
  assign G2699 = G2100;
  assign G2702 = G2096;
  assign G158 = ~G157;
  assign G259 = ~G258;
  assign G487 = ~G486;
  assign G391 = G654;
  assign G1475 = ~G2430 | ~G2433;
  assign G1476 = ~G2427 | ~G2434;
  assign G1484 = ~G2438 | ~G2441;
  assign G1485 = ~G2435 | ~G2442;
  assign G1493 = ~G2446 | ~G2449;
  assign G1494 = ~G2443 | ~G2450;
  assign G2459 = ~G2454 | ~G2457;
  assign G2460 = ~G2451 | ~G2458;
  assign G173 = G94 & G654;
  assign G216 = G2106 & G1955;
  assign G223 = ~G1955;
  assign G234 = ~G567 | ~G1955;
  assign G1253 = ~G1251;
  assign G1256 = ~G1254;
  assign G558 = G1254 & G1251;
  assign G748 = G655;
  assign G784 = ~G772;
  assign G807 = ~G795;
  assign G821 = G795 & G80 & G772;
  assign G825 = G795 & G68 & G772;
  assign G829 = G795 & G79 & G772;
  assign G833 = G795 & G78 & G772;
  assign G837 = G795 & G77 & G772;
  assign G881 = G11 & G875;
  assign G994 = G655;
  assign G1273 = ~G1261;
  assign G1296 = ~G1284;
  assign G1310 = G1284 & G76 & G1261;
  assign G1314 = G1284 & G75 & G1261;
  assign G1318 = G1284 & G74 & G1261;
  assign G1322 = G1284 & G73 & G1261;
  assign G1326 = G1284 & G72 & G1261;
  assign G1406 = ~G1394;
  assign G1430 = ~G1418;
  assign G1444 = G1418 & G114 & G1394;
  assign G1448 = G1418 & G113 & G1394;
  assign G1452 = G1418 & G112 & G1394;
  assign G1456 = G1418 & G111 & G1394;
  assign G1460 = G1394 & G1418;
  assign G1477 = ~G1475 | ~G1476;
  assign G1486 = ~G1484 | ~G1485;
  assign G1495 = ~G1493 | ~G1494;
  assign G2477 = ~G2471;
  assign G1499 = ~G2471 | ~G2478;
  assign G2485 = ~G2479;
  assign G2486 = ~G2482;
  assign G2493 = ~G2487;
  assign G2494 = ~G2490;
  assign G1643 = ~G1631;
  assign G1667 = ~G1655;
  assign G1681 = G1655 & G118 & G1631;
  assign G1685 = G1655 & G107 & G1631;
  assign G1689 = G1655 & G117 & G1631;
  assign G1693 = G1655 & G116 & G1631;
  assign G1697 = G1655 & G115 & G1631;
  assign G1716 = ~G1710;
  assign G1728 = ~G1721;
  assign G2681 = ~G2675;
  assign G1776 = ~G2675 | ~G2682;
  assign G2689 = ~G2683;
  assign G2690 = ~G2686;
  assign G2697 = ~G2691;
  assign G2698 = ~G2694;
  assign G1831 = G658;
  assign G1893 = G658;
  assign G2007 = ~G2001;
  assign G2018 = ~G2012;
  assign G2467 = ~G2461;
  assign G2468 = ~G2464;
  assign G2501 = ~G2495;
  assign G2502 = ~G2498;
  assign G2511 = ~G2505;
  assign G2512 = ~G2508;
  assign G2518 = ~G2459 | ~G2460;
  assign G2551 = G1344;
  assign G2559 = G1351;
  assign G2567 = G1959;
  assign G2575 = G1964;
  assign G2583 = G1969;
  assign G2591 = G1974;
  assign G2599 = G1979;
  assign G2607 = G1984;
  assign G2615 = G1989;
  assign G2623 = G1994;
  assign G2705 = ~G2699;
  assign G2706 = ~G2702;
  assign G2735 = G1999;
  assign G2743 = G2070;
  assign G2751 = G2076;
  assign G2759 = G2082;
  assign G2767 = G2088;
  assign G2775 = G2094;
  assign G217 = ~G216;
  assign G550 = G2106 & G1253;
  assign G552 = G567 & G1256;
  assign G325 = G558;
  assign G894 = G881 | G882;
  assign G1498 = ~G2474 | ~G2477;
  assign G1507 = ~G2482 | ~G2485;
  assign G1508 = ~G2479 | ~G2486;
  assign G1516 = ~G2490 | ~G2493;
  assign G1517 = ~G2487 | ~G2494;
  assign G1775 = ~G2678 | ~G2681;
  assign G1784 = ~G2686 | ~G2689;
  assign G1785 = ~G2683 | ~G2690;
  assign G1793 = ~G2694 | ~G2697;
  assign G1794 = ~G2691 | ~G2698;
  assign G2469 = ~G2464 | ~G2467;
  assign G2470 = ~G2461 | ~G2468;
  assign G2503 = ~G2498 | ~G2501;
  assign G2504 = ~G2495 | ~G2502;
  assign G2513 = ~G2508 | ~G2511;
  assign G2514 = ~G2505 | ~G2512;
  assign G2707 = ~G2702 | ~G2705;
  assign G2708 = ~G2699 | ~G2706;
  assign G261 = ~G558;
  assign G551 = ~G550;
  assign G553 = ~G552;
  assign G818 = G807 & G93 & G784;
  assign G819 = G807 & G55 & G772;
  assign G820 = G795 & G67 & G784;
  assign G822 = G807 & G81 & G784;
  assign G823 = G807 & G43 & G772;
  assign G824 = G795 & G56 & G784;
  assign G826 = G807 & G92 & G784;
  assign G827 = G807 & G54 & G772;
  assign G828 = G795 & G66 & G784;
  assign G830 = G807 & G91 & G784;
  assign G831 = G807 & G53 & G772;
  assign G832 = G795 & G65 & G784;
  assign G834 = G807 & G90 & G784;
  assign G835 = G807 & G52 & G772;
  assign G836 = G795 & G64 & G784;
  assign G1307 = G1296 & G89 & G1273;
  assign G1308 = G1296 & G51 & G1261;
  assign G1309 = G1284 & G63 & G1273;
  assign G1311 = G1296 & G88 & G1273;
  assign G1312 = G1296 & G50 & G1261;
  assign G1313 = G1284 & G62 & G1273;
  assign G1315 = G1296 & G87 & G1273;
  assign G1316 = G1296 & G49 & G1261;
  assign G1317 = G1273 & G1284;
  assign G1319 = G1296 & G86 & G1273;
  assign G1320 = G1296 & G48 & G1261;
  assign G1321 = G1284 & G61 & G1273;
  assign G1323 = G1296 & G85 & G1273;
  assign G1324 = G1296 & G47 & G1261;
  assign G1325 = G1284 & G60 & G1273;
  assign G1441 = G1430 & G138 & G1406;
  assign G1442 = G1430 & G102 & G1394;
  assign G1443 = G1418 & G126 & G1406;
  assign G1445 = G1430 & G137 & G1406;
  assign G1446 = G1430 & G101 & G1394;
  assign G1447 = G1418 & G125 & G1406;
  assign G1449 = G1430 & G136 & G1406;
  assign G1450 = G1430 & G100 & G1394;
  assign G1451 = G1418 & G124 & G1406;
  assign G1453 = G1430 & G135 & G1406;
  assign G1454 = G1430 & G99 & G1394;
  assign G1455 = G1418 & G123 & G1406;
  assign G1457 = G1406 & G1430;
  assign G1458 = G1394 & G1430;
  assign G1459 = G1406 & G1418;
  assign G1481 = ~G1477;
  assign G1490 = ~G1486;
  assign G1500 = ~G1498 | ~G1499;
  assign G1509 = ~G1507 | ~G1508;
  assign G1518 = ~G1516 | ~G1517;
  assign G1521 = G1495;
  assign G1525 = G1495;
  assign G2557 = ~G2551;
  assign G2565 = ~G2559;
  assign G2573 = ~G2567;
  assign G2581 = ~G2575;
  assign G2589 = ~G2583;
  assign G2597 = ~G2591;
  assign G2605 = ~G2599;
  assign G2613 = ~G2607;
  assign G2621 = ~G2615;
  assign G2629 = ~G2623;
  assign G1678 = G1667 & G142 & G1643;
  assign G1679 = G1667 & G106 & G1631;
  assign G1680 = G1655 & G130 & G1643;
  assign G1682 = G1667 & G131 & G1643;
  assign G1683 = G1667 & G95 & G1631;
  assign G1684 = G1655 & G119 & G1643;
  assign G1686 = G1667 & G141 & G1643;
  assign G1687 = G1667 & G105 & G1631;
  assign G1688 = G1655 & G129 & G1643;
  assign G1690 = G1667 & G140 & G1643;
  assign G1691 = G1667 & G104 & G1631;
  assign G1692 = G1655 & G128 & G1643;
  assign G1694 = G1667 & G139 & G1643;
  assign G1695 = G1667 & G103 & G1631;
  assign G1696 = G1655 & G127 & G1643;
  assign G1734 = G19 & G1716;
  assign G1736 = G4 & G1716;
  assign G1738 = G20 & G1716;
  assign G1740 = G5 & G1716;
  assign G1742 = G21 & G1728;
  assign G1744 = G22 & G1728;
  assign G1746 = G23 & G1728;
  assign G1748 = G6 & G1728;
  assign G1750 = G24 & G1728;
  assign G1777 = ~G1775 | ~G1776;
  assign G1786 = ~G1784 | ~G1785;
  assign G1795 = ~G1793 | ~G1794;
  assign G2023 = G25 & G2007;
  assign G2025 = G32 & G2007;
  assign G2027 = G26 & G2007;
  assign G2029 = G33 & G2007;
  assign G2031 = G27 & G2018;
  assign G2033 = G34 & G2018;
  assign G2035 = G35 & G2018;
  assign G2037 = G28 & G2018;
  assign G2741 = ~G2735;
  assign G2749 = ~G2743;
  assign G2757 = ~G2751;
  assign G2765 = ~G2759;
  assign G2773 = ~G2767;
  assign G2781 = ~G2775;
  assign G2515 = ~G2469 | ~G2470;
  assign G2522 = ~G2518;
  assign G2525 = ~G2513 | ~G2514;
  assign G2528 = ~G2503 | ~G2504;
  assign G2730 = ~G2707 | ~G2708;
  assign G554 = G551 & G553;
  assign G838 = G821 | G820 | G818 | G819;
  assign G841 = G825 | G824 | G822 | G823;
  assign G846 = G829 | G828 | G826 | G827;
  assign G854 = G833 | G832 | G830 | G831;
  assign G857 = G837 | G836 | G834 | G835;
  assign G1327 = G1310 | G1309 | G1307 | G1308;
  assign G1329 = G1314 | G1313 | G1311 | G1312;
  assign G1331 = G1318 | G1317 | G1315 | G1316;
  assign G1333 = G1322 | G1321 | G1319 | G1320;
  assign G1335 = G1326 | G1325 | G1323 | G1324;
  assign G1461 = G1444 | G1443 | G1441 | G1442;
  assign G1464 = G1448 | G1447 | G1445 | G1446;
  assign G1467 = G1452 | G1451 | G1449 | G1450;
  assign G1470 = G1456 | G1455 | G1453 | G1454;
  assign G1473 = G1460 | G1459 | G1457 | G1458;
  assign G1698 = G1685 | G1684 | G1682 | G1683;
  assign G1701 = G1689 | G1688 | G1686 | G1687;
  assign G1704 = G1693 | G1692 | G1690 | G1691;
  assign G1707 = G1697 | G1696 | G1694 | G1695;
  assign G2634 = G1681 | G1680 | G1678 | G1679;
  assign G319 = G554;
  assign G1504 = ~G1500;
  assign G1513 = ~G1509;
  assign G1524 = ~G1521;
  assign G1528 = ~G1525;
  assign G1529 = G1518;
  assign G1533 = G1518;
  assign G1538 = G1521 & G1486 & G1477;
  assign G1541 = G1525 & G1490 & G1481;
  assign G1781 = ~G1777;
  assign G1790 = ~G1786;
  assign G1806 = G1795;
  assign G1810 = G1795;
  assign G2734 = ~G2730;
  assign G2521 = ~G2515;
  assign G2524 = ~G2515 | ~G2522;
  assign G2531 = ~G2525;
  assign G2532 = ~G2528;
  assign G144 = G838 & G860;
  assign G147 = G846 & G860;
  assign G152 = G841 & G860;
  assign G160 = ~G1464;
  assign G162 = ~G1467;
  assign G164 = ~G1461;
  assign G166 = ~G1329;
  assign G168 = ~G1327;
  assign G171 = ~G857;
  assign G175 = G554 & G36 & G480 & G483;
  assign G187 = G547 & G554 & G480 & G483;
  assign G516 = G838;
  assign G852 = ~G846;
  assign G885 = G841 & G875;
  assign G887 = G846 & G875;
  assign G893 = G1327 & G868;
  assign G1028 = ~G838;
  assign G1031 = ~G841;
  assign G1035 = ~G846;
  assign G1041 = G854;
  assign G1049 = G857;
  assign G1057 = G1327;
  assign G1060 = G1329;
  assign G1066 = G1331;
  assign G1072 = G1333;
  assign G1078 = G1335;
  assign G1213 = ~G2099 | ~G1470;
  assign G1218 = ~G2103 | ~G1473;
  assign G1250 = G1704;
  assign G1387 = G1461 & G1385;
  assign G1389 = ~G1464;
  assign G1537 = G1524 & G1481 & G1486;
  assign G1540 = G1528 & G1477 & G1490;
  assign G1735 = G841 & G1710;
  assign G1737 = G846 & G1710;
  assign G1739 = G854 & G1710;
  assign G1741 = G857 & G1710;
  assign G1743 = G1327 & G1721;
  assign G1745 = G1329 & G1721;
  assign G1747 = G1331 & G1721;
  assign G1749 = G1333 & G1721;
  assign G1751 = G1335 & G1721;
  assign G2638 = ~G2634;
  assign G2024 = G1698 & G2001;
  assign G2026 = G1701 & G2001;
  assign G2028 = G1704 & G2001;
  assign G2030 = G1707 & G2001;
  assign G2032 = G1461 & G2012;
  assign G2034 = G1464 & G2012;
  assign G2036 = G1467 & G2012;
  assign G2038 = G1470 & G2012;
  assign G2154 = G841;
  assign G2523 = ~G2518 | ~G2521;
  assign G2533 = ~G2528 | ~G2531;
  assign G2534 = ~G2525 | ~G2532;
  assign G2631 = G1698;
  assign G2639 = G1704;
  assign G2642 = G1701;
  assign G2647 = G1461;
  assign G2650 = G1707;
  assign G2655 = G1467;
  assign G2658 = G1464;
  assign G2665 = G1473;
  assign G2668 = G1470;
  assign G153 = G865 | G152;
  assign G176 = ~G175;
  assign G188 = ~G187;
  assign G299 = G1041;
  assign G301 = G1049;
  assign G286 = G1057;
  assign G303 = G1060;
  assign G288 = G1066;
  assign G305 = G1072;
  assign G290 = G1078;
  assign G1532 = ~G1529;
  assign G1536 = ~G1533;
  assign G1539 = ~G1537 & ~G1538;
  assign G1542 = ~G1540 & ~G1541;
  assign G1544 = G1529 & G1509 & G1500;
  assign G1547 = G1533 & G1513 & G1504;
  assign G2065 = G2037 | G2038;
  assign G1809 = ~G1806;
  assign G1813 = ~G1810;
  assign G1821 = G1806 & G1786 & G1777;
  assign G1824 = G1810 & G1790 & G1781;
  assign G2538 = ~G2523 | ~G2524;
  assign G2546 = ~G2533 | ~G2534;
  assign G2554 = G1734 | G1735;
  assign G2562 = G1736 | G1737;
  assign G2570 = G1738 | G1739;
  assign G2578 = G1740 | G1741;
  assign G2586 = G1742 | G1743;
  assign G2594 = G1744 | G1745;
  assign G2602 = G1746 | G1747;
  assign G2610 = G1748 | G1749;
  assign G2618 = G1750 | G1751;
  assign G2626 = G2023 | G2024;
  assign G2738 = G2025 | G2026;
  assign G2746 = G2027 | G2028;
  assign G2754 = G2029 | G2030;
  assign G2762 = G2031 | G2032;
  assign G2770 = G2033 | G2034;
  assign G2778 = G2035 | G2036;
  assign G456 = G40 & G1389 & G1387;
  assign G466 = ~G1387;
  assign G562 = ~G560 | ~G852;
  assign G883 = G516 & G875;
  assign G889 = G1049 & G868;
  assign G891 = G1041 & G875;
  assign G1043 = ~G1041;
  assign G1051 = ~G1049;
  assign G1062 = ~G1060;
  assign G1068 = ~G1066;
  assign G1074 = ~G1072;
  assign G1080 = ~G1078;
  assign G1225 = G2099 & G1213;
  assign G1227 = G1213 & G1470;
  assign G1232 = G2103 & G1218;
  assign G1234 = G1218 & G1473;
  assign G1543 = G1532 & G1504 & G1509;
  assign G1546 = G1536 & G1500 & G1513;
  assign G2637 = ~G2631;
  assign G1753 = ~G2631 | ~G2638;
  assign G2645 = ~G2639;
  assign G2646 = ~G2642;
  assign G2653 = ~G2647;
  assign G2654 = ~G2650;
  assign G1820 = G1809 & G1781 & G1786;
  assign G1823 = G1813 & G1777 & G1790;
  assign G2107 = G1031;
  assign G2110 = G1028;
  assign G2118 = G1035;
  assign G2123 = ~G1057;
  assign G2151 = ~G852;
  assign G2158 = ~G2154;
  assign G2161 = G1031;
  assign G2164 = G1028;
  assign G2172 = G1035;
  assign G2235 = G516;
  assign G2262 = G1035;
  assign G2350 = G1035;
  assign G2535 = ~G1542 | ~G1539;
  assign G2661 = ~G2655;
  assign G2662 = ~G2658;
  assign G2671 = ~G2665;
  assign G2672 = ~G2668;
  assign G468 = G466 & G40 & G1389;
  assign G897 = G887 | G889;
  assign G898 = G891 | G893;
  assign G1228 = G1225 | G1227;
  assign G1235 = G1232 | G1234;
  assign G1545 = ~G1543 & ~G1544;
  assign G1548 = ~G1546 & ~G1547;
  assign G2542 = ~G2538;
  assign G2550 = ~G2546;
  assign G1561 = ~G2554 | ~G2557;
  assign G2558 = ~G2554;
  assign G1565 = ~G2562 | ~G2565;
  assign G2566 = ~G2562;
  assign G1569 = ~G2570 | ~G2573;
  assign G2574 = ~G2570;
  assign G1573 = ~G2578 | ~G2581;
  assign G2582 = ~G2578;
  assign G1577 = ~G2586 | ~G2589;
  assign G2590 = ~G2586;
  assign G1581 = ~G2594 | ~G2597;
  assign G2598 = ~G2594;
  assign G1585 = ~G2602 | ~G2605;
  assign G2606 = ~G2602;
  assign G1589 = ~G2610 | ~G2613;
  assign G2614 = ~G2610;
  assign G1593 = ~G2618 | ~G2621;
  assign G2622 = ~G2618;
  assign G1597 = ~G2626 | ~G2629;
  assign G2630 = ~G2626;
  assign G1752 = ~G2634 | ~G2637;
  assign G1761 = ~G2642 | ~G2645;
  assign G1762 = ~G2639 | ~G2646;
  assign G1770 = ~G2650 | ~G2653;
  assign G1771 = ~G2647 | ~G2654;
  assign G1822 = ~G1820 & ~G1821;
  assign G1825 = ~G1823 & ~G1824;
  assign G2039 = ~G2738 | ~G2741;
  assign G2742 = ~G2738;
  assign G2043 = ~G2746 | ~G2749;
  assign G2750 = ~G2746;
  assign G2047 = ~G2754 | ~G2757;
  assign G2758 = ~G2754;
  assign G2051 = ~G2762 | ~G2765;
  assign G2766 = ~G2762;
  assign G2055 = ~G2770 | ~G2773;
  assign G2774 = ~G2770;
  assign G2059 = ~G2778 | ~G2781;
  assign G2782 = ~G2778;
  assign G2663 = ~G2658 | ~G2661;
  assign G2664 = ~G2655 | ~G2662;
  assign G2673 = ~G2668 | ~G2671;
  assign G2674 = ~G2665 | ~G2672;
  assign G146 = G562 & G865;
  assign G462 = ~G456;
  assign G2113 = ~G2107;
  assign G2114 = ~G2110;
  assign G2122 = ~G2118;
  assign G2129 = ~G2123;
  assign G592 = G562;
  assign G2167 = ~G2161;
  assign G2168 = ~G2164;
  assign G2176 = ~G2172;
  assign G2241 = ~G2235;
  assign G2266 = ~G2262;
  assign G743 = ~G456;
  assign G749 = G456;
  assign G886 = G562 & G868;
  assign G284 = G897;
  assign G321 = G897;
  assign G297 = G898;
  assign G280 = G898;
  assign G995 = G456;
  assign G1006 = ~G456;
  assign G1550 = ~G2535 | ~G2542;
  assign G2354 = ~G2350;
  assign G2541 = ~G2535;
  assign G1562 = ~G2551 | ~G2558;
  assign G1566 = ~G2559 | ~G2566;
  assign G1570 = ~G2567 | ~G2574;
  assign G1574 = ~G2575 | ~G2582;
  assign G1578 = ~G2583 | ~G2590;
  assign G1582 = ~G2591 | ~G2598;
  assign G1586 = ~G2599 | ~G2606;
  assign G1590 = ~G2607 | ~G2614;
  assign G1594 = ~G2615 | ~G2622;
  assign G1598 = ~G2623 | ~G2630;
  assign G1754 = ~G1752 | ~G1753;
  assign G1763 = ~G1761 | ~G1762;
  assign G1772 = ~G1770 | ~G1771;
  assign G2040 = ~G2735 | ~G2742;
  assign G2044 = ~G2743 | ~G2750;
  assign G2048 = ~G2751 | ~G2758;
  assign G2052 = ~G2759 | ~G2766;
  assign G2056 = ~G2767 | ~G2774;
  assign G2060 = ~G2775 | ~G2782;
  assign G2115 = G1043;
  assign G2126 = G1051;
  assign G2131 = G1068;
  assign G2134 = G1062;
  assign G2141 = G1080;
  assign G2144 = G1074;
  assign G2157 = ~G2151;
  assign G2160 = ~G2151 | ~G2158;
  assign G2169 = G1043;
  assign G2177 = G1068;
  assign G2180 = G1062;
  assign G2187 = G1080;
  assign G2190 = G1074;
  assign G2207 = ~G562;
  assign G2254 = G1043;
  assign G2334 = G1051;
  assign G2342 = G1043;
  assign G2422 = G1051;
  assign G2543 = ~G1548 | ~G1545;
  assign G2709 = ~G2673 | ~G2674;
  assign G2712 = ~G2663 | ~G2664;
  assign G2727 = ~G1825 | ~G1822;
  assign G148 = G146 | G147;
  assign G569 = ~G2110 | ~G2113;
  assign G570 = ~G2107 | ~G2114;
  assign G599 = ~G2164 | ~G2167;
  assign G600 = ~G2161 | ~G2168;
  assign G896 = G885 | G886;
  assign G1549 = ~G2538 | ~G2541;
  assign G1243 = ~G1228;
  assign G1245 = ~G1235;
  assign G1257 = G468;
  assign G1258 = G468;
  assign G1563 = ~G1561 | ~G1562;
  assign G1567 = ~G1565 | ~G1566;
  assign G1571 = ~G1569 | ~G1570;
  assign G1575 = ~G1573 | ~G1574;
  assign G1579 = ~G1577 | ~G1578;
  assign G1583 = ~G1581 | ~G1582;
  assign G1587 = ~G1585 | ~G1586;
  assign G1591 = ~G1589 | ~G1590;
  assign G1595 = ~G1593 | ~G1594;
  assign G1599 = ~G1597 | ~G1598;
  assign G2041 = ~G2039 | ~G2040;
  assign G2045 = ~G2043 | ~G2044;
  assign G2049 = ~G2047 | ~G2048;
  assign G2053 = ~G2051 | ~G2052;
  assign G2057 = ~G2055 | ~G2056;
  assign G2061 = ~G2059 | ~G2060;
  assign G2159 = ~G2154 | ~G2157;
  assign G475 = G462;
  assign G490 = G1078 & G743;
  assign G496 = G1698 & G743;
  assign G502 = G1701 & G743;
  assign G508 = G1250 & G743;
  assign G765 = G1057 & G749;
  assign G769 = G1060 & G749;
  assign G571 = ~G569 | ~G570;
  assign G2121 = ~G2115;
  assign G579 = ~G2115 | ~G2122;
  assign G587 = ~G2126 | ~G2129;
  assign G2130 = ~G2126;
  assign G596 = ~G592;
  assign G601 = ~G599 | ~G600;
  assign G2175 = ~G2169;
  assign G609 = ~G2169 | ~G2176;
  assign G2258 = ~G2254;
  assign G1014 = G1057 & G995;
  assign G1018 = G1060 & G995;
  assign G717 = G1078 & G1006;
  assign G723 = G1698 & G1006;
  assign G729 = G1701 & G1006;
  assign G735 = G1250 & G1006;
  assign G753 = ~G749;
  assign G282 = G896;
  assign G323 = G896;
  assign G2338 = ~G2334;
  assign G999 = ~G995;
  assign G1091 = ~G1549 | ~G1550;
  assign G2346 = ~G2342;
  assign G2426 = ~G2422;
  assign G1337 = G462;
  assign G2549 = ~G2543;
  assign G1552 = ~G2543 | ~G2550;
  assign G1600 = ~G1599;
  assign G1596 = ~G1595;
  assign G1592 = ~G1591;
  assign G1588 = ~G1587;
  assign G1584 = ~G1583;
  assign G1580 = ~G1579;
  assign G1576 = ~G1575;
  assign G1572 = ~G1571;
  assign G1568 = ~G1567;
  assign G1564 = ~G1563;
  assign G2062 = ~G2061;
  assign G2058 = ~G2057;
  assign G2054 = ~G2053;
  assign G2050 = ~G2049;
  assign G2046 = ~G2045;
  assign G2042 = ~G2041;
  assign G1758 = ~G1754;
  assign G1767 = ~G1763;
  assign G1798 = G1772;
  assign G1802 = G1772;
  assign G2733 = ~G2727;
  assign G1829 = ~G2727 | ~G2734;
  assign G2137 = ~G2131;
  assign G2138 = ~G2134;
  assign G2147 = ~G2141;
  assign G2148 = ~G2144;
  assign G2183 = ~G2177;
  assign G2184 = ~G2180;
  assign G2193 = ~G2187;
  assign G2194 = ~G2190;
  assign G2210 = ~G2159 | ~G2160;
  assign G2213 = ~G2207;
  assign G2715 = ~G2709;
  assign G2716 = ~G2712;
  assign G1094 = G1235 & G1245;
  assign G1096 = G1228 & G1243;
  assign G578 = ~G2118 | ~G2121;
  assign G588 = ~G2123 | ~G2130;
  assign G608 = ~G2172 | ~G2175;
  assign G742 = G1257;
  assign G1005 = G1257;
  assign G1092 = ~G1091;
  assign G1551 = ~G2546 | ~G2549;
  assign G1554 = G1584 & G1588 & G1592 & G1600 & G1596;
  assign G1555 = G1564 & G1568 & G1572 & G1580 & G1576;
  assign G1557 = G2065 & G2062;
  assign G1558 = G2042 & G2046 & G2050 & G2058 & G2054;
  assign G1828 = ~G2730 | ~G2733;
  assign G1845 = G1258;
  assign G1907 = G1258;
  assign G2139 = ~G2134 | ~G2137;
  assign G2140 = ~G2131 | ~G2138;
  assign G2149 = ~G2144 | ~G2147;
  assign G2150 = ~G2141 | ~G2148;
  assign G2185 = ~G2180 | ~G2183;
  assign G2186 = ~G2177 | ~G2184;
  assign G2195 = ~G2190 | ~G2193;
  assign G2196 = ~G2187 | ~G2194;
  assign G2717 = ~G2712 | ~G2715;
  assign G2718 = ~G2709 | ~G2716;
  assign G154 = G1094 | G1245;
  assign G155 = G1096 | G1243;
  assign G763 = G1057 & G753;
  assign G767 = G1060 & G753;
  assign G531 = G1066 & G753;
  assign G537 = G1072 & G753;
  assign G575 = ~G571;
  assign G580 = ~G578 | ~G579;
  assign G589 = ~G587 | ~G588;
  assign G605 = ~G601;
  assign G610 = ~G608 | ~G609;
  assign G1012 = G1057 & G999;
  assign G1016 = G1060 & G999;
  assign G705 = G1066 & G999;
  assign G711 = G1072 & G999;
  assign G1093 = G1092 & G14;
  assign G1355 = G475;
  assign G1553 = ~G1551 | ~G1552;
  assign G1556 = G1554 & G1555;
  assign G1559 = G1557 & G1558;
  assign G1601 = G1337;
  assign G1801 = ~G1798;
  assign G1805 = ~G1802;
  assign G1815 = G1798 & G1763 & G1754;
  assign G1818 = G1802 & G1767 & G1758;
  assign G1830 = ~G1828 | ~G1829;
  assign G1836 = G475;
  assign G1850 = G475;
  assign G1898 = G1337;
  assign G1912 = G1337;
  assign G2197 = ~G2149 | ~G2150;
  assign G2200 = ~G2139 | ~G2140;
  assign G2214 = ~G2210;
  assign G2215 = ~G2210 | ~G2213;
  assign G2217 = ~G2195 | ~G2196;
  assign G2220 = ~G2185 | ~G2186;
  assign G2722 = ~G2717 | ~G2718;
  assign G156 = ~G154 | ~G155;
  assign G492 = G490 & G742;
  assign G498 = G496 & G742;
  assign G504 = G502 & G742;
  assign G510 = G508 & G742;
  assign G519 = G763 | G765;
  assign G525 = G767 | G769;
  assign G533 = G531 & G748;
  assign G539 = G537 & G748;
  assign G693 = G1012 | G1014;
  assign G699 = G1016 | G1018;
  assign G707 = G705 & G994;
  assign G713 = G711 & G994;
  assign G719 = G717 & G1005;
  assign G725 = G723 & G1005;
  assign G731 = G729 & G1005;
  assign G737 = G735 & G1005;
  assign G401 = G1093;
  assign G1560 = G894 & G1556 & G1559;
  assign G1814 = G1801 & G1758 & G1763;
  assign G1817 = G1805 & G1754 & G1767;
  assign G2216 = ~G2207 | ~G2214;
  assign G227 = ~G1830;
  assign G229 = ~G1553;
  assign G493 = ~G492;
  assign G499 = ~G498;
  assign G505 = ~G504;
  assign G511 = ~G510;
  assign G521 = G519 & G748;
  assign G527 = G525 & G748;
  assign G534 = ~G533;
  assign G540 = ~G539;
  assign G584 = ~G580;
  assign G613 = G589;
  assign G617 = G589;
  assign G621 = G610;
  assign G625 = G610;
  assign G676 = G1344 & G1355;
  assign G695 = G693 & G994;
  assign G701 = G699 & G994;
  assign G708 = ~G707;
  assign G714 = ~G713;
  assign G720 = ~G719;
  assign G726 = ~G725;
  assign G732 = ~G731;
  assign G738 = ~G737;
  assign G1087 = ~G1093;
  assign G1108 = G1344 & G1601;
  assign G1361 = ~G1355;
  assign G1369 = G1351 & G1355;
  assign G1373 = G1959 & G1355;
  assign G1377 = G1964 & G1355;
  assign G311 = G1560;
  assign G1607 = ~G1601;
  assign G1615 = G1351 & G1601;
  assign G1619 = G1959 & G1601;
  assign G1623 = G1964 & G1601;
  assign G1816 = ~G1814 & ~G1815;
  assign G1819 = ~G1817 & ~G1818;
  assign G2726 = ~G2722;
  assign G1842 = ~G1836;
  assign G1858 = G1969 & G1836;
  assign G1863 = G1974 & G1836;
  assign G1866 = G1979 & G1836;
  assign G1868 = G1984 & G1836;
  assign G1870 = G1989 & G1850;
  assign G1872 = G1994 & G1850;
  assign G1874 = G1999 & G1850;
  assign G1876 = G2070 & G1850;
  assign G1904 = ~G1898;
  assign G1920 = G1969 & G1898;
  assign G1925 = G1974 & G1898;
  assign G1928 = G1979 & G1898;
  assign G1930 = G1984 & G1898;
  assign G1932 = G1989 & G1912;
  assign G1934 = G1994 & G1912;
  assign G1936 = G1999 & G1912;
  assign G1938 = G2070 & G1912;
  assign G2203 = ~G2197;
  assign G2204 = ~G2200;
  assign G2223 = ~G2217;
  assign G2224 = ~G2220;
  assign G2238 = ~G2215 | ~G2216;
  assign G150 = ~G1560;
  assign G522 = ~G521;
  assign G528 = ~G527;
  assign G696 = ~G695;
  assign G702 = ~G701;
  assign G1881 = G1866 & G1831;
  assign G1883 = G1868 & G1831;
  assign G1885 = G1870 & G1845;
  assign G1887 = G1872 & G1845;
  assign G1889 = G1874 & G1845;
  assign G1891 = G1876 & G1845;
  assign G1943 = G1928 & G1893;
  assign G1945 = G1930 & G1893;
  assign G1947 = G1932 & G1907;
  assign G1949 = G1934 & G1907;
  assign G1951 = G1936 & G1907;
  assign G1953 = G1938 & G1907;
  assign G2205 = ~G2200 | ~G2203;
  assign G2206 = ~G2197 | ~G2204;
  assign G2225 = ~G2220 | ~G2223;
  assign G2226 = ~G2217 | ~G2224;
  assign G2719 = ~G1819 | ~G1816;
  assign G616 = ~G613;
  assign G620 = ~G617;
  assign G624 = ~G621;
  assign G628 = ~G625;
  assign G630 = G613 & G580 & G571;
  assign G633 = G617 & G584 & G575;
  assign G636 = G621 & G601 & G592;
  assign G639 = G625 & G605 & G596;
  assign G645 = ~G2238 | ~G2241;
  assign G2242 = ~G2238;
  assign G675 = G1999 & G1361;
  assign G1107 = G1999 & G1607;
  assign G1368 = G2070 & G1361;
  assign G1371 = G2076 & G1361;
  assign G1375 = G2082 & G1361;
  assign G1614 = G2070 & G1607;
  assign G1617 = G2076 & G1607;
  assign G1621 = G2082 & G1607;
  assign G1856 = G2088 & G1842;
  assign G1861 = G2094 & G1842;
  assign G1918 = G2088 & G1904;
  assign G1923 = G2094 & G1904;
  assign G2230 = ~G2205 | ~G2206;
  assign G2246 = ~G2225 | ~G2226;
  assign G2270 = G511;
  assign G2278 = G505;
  assign G2286 = G499;
  assign G2294 = G493;
  assign G2302 = G540;
  assign G2310 = G534;
  assign G2358 = G738;
  assign G2366 = G732;
  assign G2374 = G726;
  assign G2382 = G720;
  assign G2390 = G714;
  assign G2398 = G708;
  assign G629 = G616 & G575 & G580;
  assign G632 = G620 & G571 & G584;
  assign G635 = G624 & G596 & G601;
  assign G638 = G628 & G592 & G605;
  assign G646 = ~G2235 | ~G2242;
  assign G677 = G675 | G676;
  assign G1827 = ~G2719 | ~G2726;
  assign G907 = G1891 & G511;
  assign G915 = G1889 & G505;
  assign G922 = G1887 & G499;
  assign G924 = G493 & G1885;
  assign G937 = G1883 & G540;
  assign G946 = G1881 & G534;
  assign G1109 = G1107 | G1108;
  assign G1125 = G1953 & G738;
  assign G1133 = G1951 & G732;
  assign G1140 = G1949 & G726;
  assign G1142 = G720 & G1947;
  assign G1155 = G1945 & G714;
  assign G1164 = G1943 & G708;
  assign G1378 = G1368 | G1369;
  assign G1380 = G1371 | G1373;
  assign G1382 = G1375 | G1377;
  assign G1624 = G1614 | G1615;
  assign G1626 = G1617 | G1619;
  assign G1628 = G1621 | G1623;
  assign G2725 = ~G2719;
  assign G1859 = G1856 | G1858;
  assign G1864 = G1861 | G1863;
  assign G1921 = G1918 | G1920;
  assign G1926 = G1923 | G1925;
  assign G2267 = G1891;
  assign G2275 = G1889;
  assign G2283 = G1887;
  assign G2291 = G1885;
  assign G2299 = G1883;
  assign G2307 = G1881;
  assign G2318 = G528;
  assign G2326 = G522;
  assign G2355 = G1953;
  assign G2363 = G1951;
  assign G2371 = G1949;
  assign G2379 = G1947;
  assign G2387 = G1945;
  assign G2395 = G1943;
  assign G2406 = G702;
  assign G2414 = G696;
  assign G647 = ~G645 | ~G646;
  assign G631 = ~G629 & ~G630;
  assign G634 = ~G632 & ~G633;
  assign G637 = ~G635 & ~G636;
  assign G640 = ~G638 & ~G639;
  assign G2234 = ~G2230;
  assign G2250 = ~G2246;
  assign G679 = G677 & G1031;
  assign G1826 = ~G2722 | ~G2725;
  assign G2274 = ~G2270;
  assign G2282 = ~G2278;
  assign G2290 = ~G2286;
  assign G2298 = ~G2294;
  assign G2306 = ~G2302;
  assign G2314 = ~G2310;
  assign G1110 = G1109 & G1031;
  assign G2362 = ~G2358;
  assign G2370 = ~G2366;
  assign G2378 = ~G2374;
  assign G2386 = ~G2382;
  assign G2394 = ~G2390;
  assign G2402 = ~G2398;
  assign G1877 = G1859 & G1831;
  assign G1879 = G1864 & G1831;
  assign G1939 = G1921 & G1893;
  assign G1941 = G1926 & G1893;
  assign G143 = G647 & G865;
  assign G671 = G1380 & G1043;
  assign G674 = G1378 & G1035;
  assign G686 = ~G1826 | ~G1827;
  assign G2273 = ~G2267;
  assign G900 = ~G2267 | ~G2274;
  assign G2281 = ~G2275;
  assign G909 = ~G2275 | ~G2282;
  assign G2289 = ~G2283;
  assign G917 = ~G2283 | ~G2290;
  assign G2297 = ~G2291;
  assign G926 = ~G2291 | ~G2298;
  assign G2305 = ~G2299;
  assign G929 = ~G2299 | ~G2306;
  assign G2313 = ~G2307;
  assign G939 = ~G2307 | ~G2314;
  assign G2322 = ~G2318;
  assign G2330 = ~G2326;
  assign G967 = G1382 & G1051;
  assign G1104 = G1626 & G1043;
  assign G1106 = G1624 & G1035;
  assign G2361 = ~G2355;
  assign G1118 = ~G2355 | ~G2362;
  assign G2369 = ~G2363;
  assign G1127 = ~G2363 | ~G2370;
  assign G2377 = ~G2371;
  assign G1135 = ~G2371 | ~G2378;
  assign G2385 = ~G2379;
  assign G1144 = ~G2379 | ~G2386;
  assign G2393 = ~G2387;
  assign G1147 = ~G2387 | ~G2394;
  assign G2401 = ~G2395;
  assign G1157 = ~G2395 | ~G2402;
  assign G2410 = ~G2406;
  assign G2418 = ~G2414;
  assign G1184 = G1628 & G1051;
  assign G2227 = ~G634 | ~G631;
  assign G2243 = ~G640 | ~G637;
  assign G2251 = G1380;
  assign G2259 = G1378;
  assign G2331 = G1382;
  assign G2339 = G1626;
  assign G2347 = G1624;
  assign G2419 = G1628;
  assign G145 = G143 | G144;
  assign G687 = ~G686;
  assign G899 = ~G2270 | ~G2273;
  assign G908 = ~G2278 | ~G2281;
  assign G916 = ~G2286 | ~G2289;
  assign G925 = ~G2294 | ~G2297;
  assign G928 = ~G2302 | ~G2305;
  assign G938 = ~G2310 | ~G2313;
  assign G954 = G1879 & G528;
  assign G961 = G1877 & G522;
  assign G1117 = ~G2358 | ~G2361;
  assign G1126 = ~G2366 | ~G2369;
  assign G1134 = ~G2374 | ~G2377;
  assign G1143 = ~G2382 | ~G2385;
  assign G1146 = ~G2390 | ~G2393;
  assign G1156 = ~G2398 | ~G2401;
  assign G1172 = G1941 & G702;
  assign G1179 = G1939 & G696;
  assign G2315 = G1879;
  assign G2323 = G1877;
  assign G2403 = G1941;
  assign G2411 = G1939;
  assign G2233 = ~G2227;
  assign G642 = ~G2227 | ~G2234;
  assign G2249 = ~G2243;
  assign G649 = ~G2243 | ~G2250;
  assign G2257 = ~G2251;
  assign G665 = ~G2251 | ~G2258;
  assign G684 = ~G2259 | ~G2266;
  assign G2265 = ~G2259;
  assign G688 = G687 & G487;
  assign G901 = ~G899 | ~G900;
  assign G910 = ~G908 | ~G909;
  assign G918 = ~G916 | ~G917;
  assign G927 = ~G925 | ~G926;
  assign G930 = ~G928 | ~G929;
  assign G940 = ~G938 | ~G939;
  assign G2337 = ~G2331;
  assign G963 = ~G2331 | ~G2338;
  assign G2345 = ~G2339;
  assign G1099 = ~G2339 | ~G2346;
  assign G1115 = ~G2347 | ~G2354;
  assign G2353 = ~G2347;
  assign G1119 = ~G1117 | ~G1118;
  assign G1128 = ~G1126 | ~G1127;
  assign G1136 = ~G1134 | ~G1135;
  assign G1145 = ~G1143 | ~G1144;
  assign G1148 = ~G1146 | ~G1147;
  assign G1158 = ~G1156 | ~G1157;
  assign G2425 = ~G2419;
  assign G1181 = ~G2419 | ~G2426;
  assign G641 = ~G2230 | ~G2233;
  assign G648 = ~G2246 | ~G2249;
  assign G664 = ~G2254 | ~G2257;
  assign G683 = ~G2262 | ~G2265;
  assign G395 = G688;
  assign G2321 = ~G2315;
  assign G948 = ~G2315 | ~G2322;
  assign G2329 = ~G2323;
  assign G956 = ~G2323 | ~G2330;
  assign G962 = ~G2334 | ~G2337;
  assign G1098 = ~G2342 | ~G2345;
  assign G1114 = ~G2350 | ~G2353;
  assign G2409 = ~G2403;
  assign G1166 = ~G2403 | ~G2410;
  assign G2417 = ~G2411;
  assign G1174 = ~G2411 | ~G2418;
  assign G1180 = ~G2422 | ~G2425;
  assign G643 = ~G641 | ~G642;
  assign G650 = ~G648 | ~G649;
  assign G666 = ~G664 | ~G665;
  assign G681 = ~G683 | ~G684;
  assign G690 = ~G688;
  assign G947 = ~G2318 | ~G2321;
  assign G955 = ~G2326 | ~G2329;
  assign G964 = ~G962 | ~G963;
  assign G968 = G901 & G918 & G910 & G927;
  assign G970 = G901 & G915;
  assign G971 = G922 & G910 & G901;
  assign G972 = G910 & G924 & G918 & G901;
  assign G978 = G930 & G946;
  assign G979 = G954 & G940 & G930;
  assign G1100 = ~G1098 | ~G1099;
  assign G1112 = ~G1114 | ~G1115;
  assign G1165 = ~G2406 | ~G2409;
  assign G1173 = ~G2414 | ~G2417;
  assign G1182 = ~G1180 | ~G1181;
  assign G1185 = G1119 & G1136 & G1128 & G1145;
  assign G1187 = G1119 & G1133;
  assign G1188 = G1140 & G1128 & G1119;
  assign G1189 = G1128 & G1142 & G1136 & G1119;
  assign G1195 = G1148 & G1164;
  assign G1196 = G1172 & G1158 & G1148;
  assign G644 = ~G643;
  assign G884 = G650 & G868;
  assign G949 = ~G947 | ~G948;
  assign G957 = ~G955 | ~G956;
  assign G969 = ~G968;
  assign G973 = G972 | G971 | G907 | G970;
  assign G1167 = ~G1165 | ~G1166;
  assign G1175 = ~G1173 | ~G1174;
  assign G1186 = ~G1185;
  assign G1190 = G1189 | G1188 | G1125 | G1187;
  assign G680 = G666 & G674;
  assign G682 = G679 & G681 & G666;
  assign G895 = G883 | G884;
  assign G1025 = G644 & G487;
  assign G1111 = G1100 & G1106;
  assign G1113 = G1110 & G1112 & G1100;
  assign G685 = G682 | G671 | G680;
  assign G295 = G895;
  assign G331 = G895;
  assign G976 = ~G973;
  assign G977 = G957 & G930 & G949 & G940 & G964;
  assign G980 = G940 & G961 & G949 & G930;
  assign G981 = G940 & G967 & G930 & G957 & G949;
  assign G397 = G1025;
  assign G1116 = G1113 | G1104 | G1111;
  assign G1193 = ~G1190;
  assign G1194 = G1175 & G1148 & G1167 & G1158 & G1182;
  assign G1197 = G1158 & G1179 & G1167 & G1148;
  assign G1198 = G1158 & G1184 & G1148 & G1175 & G1167;
  assign G982 = G981 | G980 | G979 | G937 | G978;
  assign G983 = G977 & G685;
  assign G988 = ~G976 | ~G969;
  assign G1027 = ~G1025;
  assign G1199 = G1198 | G1197 | G1196 | G1155 | G1195;
  assign G1200 = G1194 & G1116;
  assign G1205 = ~G1193 | ~G1186;
  assign G984 = G982 | G983;
  assign G1085 = G1830 & G690 & G1027;
  assign G1201 = G1199 | G1200;
  assign G987 = ~G984;
  assign G990 = G988 & G984;
  assign G1204 = ~G1201;
  assign G1207 = G1205 & G1201;
  assign G989 = G973 & G987;
  assign G1206 = G1190 & G1204;
  assign G991 = G989 | G990;
  assign G1208 = G1206 | G1207;
  assign G329 = G1208;
  assign G1221 = ~G1208 | ~G991;
  assign G1238 = G1208 & G1221;
  assign G1239 = G1221 & G991;
  assign G1240 = G1238 | G1239;
  assign G1247 = ~G1240;
  assign G471 = G1240 & G1247;
  assign G473 = G471 | G1247;
  assign G231 = ~G473;
  assign G1088 = G473 & G1553 & G1087;
  assign G1089 = G554 & G1085 & G1088;
  assign G308 = G1089;
  assign G225 = ~G1089;
endmodule


