// Benchmark "c7552_lock" written by ABC on Thu May 13 23:36:26 2021

module c7552_lock ( 
    keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
    keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
    keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
    keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
    keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
    keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
    keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
    keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
    keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
    keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
    keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
    keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
    keyinput_61, keyinput_62, keyinput_63, G9, G12, G18, G23, G26, G29,
    G32, G35, G41, G44, G47, G50, G53, G54, G55, G56, G58, G59, G60, G61,
    G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79,
    G80, G81, G82, G83, G84, G85, G86, G87, G88, G94, G97, G100, G103,
    G106, G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127,
    G130, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155,
    G156, G157, G158, G159, G160, G161, G162, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    G339, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204,
    G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256,
    G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749,
    G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437,
    G418  );
  input  keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4,
    keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9,
    keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14,
    keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19,
    keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24,
    keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29,
    keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34,
    keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39,
    keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44,
    keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49,
    keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54,
    keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59,
    keyinput_60, keyinput_61, keyinput_62, keyinput_63, G9, G12, G18, G23,
    G26, G29, G32, G35, G41, G44, G47, G50, G53, G54, G55, G56, G58, G59,
    G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77,
    G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G94, G97, G100,
    G103, G106, G109, G110, G111, G112, G113, G114, G115, G118, G121, G124,
    G127, G130, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G164, G165, G166, G167,
    G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179,
    G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191,
    G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203,
    G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215,
    G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227,
    G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239,
    G240, G339, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496,
    G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253,
    G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743,
    G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432,
    G4437;
  output G418;
  wire n1960, n2028, n1111, n1110, G406, n1113, n1112, G404, n1115, n1114,
    G408, n1117, n1116, G410, n2067, n1203, n1207, n1120, n2034, n1121,
    n1214, n2032, n1122, n1209, n2033, n1210, n1123, n1220, n1181, n1185,
    n1134, n2044, n1135, n2062, n1186, n2027, n1136, n1190, n2043, n1196,
    n1200, n1137, n2029, n1165, n1164, n1934, n1166, n1415, n2092, n1430,
    n1167, n2095, n1449, n1169, n1168, n1931, n1171, n1170, n1935, n1438,
    n1172, n2091, n1174, n1173, n1922, n1440, n1175, n2088, n1177, n1176,
    n1924, n1442, n1178, n2085, n1183, n1182, n1941, n1184, n2077, n1187,
    n2082, n1189, n1188, n1954, n1191, n2069, n1193, n1192, n1940, n1198,
    n1197, n1943, n1199, n2078, n1205, n1204, n1956, n1206, n2084, n1208,
    n2071, n1212, n1211, n1947, n1213, n2073, n1216, n1215, n1942, n1222,
    n1221, n1946, n1436, n1263, n2090, n1265, n1264, n1923, n1277, n1428,
    n1276, n1925, n1419, n1278, n2086, n1282, n1281, n1930, n1283, n1421,
    n2097, n1903, n1305, n1520, n1304, n1913, n2051, n1999, n1306, n2110,
    n1308, n1307, n1911, n1309, n2112, n1313, n1312, n1912, n1314, n2114,
    n1317, n2109, n1321, n1320, n1910, n1506, n2131, n1324, n1464, n1323,
    n1963, n1325, n2128, n1327, n1470, n1326, n1966, n1328, n2123, n1332,
    n1462, n1331, n1974, n1333, n2127, n1339, n2126, n1341, n1472, n1340,
    n1970, n1475, n1342, n2118, n1344, n1343, n1967, n1345, n1477, n2119,
    n1347, n1346, n1969, n1460, n1351, n1350, n1965, n1458, n1352, n2120,
    n1473, n1361, n2117, n1363, n1362, n1968, n1384, n1383, n1388, n1975,
    n1904, n1416, n2018, n1420, n2010, n1422, n2017, n1429, n2021, n1435,
    n2012, n1437, n2011, n1439, n2022, n1441, n2009, n1457, n1985, n2001,
    n1461, n1995, n1463, n1992, n1465, n1512, n1987, n1471, n1998, n1474,
    n1989, n1476, n1991, n1478, n1986, n1505, n2055, n1507, n2049, n1513,
    n2048, n1515, n2047, n1898, n1901, n1899, n1900, n1909, n1902, n1907,
    n1905, n1906, n1908, n1917, n1915, n1914, n1916, n1939, n1918, n1921,
    n1919, n1920, n1929, n1927, n1926, n1928, n1933, n1932, n1937, n1936,
    n1938, n1984, n1945, n1944, n1959, n1953, n1948, n1951, n1949, n1950,
    n1952, n1955, n1957, n1958, n1982, n1962, n1961, n1964, n1980, n1978,
    n1972, n1971, n1973, n1976, n1977, n1979, n1981, n1983, G414, n1988,
    n1990, n1994, n1993, n1996, n1997, n2005, n2000, n2134, n2002, n2003,
    n2004, n2026, n2006, n2101, n2007, n2008, n2016, n2014, n2013, n2015,
    n2020, n2019, n2024, n2023, n2025, n2061, n2030, n2031, n2036, n2035,
    n2042, n2037, n2040, n2038, n2039, n2041, n2046, n2045, n2059, n2050,
    n2057, n2108, n2052, n2053, n2054, n2056, n2058, n2060, G412, n2063,
    n2066, n2064, n2065, n2076, n2068, n2070, n2072, n2074, n2075, n2080,
    n2079, n2081, n2083, n2105, n2087, n2089, n2094, n2093, n2096, n2098,
    n2103, n2099, n2100, n2102, n2104, n2140, n2106, n2107, n2116, n2111,
    n2113, n2115, n2138, n2122, n2121, n2124, n2125, n2130, n2129, n2136,
    n2132, n2133, n2135, n2137, n2139, G416, n2142, n2141, n2143, n2145,
    n2144, G418_Lock, input_0, input_1, AND_1, input_2, OR_2, input_3,
    AND_3, input_4, OR_4, input_5, AND_5, input_6, AND_6, input_7, AND_7,
    input_8, OR_8, input_9, AND_9, input_10, AND_10, input_11, OR_11,
    input_12, AND_12, input_13, AND_13, input_14, AND_14, input_15, OR_15,
    input_16, AND_16, input_17, AND_17, input_18, OR_18, input_19, AND_19,
    input_20, AND_20, input_21, OR_21, input_22, AND_22, input_23, OR_23,
    input_24, OR_24, input_25, OR_25, input_26, AND_26, input_27, AND_27,
    input_28, OR_28, input_29, OR_29, input_30, OR_30, input_31, OR_31,
    input_32, input_33, AND_33, input_34, OR_34, input_35, AND_35,
    input_36, OR_36, input_37, AND_37, input_38, AND_38, input_39, AND_39,
    input_40, OR_40, input_41, AND_41, input_42, AND_42, input_43, OR_43,
    input_44, AND_44, input_45, AND_45, input_46, AND_46, input_47, OR_47,
    input_48, AND_48, input_49, AND_49, input_50, OR_50, input_51, AND_51,
    input_52, AND_52, input_53, OR_53, input_54, AND_54, input_55, OR_55,
    input_56, OR_56, input_57, OR_57, input_58, AND_58, input_59, AND_59,
    input_60, OR_60, input_61, OR_61, input_62, OR_62, input_63, OR_63,
    OR_63_INV, CASOP;
  assign n1960 = ~G18;
  assign n2028 = n1123 & n1220;
  assign n1111 = ~G152 | ~G210;
  assign n1110 = ~G218 | ~G230;
  assign G406 = n1111 | n1110;
  assign n1113 = ~G184 | ~G150;
  assign n1112 = ~G228 | ~G240;
  assign G404 = n1113 | n1112;
  assign n1115 = ~G182 | ~G183;
  assign n1114 = ~G185 | ~G186;
  assign G408 = n1115 | n1114;
  assign n1117 = ~G172 | ~G162;
  assign n1116 = ~G188 | ~G199;
  assign G410 = n1117 | n1116;
  assign n2067 = ~n2062 | ~G41;
  assign n1203 = ~G3723;
  assign n1207 = ~G103 | ~n2062;
  assign n1120 = ~G18 | ~G235;
  assign n2034 = ~n1207 | ~n1120;
  assign n1121 = ~G236 | ~G18;
  assign n1214 = ~G23 | ~n2062;
  assign n2032 = n1121 & n1214;
  assign n1122 = ~G237 | ~G18;
  assign n1209 = ~G26 | ~n2062;
  assign n2033 = ~n1122 | ~n1209;
  assign n1210 = ~G3711;
  assign n1123 = ~G238 | ~G18;
  assign n1220 = ~G29 | ~n1960;
  assign n1181 = ~G3749;
  assign n1185 = ~G100 | ~n1960;
  assign n1134 = ~G18 | ~G231;
  assign n2044 = ~n1185 | ~n1134;
  assign n1135 = ~G232 | ~G18;
  assign n2062 = ~G18;
  assign n1186 = ~G124 | ~n2062;
  assign n2027 = n1135 & n1186;
  assign n1136 = ~G233 | ~G18;
  assign n1190 = ~G127 | ~n1960;
  assign n2043 = n1136 & n1190;
  assign n1196 = ~G3729;
  assign n1200 = ~G130 | ~n1960;
  assign n1137 = ~G18 | ~G234;
  assign n2029 = ~n1200 | ~n1137;
  assign n1165 = ~G18 | ~G4437;
  assign n1164 = G18 | G62;
  assign n1934 = n1165 & n1164;
  assign n1166 = ~G189 | ~G18;
  assign n1415 = ~G66 | ~n1960;
  assign n2092 = ~n1166 | ~n1415;
  assign n1430 = ~G47 | ~n1960;
  assign n1167 = ~G18 | ~G193;
  assign n2095 = ~n1430 | ~n1167;
  assign n1449 = ~G4415;
  assign n1169 = ~G18 | ~n1449;
  assign n1168 = ~G80 | ~n1960;
  assign n1931 = ~n1169 | ~n1168;
  assign n1171 = ~G18 & ~G59;
  assign n1170 = G4405 & G18;
  assign n1935 = ~n1171 & ~n1170;
  assign n1438 = ~G94 | ~n1960;
  assign n1172 = ~G18 | ~G195;
  assign n2091 = ~n1438 | ~n1172;
  assign n1174 = ~G18 & ~G78;
  assign n1173 = G4400 & G18;
  assign n1922 = ~n1174 & ~n1173;
  assign n1440 = ~G97 | ~n2062;
  assign n1175 = ~G18 | ~G196;
  assign n2088 = ~n1440 | ~n1175;
  assign n1177 = ~G18 & ~G77;
  assign n1176 = G4394 & G18;
  assign n1924 = ~n1177 & ~n1176;
  assign n1442 = ~G118 | ~n2062;
  assign n1178 = ~G18 | ~G187;
  assign n2085 = ~n1442 | ~n1178;
  assign n1183 = ~G18 & ~G56;
  assign n1182 = ~n1181 & ~n2062;
  assign n1941 = ~n1183 & ~n1182;
  assign n1184 = ~G18 | ~G200;
  assign n2077 = ~n1185 | ~n1184;
  assign n1187 = ~G201 | ~G18;
  assign n2082 = n1187 & n1186;
  assign n1189 = ~G18 | ~G3743;
  assign n1188 = G18 | G55;
  assign n1954 = ~n1189 | ~n1188;
  assign n1191 = ~G202 | ~G18;
  assign n2069 = ~n1191 | ~n1190;
  assign n1193 = ~G18 | ~G3737;
  assign n1192 = G18 | G54;
  assign n1940 = n1193 & n1192;
  assign n1198 = ~G18 & ~G53;
  assign n1197 = ~n1196 & ~n2062;
  assign n1943 = ~n1198 & ~n1197;
  assign n1199 = ~G18 | ~G203;
  assign n2078 = ~n1200 | ~n1199;
  assign n1205 = ~G18 | ~n1203;
  assign n1204 = ~G73 | ~n2062;
  assign n1956 = ~n1205 | ~n1204;
  assign n1206 = ~G18 | ~G204;
  assign n2084 = ~n1207 | ~n1206;
  assign n1208 = ~G18 | ~G206;
  assign n2071 = ~n1209 | ~n1208;
  assign n1212 = ~G18 & ~G76;
  assign n1211 = ~n1210 & ~n2062;
  assign n1947 = ~n1212 & ~n1211;
  assign n1213 = ~G18 | ~G205;
  assign n2073 = ~n1214 | ~n1213;
  assign n1216 = ~G18 & ~G75;
  assign n1215 = G3717 & G18;
  assign n1942 = ~n1216 & ~n1215;
  assign n1222 = n1960 | G3705;
  assign n1221 = ~G74 | ~n2062;
  assign n1946 = ~n1222 | ~n1221;
  assign n1436 = ~G121 | ~n2062;
  assign n1263 = ~G18 | ~G194;
  assign n2090 = ~n1436 | ~n1263;
  assign n1265 = ~G18 & ~G81;
  assign n1264 = G4410 & G18;
  assign n1923 = ~n1265 & ~n1264;
  assign n1277 = ~G18 & ~G79;
  assign n1428 = ~G4420;
  assign n1276 = ~n1428 & ~n2062;
  assign n1925 = ~n1277 & ~n1276;
  assign n1419 = ~G35 | ~n2062;
  assign n1278 = ~G18 | ~G192;
  assign n2086 = ~n1419 | ~n1278;
  assign n1282 = ~G18 | ~G4427;
  assign n1281 = G18 | G60;
  assign n1930 = ~n1282 | ~n1281;
  assign n1283 = ~G191 | ~G18;
  assign n1421 = ~G32 | ~n2062;
  assign n2097 = n1283 & n1421;
  assign n1903 = ~G2204 & ~G1455;
  assign n1305 = ~G18 & ~G88;
  assign n1520 = ~G1486;
  assign n1304 = ~n1520 & ~n2062;
  assign n1913 = ~n1305 & ~n1304;
  assign n2051 = ~G12 | ~G9;
  assign n1999 = ~n2051;
  assign n1306 = ~G166 & ~n2062;
  assign n2110 = ~n1999 & ~n1306;
  assign n1308 = ~G18 & ~G112;
  assign n1307 = G1480 & G18;
  assign n1911 = ~n1308 & ~n1307;
  assign n1309 = ~G167 & ~n2062;
  assign n2112 = ~n1999 & ~n1309;
  assign n1313 = ~G18 & ~G111;
  assign n1312 = G1469 & G18;
  assign n1912 = ~n1313 & ~n1312;
  assign n1314 = ~G169 & ~n2062;
  assign n2114 = ~n1999 & ~n1314;
  assign n1317 = ~G168 & ~n2062;
  assign n2109 = ~n1999 & ~n1317;
  assign n1321 = ~G18 | ~G1462;
  assign n1320 = G18 | G113;
  assign n1910 = ~n1321 | ~n1320;
  assign n1506 = ~G18 & ~n1999;
  assign n2131 = G173 & n2051;
  assign n1324 = ~G18 & ~G86;
  assign n1464 = ~G2247;
  assign n1323 = ~n1464 & ~n2062;
  assign n1963 = ~n1324 & ~n1323;
  assign n1325 = ~G175 & ~n2062;
  assign n2128 = ~n1999 & ~n1325;
  assign n1327 = ~G18 & ~G63;
  assign n1470 = ~G2239;
  assign n1326 = ~n1470 & ~n2062;
  assign n1966 = ~n1327 & ~n1326;
  assign n1328 = ~G176 & ~n2062;
  assign n2123 = ~n1999 & ~n1328;
  assign n1332 = ~G18 & ~G109;
  assign n1462 = ~G2253;
  assign n1331 = ~n1462 & ~n2062;
  assign n1974 = ~n1332 & ~n1331;
  assign n1333 = ~G174 & ~n2062;
  assign n2127 = ~n1999 & ~n1333;
  assign n1339 = ~G177 & ~n2062;
  assign n2126 = ~n1999 & ~n1339;
  assign n1341 = ~G18 & ~G64;
  assign n1472 = ~G2236;
  assign n1340 = ~n1472 & ~n2062;
  assign n1970 = ~n1341 & ~n1340;
  assign n1475 = ~G144 | ~n1960;
  assign n1342 = ~G18 | ~G179;
  assign n2118 = ~n1475 | ~n1342;
  assign n1344 = ~G18 & ~G84;
  assign n1343 = G2224 & G18;
  assign n1967 = ~n1344 & ~n1343;
  assign n1345 = ~G180 | ~G18;
  assign n1477 = ~G138 | ~n1960;
  assign n2119 = ~n1345 | ~n1477;
  assign n1347 = ~G18 | ~G2218;
  assign n1346 = G18 | G83;
  assign n1969 = n1347 & n1346;
  assign n1460 = ~G2211;
  assign n1351 = ~G18 | ~n1460;
  assign n1350 = ~G65 | ~n1960;
  assign n1965 = ~n1351 | ~n1350;
  assign n1458 = ~G147 | ~n1960;
  assign n1352 = ~G18 | ~G171;
  assign n2120 = ~n1458 | ~n1352;
  assign n1473 = ~G135 | ~n2062;
  assign n1361 = ~G18 | ~G178;
  assign n2117 = ~n1473 | ~n1361;
  assign n1363 = ~G18 & ~G85;
  assign n1362 = G2230 & G18;
  assign n1968 = ~n1363 & ~n1362;
  assign n1384 = ~G18 | ~G2256;
  assign n1383 = G18 | G110;
  assign n1388 = ~n1384 | ~n1383;
  assign n1975 = ~n1388;
  assign n1904 = G2204 & G1455;
  assign n1416 = ~G219 | ~G18;
  assign n2018 = ~n1416 | ~n1415;
  assign n1420 = ~G222 | ~G18;
  assign n2010 = ~n1420 | ~n1419;
  assign n1422 = ~G221 | ~G18;
  assign n2017 = n1422 & n1421;
  assign n1429 = ~G18 | ~G223;
  assign n2021 = ~n1430 | ~n1429;
  assign n1435 = ~G18 | ~G224;
  assign n2012 = n1436 & n1435;
  assign n1437 = ~G18 | ~G225;
  assign n2011 = n1438 & n1437;
  assign n1439 = ~G18 | ~G226;
  assign n2022 = n1440 & n1439;
  assign n1441 = ~G18 | ~G217;
  assign n2009 = n1442 & n1441;
  assign n1457 = ~G18 | ~G151;
  assign n1985 = ~n1458 | ~n1457;
  assign n2001 = G153 & n2051;
  assign n1461 = ~G154 & ~n2062;
  assign n1995 = ~n1999 & ~n1461;
  assign n1463 = ~G155 & ~n2062;
  assign n1992 = ~n1999 & ~n1463;
  assign n1465 = ~n2051 | ~G156;
  assign n1512 = ~n1506;
  assign n1987 = ~n1465 | ~n1512;
  assign n1471 = ~G157 & ~n2062;
  assign n1998 = ~n1999 & ~n1471;
  assign n1474 = ~G158 | ~G18;
  assign n1989 = ~n1474 | ~n1473;
  assign n1476 = ~G159 | ~G18;
  assign n1991 = ~n1476 | ~n1475;
  assign n1478 = ~G160 | ~G18;
  assign n1986 = n1478 & n1477;
  assign n1505 = n1506 | G215;
  assign n2055 = ~n2051 | ~n1505;
  assign n1507 = n1506 | G216;
  assign n2049 = ~n2051 | ~n1507;
  assign n1513 = ~n2051 | ~G214;
  assign n2048 = n1513 & n1512;
  assign n1515 = ~G213 & ~n2062;
  assign n2047 = ~n1999 & ~n1515;
  assign n1898 = ~G1459 ^ G106;
  assign n1901 = ~n1898 | ~G18;
  assign n1899 = ~G87 ^ G114;
  assign n1900 = ~n1960 | ~n1899;
  assign n1909 = ~n1901 | ~n1900;
  assign n1902 = G1492 ^ G1496;
  assign n1907 = ~n2062 & ~n1902;
  assign n1905 = ~n1904 & ~n1903;
  assign n1906 = ~G18 & ~n1905;
  assign n1908 = ~n1907 & ~n1906;
  assign n1917 = ~n1909 ^ n1908;
  assign n1915 = ~n1911 ^ n1910;
  assign n1914 = ~n1913 ^ n1912;
  assign n1916 = ~n1915 ^ n1914;
  assign n1939 = ~n1917 ^ n1916;
  assign n1918 = G4432 ^ G4393;
  assign n1921 = ~n1918 | ~G18;
  assign n1919 = G61 ^ G58;
  assign n1920 = ~n2062 | ~n1919;
  assign n1929 = ~n1921 | ~n1920;
  assign n1927 = n1923 ^ n1922;
  assign n1926 = ~n1925 ^ n1924;
  assign n1928 = ~n1927 ^ n1926;
  assign n1933 = ~n1929 ^ n1928;
  assign n1932 = n1931 ^ n1930;
  assign n1937 = ~n1933 ^ n1932;
  assign n1936 = ~n1935 ^ n1934;
  assign n1938 = ~n1937 ^ n1936;
  assign n1984 = ~n1939 & ~n1938;
  assign n1945 = n1941 ^ n1940;
  assign n1944 = ~n1943 ^ n1942;
  assign n1959 = ~n1945 ^ n1944;
  assign n1953 = ~n1947 ^ n1946;
  assign n1948 = ~G3698 ^ G3701;
  assign n1951 = ~n1948 | ~G18;
  assign n1949 = ~G70 ^ G69;
  assign n1950 = ~n2062 | ~n1949;
  assign n1952 = ~n1951 | ~n1950;
  assign n1955 = ~n1953 ^ n1952;
  assign n1957 = ~n1955 ^ n1954;
  assign n1958 = ~n1957 ^ n1956;
  assign n1982 = ~n1959 ^ n1958;
  assign n1962 = G2208 | n1960;
  assign n1961 = ~G82 | ~n2062;
  assign n1964 = ~n1962 | ~n1961;
  assign n1980 = ~n1964 ^ n1963;
  assign n1978 = ~n1966 ^ n1965;
  assign n1972 = n1968 ^ n1967;
  assign n1971 = ~n1970 ^ n1969;
  assign n1973 = ~n1972 ^ n1971;
  assign n1976 = ~n1974 ^ n1973;
  assign n1977 = n1976 ^ n1975;
  assign n1979 = ~n1978 ^ n1977;
  assign n1981 = ~n1980 ^ n1979;
  assign n1983 = ~n1982 & ~n1981;
  assign G414 = ~n1984 | ~n1983;
  assign n1988 = n1986 ^ n1985;
  assign n1990 = n1988 ^ n1987;
  assign n1994 = ~n1990 ^ n1989;
  assign n1993 = n1992 ^ n1991;
  assign n1996 = ~n1994 ^ n1993;
  assign n1997 = n1996 ^ n1995;
  assign n2005 = ~n1998 ^ n1997;
  assign n2000 = G141 ^ n1999;
  assign n2134 = ~G18 & ~n2000;
  assign n2002 = ~G161 ^ n2001;
  assign n2003 = ~n1960 & ~n2002;
  assign n2004 = ~n2134 & ~n2003;
  assign n2026 = n2005 ^ n2004;
  assign n2006 = ~G50 ^ G115;
  assign n2101 = ~n2006 | ~n2062;
  assign n2007 = ~G220 ^ G227;
  assign n2008 = ~G18 | ~n2007;
  assign n2016 = ~n2101 | ~n2008;
  assign n2014 = ~n2010 ^ n2009;
  assign n2013 = ~n2012 ^ n2011;
  assign n2015 = ~n2014 ^ n2013;
  assign n2020 = ~n2016 ^ n2015;
  assign n2019 = n2018 ^ n2017;
  assign n2024 = ~n2020 ^ n2019;
  assign n2023 = ~n2022 ^ n2021;
  assign n2025 = ~n2024 ^ n2023;
  assign n2061 = ~n2026 & ~n2025;
  assign n2030 = n2028 ^ n2027;
  assign n2031 = ~n2030 ^ n2029;
  assign n2036 = ~n2032 ^ n2031;
  assign n2035 = n2034 ^ n2033;
  assign n2042 = ~n2036 ^ n2035;
  assign n2037 = ~G41 ^ G44;
  assign n2040 = ~n2037 | ~n2062;
  assign n2038 = ~G229 ^ G239;
  assign n2039 = ~G18 | ~n2038;
  assign n2041 = ~n2040 | ~n2039;
  assign n2046 = n2042 ^ n2041;
  assign n2045 = n2044 ^ n2043;
  assign n2059 = ~n2046 ^ n2045;
  assign n2050 = ~n2048 ^ n2047;
  assign n2057 = ~n2050 ^ n2049;
  assign n2108 = ~G18 | ~n2051;
  assign n2052 = ~G212 ^ G209;
  assign n2053 = ~G211 ^ n2052;
  assign n2054 = ~n2108 & ~n2053;
  assign n2056 = n2055 ^ n2054;
  assign n2058 = ~n2057 ^ n2056;
  assign n2060 = ~n2059 & ~n2058;
  assign G412 = ~n2061 | ~n2060;
  assign n2063 = ~G29 ^ G44;
  assign n2066 = ~n2063 | ~n2062;
  assign n2064 = ~G207 ^ G208;
  assign n2065 = ~G18 | ~n2064;
  assign n2076 = ~n2066 | ~n2065;
  assign n2068 = ~G198 | ~G18;
  assign n2070 = ~n2068 | ~n2067;
  assign n2072 = n2070 ^ n2069;
  assign n2074 = ~n2072 ^ n2071;
  assign n2075 = ~n2074 ^ n2073;
  assign n2080 = ~n2076 ^ n2075;
  assign n2079 = n2078 ^ n2077;
  assign n2081 = ~n2080 ^ n2079;
  assign n2083 = n2082 ^ n2081;
  assign n2105 = ~n2084 ^ n2083;
  assign n2087 = n2086 ^ n2085;
  assign n2089 = ~n2088 ^ n2087;
  assign n2094 = ~n2090 ^ n2089;
  assign n2093 = ~n2092 ^ n2091;
  assign n2096 = ~n2094 ^ n2093;
  assign n2098 = ~n2096 ^ n2095;
  assign n2103 = n2098 ^ n2097;
  assign n2099 = ~G190 ^ G197;
  assign n2100 = ~G18 | ~n2099;
  assign n2102 = ~n2101 | ~n2100;
  assign n2104 = n2103 ^ n2102;
  assign n2140 = ~n2105 & ~n2104;
  assign n2106 = ~G170 ^ G164;
  assign n2107 = ~n2106 ^ G165;
  assign n2116 = ~n2108 & ~n2107;
  assign n2111 = n2110 ^ n2109;
  assign n2113 = ~n2112 ^ n2111;
  assign n2115 = n2114 ^ n2113;
  assign n2138 = ~n2116 ^ n2115;
  assign n2122 = ~n2118 ^ n2117;
  assign n2121 = n2120 ^ n2119;
  assign n2124 = ~n2122 ^ n2121;
  assign n2125 = n2124 ^ n2123;
  assign n2130 = ~n2126 ^ n2125;
  assign n2129 = n2128 ^ n2127;
  assign n2136 = ~n2130 ^ n2129;
  assign n2132 = ~G181 ^ n2131;
  assign n2133 = ~n2062 & ~n2132;
  assign n2135 = ~n2134 & ~n2133;
  assign n2137 = n2136 ^ n2135;
  assign n2139 = ~n2138 & ~n2137;
  assign G416 = ~n2140 | ~n2139;
  assign n2142 = ~G410 & ~G408;
  assign n2141 = ~G404 & ~G406;
  assign n2143 = ~n2142 | ~n2141;
  assign n2145 = ~G414 & ~n2143;
  assign n2144 = ~G412 & ~G416;
  assign G418_Lock = ~n2145 | ~n2144;
  assign input_0 = keyinput_0 ^ G9;
  assign input_1 = keyinput_1 ^ G12;
  assign AND_1 = input_0 & input_1;
  assign input_2 = ~keyinput_2 ^ G18;
  assign OR_2 = input_2 | AND_1;
  assign input_3 = keyinput_3 ^ G23;
  assign AND_3 = input_3 & OR_2;
  assign input_4 = keyinput_4 ^ G26;
  assign OR_4 = input_4 | AND_3;
  assign input_5 = keyinput_5 ^ G29;
  assign AND_5 = input_5 & OR_4;
  assign input_6 = ~keyinput_6 ^ G32;
  assign AND_6 = input_6 & AND_5;
  assign input_7 = ~keyinput_7 ^ G35;
  assign AND_7 = input_7 & AND_6;
  assign input_8 = keyinput_8 ^ G41;
  assign OR_8 = input_8 | AND_7;
  assign input_9 = keyinput_9 ^ G44;
  assign AND_9 = input_9 & OR_8;
  assign input_10 = keyinput_10 ^ G47;
  assign AND_10 = input_10 & AND_9;
  assign input_11 = ~keyinput_11 ^ G50;
  assign OR_11 = input_11 | AND_10;
  assign input_12 = ~keyinput_12 ^ G53;
  assign AND_12 = input_12 & OR_11;
  assign input_13 = ~keyinput_13 ^ G54;
  assign AND_13 = input_13 & AND_12;
  assign input_14 = ~keyinput_14 ^ G55;
  assign AND_14 = input_14 & AND_13;
  assign input_15 = ~keyinput_15 ^ G56;
  assign OR_15 = input_15 | AND_14;
  assign input_16 = ~keyinput_16 ^ G58;
  assign AND_16 = input_16 & OR_15;
  assign input_17 = ~keyinput_17 ^ G59;
  assign AND_17 = input_17 & AND_16;
  assign input_18 = keyinput_18 ^ G60;
  assign OR_18 = input_18 | AND_17;
  assign input_19 = keyinput_19 ^ G61;
  assign AND_19 = input_19 & OR_18;
  assign input_20 = ~keyinput_20 ^ G62;
  assign AND_20 = input_20 & AND_19;
  assign input_21 = ~keyinput_21 ^ G63;
  assign OR_21 = input_21 | AND_20;
  assign input_22 = keyinput_22 ^ G64;
  assign AND_22 = input_22 & OR_21;
  assign input_23 = keyinput_23 ^ G65;
  assign OR_23 = input_23 | AND_22;
  assign input_24 = ~keyinput_24 ^ G66;
  assign OR_24 = input_24 | OR_23;
  assign input_25 = ~keyinput_25 ^ G69;
  assign OR_25 = input_25 | OR_24;
  assign input_26 = keyinput_26 ^ G70;
  assign AND_26 = input_26 & OR_25;
  assign input_27 = keyinput_27 ^ G73;
  assign AND_27 = input_27 & AND_26;
  assign input_28 = keyinput_28 ^ G74;
  assign OR_28 = input_28 | AND_27;
  assign input_29 = ~keyinput_29 ^ G75;
  assign OR_29 = input_29 | OR_28;
  assign input_30 = keyinput_30 ^ G76;
  assign OR_30 = input_30 | OR_29;
  assign input_31 = ~keyinput_31 ^ G77;
  assign OR_31 = input_31 | OR_30;
  assign input_32 = keyinput_32 ^ G9;
  assign input_33 = keyinput_33 ^ G12;
  assign AND_33 = input_32 & input_33;
  assign input_34 = keyinput_34 ^ G18;
  assign OR_34 = input_34 | AND_33;
  assign input_35 = keyinput_35 ^ G23;
  assign AND_35 = input_35 & OR_34;
  assign input_36 = keyinput_36 ^ G26;
  assign OR_36 = input_36 | AND_35;
  assign input_37 = ~keyinput_37 ^ G29;
  assign AND_37 = input_37 & OR_36;
  assign input_38 = ~keyinput_38 ^ G32;
  assign AND_38 = input_38 & AND_37;
  assign input_39 = ~keyinput_39 ^ G35;
  assign AND_39 = input_39 & AND_38;
  assign input_40 = ~keyinput_40 ^ G41;
  assign OR_40 = input_40 | AND_39;
  assign input_41 = keyinput_41 ^ G44;
  assign AND_41 = input_41 & OR_40;
  assign input_42 = ~keyinput_42 ^ G47;
  assign AND_42 = input_42 & AND_41;
  assign input_43 = keyinput_43 ^ G50;
  assign OR_43 = input_43 | AND_42;
  assign input_44 = keyinput_44 ^ G53;
  assign AND_44 = input_44 & OR_43;
  assign input_45 = ~keyinput_45 ^ G54;
  assign AND_45 = input_45 & AND_44;
  assign input_46 = keyinput_46 ^ G55;
  assign AND_46 = input_46 & AND_45;
  assign input_47 = keyinput_47 ^ G56;
  assign OR_47 = input_47 | AND_46;
  assign input_48 = keyinput_48 ^ G58;
  assign AND_48 = input_48 & OR_47;
  assign input_49 = ~keyinput_49 ^ G59;
  assign AND_49 = input_49 & AND_48;
  assign input_50 = ~keyinput_50 ^ G60;
  assign OR_50 = input_50 | AND_49;
  assign input_51 = keyinput_51 ^ G61;
  assign AND_51 = input_51 & OR_50;
  assign input_52 = ~keyinput_52 ^ G62;
  assign AND_52 = input_52 & AND_51;
  assign input_53 = keyinput_53 ^ G63;
  assign OR_53 = input_53 | AND_52;
  assign input_54 = ~keyinput_54 ^ G64;
  assign AND_54 = input_54 & OR_53;
  assign input_55 = ~keyinput_55 ^ G65;
  assign OR_55 = input_55 | AND_54;
  assign input_56 = ~keyinput_56 ^ G66;
  assign OR_56 = input_56 | OR_55;
  assign input_57 = keyinput_57 ^ G69;
  assign OR_57 = input_57 | OR_56;
  assign input_58 = ~keyinput_58 ^ G70;
  assign AND_58 = input_58 & OR_57;
  assign input_59 = ~keyinput_59 ^ G73;
  assign AND_59 = input_59 & AND_58;
  assign input_60 = ~keyinput_60 ^ G74;
  assign OR_60 = input_60 | AND_59;
  assign input_61 = keyinput_61 ^ G75;
  assign OR_61 = input_61 | OR_60;
  assign input_62 = ~keyinput_62 ^ G76;
  assign OR_62 = input_62 | OR_61;
  assign input_63 = keyinput_63 ^ G77;
  assign OR_63 = input_63 | OR_62;
  assign OR_63_INV = ~OR_63;
  assign CASOP = OR_31 & OR_63_INV;
  assign G418 = G418_Lock ^ CASOP;
endmodule


