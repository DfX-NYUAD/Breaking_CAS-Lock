// Benchmark "b15_C_lock" written by ABC on Thu May 13 23:39:34 2021

module b15_C_lock ( 
    READY_N, STATEBS16_REG_SCAN_IN, REIP_REG_31__SCAN_IN,
    REIP_REG_30__SCAN_IN, REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN,
    REIP_REG_27__SCAN_IN, REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN,
    REIP_REG_24__SCAN_IN, REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN,
    REIP_REG_21__SCAN_IN, REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN,
    REIP_REG_18__SCAN_IN, REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN,
    STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN,
    STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN,
    STATE2_REG_0__SCAN_IN, INSTQUEUE_REG_15__7__SCAN_IN,
    INSTQUEUE_REG_15__6__SCAN_IN, INSTQUEUE_REG_15__5__SCAN_IN,
    INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUE_REG_15__3__SCAN_IN,
    INSTQUEUE_REG_15__2__SCAN_IN, INSTQUEUE_REG_15__1__SCAN_IN,
    INSTQUEUE_REG_15__0__SCAN_IN, INSTQUEUE_REG_14__7__SCAN_IN,
    INSTQUEUE_REG_14__6__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN,
    INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUE_REG_14__3__SCAN_IN,
    INSTQUEUE_REG_14__2__SCAN_IN, INSTQUEUE_REG_14__1__SCAN_IN,
    INSTQUEUE_REG_14__0__SCAN_IN, INSTQUEUE_REG_13__7__SCAN_IN,
    INSTQUEUE_REG_13__6__SCAN_IN, INSTQUEUE_REG_13__5__SCAN_IN,
    INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUE_REG_13__3__SCAN_IN,
    INSTQUEUE_REG_13__2__SCAN_IN, INSTQUEUE_REG_13__1__SCAN_IN,
    INSTQUEUE_REG_13__0__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN,
    INSTQUEUE_REG_12__6__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN,
    INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUE_REG_12__3__SCAN_IN,
    INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_12__1__SCAN_IN,
    INSTQUEUE_REG_12__0__SCAN_IN, INSTQUEUE_REG_11__7__SCAN_IN,
    INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUE_REG_11__5__SCAN_IN,
    INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN,
    INSTQUEUE_REG_11__2__SCAN_IN, INSTQUEUE_REG_11__1__SCAN_IN,
    INSTQUEUE_REG_11__0__SCAN_IN, INSTQUEUE_REG_10__7__SCAN_IN,
    INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUE_REG_10__5__SCAN_IN,
    INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUE_REG_10__3__SCAN_IN,
    INSTQUEUE_REG_10__2__SCAN_IN, INSTQUEUE_REG_10__1__SCAN_IN,
    INSTQUEUE_REG_10__0__SCAN_IN, INSTQUEUE_REG_9__7__SCAN_IN,
    INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN,
    INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN,
    INSTQUEUE_REG_9__2__SCAN_IN, INSTQUEUE_REG_9__1__SCAN_IN,
    INSTQUEUE_REG_9__0__SCAN_IN, INSTQUEUE_REG_8__7__SCAN_IN,
    INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUE_REG_8__5__SCAN_IN,
    INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUE_REG_8__3__SCAN_IN,
    INSTQUEUE_REG_8__2__SCAN_IN, INSTQUEUE_REG_8__1__SCAN_IN,
    INSTQUEUE_REG_8__0__SCAN_IN, INSTQUEUE_REG_7__7__SCAN_IN,
    INSTQUEUE_REG_7__6__SCAN_IN, INSTQUEUE_REG_7__5__SCAN_IN,
    INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUE_REG_7__3__SCAN_IN,
    INSTQUEUE_REG_7__2__SCAN_IN, INSTQUEUE_REG_7__1__SCAN_IN,
    INSTQUEUE_REG_7__0__SCAN_IN, INSTQUEUE_REG_6__7__SCAN_IN,
    INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_6__5__SCAN_IN,
    INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUE_REG_6__3__SCAN_IN,
    INSTQUEUE_REG_6__2__SCAN_IN, INSTQUEUE_REG_6__1__SCAN_IN,
    INSTQUEUE_REG_6__0__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN,
    INSTQUEUE_REG_5__6__SCAN_IN, INSTQUEUE_REG_5__5__SCAN_IN,
    INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUE_REG_5__3__SCAN_IN,
    INSTQUEUE_REG_5__2__SCAN_IN, INSTQUEUE_REG_5__1__SCAN_IN,
    INSTQUEUE_REG_5__0__SCAN_IN, INSTQUEUE_REG_4__7__SCAN_IN,
    INSTQUEUE_REG_4__6__SCAN_IN, INSTQUEUE_REG_4__5__SCAN_IN,
    INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUE_REG_4__3__SCAN_IN,
    INSTQUEUE_REG_4__2__SCAN_IN, INSTQUEUE_REG_4__1__SCAN_IN,
    INSTQUEUE_REG_4__0__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN,
    INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUE_REG_3__5__SCAN_IN,
    INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUE_REG_3__3__SCAN_IN,
    INSTQUEUE_REG_3__2__SCAN_IN, INSTQUEUE_REG_3__1__SCAN_IN,
    INSTQUEUE_REG_3__0__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN,
    INSTQUEUE_REG_2__6__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN,
    INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUE_REG_2__3__SCAN_IN,
    INSTQUEUE_REG_2__2__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN,
    INSTQUEUE_REG_2__0__SCAN_IN, INSTQUEUE_REG_1__7__SCAN_IN,
    INSTQUEUE_REG_1__6__SCAN_IN, INSTQUEUE_REG_1__5__SCAN_IN,
    INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN,
    INSTQUEUE_REG_1__2__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN,
    INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN,
    INSTQUEUE_REG_0__6__SCAN_IN, INSTQUEUE_REG_0__5__SCAN_IN,
    INSTQUEUE_REG_0__4__SCAN_IN, INSTQUEUE_REG_0__3__SCAN_IN,
    INSTQUEUE_REG_0__2__SCAN_IN, INSTQUEUE_REG_0__1__SCAN_IN,
    INSTQUEUE_REG_0__0__SCAN_IN, INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_4__SCAN_IN, INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_2__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
    INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
    INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
    INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
    INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
    INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
    INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
    INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
    INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
    INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
    INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
    INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
    INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
    INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
    INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
    INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
    PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
    PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
    PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
    PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
    PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
    PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
    PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
    PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
    PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
    PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
    PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
    PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
    PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
    PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
    PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
    PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
    EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
    EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
    EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
    EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
    EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
    EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
    EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
    EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
    EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
    EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
    EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
    EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
    EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
    EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
    EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
    EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
    EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
    EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
    EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
    EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
    EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
    EBX_REG_31__SCAN_IN, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN,
    REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, REIP_REG_5__SCAN_IN,
    REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, REIP_REG_8__SCAN_IN,
    REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, REIP_REG_11__SCAN_IN,
    REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, REIP_REG_14__SCAN_IN,
    REIP_REG_15__SCAN_IN,
    U2796  );
  input  READY_N, STATEBS16_REG_SCAN_IN, REIP_REG_31__SCAN_IN,
    REIP_REG_30__SCAN_IN, REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN,
    REIP_REG_27__SCAN_IN, REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN,
    REIP_REG_24__SCAN_IN, REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN,
    REIP_REG_21__SCAN_IN, REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN,
    REIP_REG_18__SCAN_IN, REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN,
    STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN,
    STATE2_REG_3__SCAN_IN, STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN,
    STATE2_REG_0__SCAN_IN, INSTQUEUE_REG_15__7__SCAN_IN,
    INSTQUEUE_REG_15__6__SCAN_IN, INSTQUEUE_REG_15__5__SCAN_IN,
    INSTQUEUE_REG_15__4__SCAN_IN, INSTQUEUE_REG_15__3__SCAN_IN,
    INSTQUEUE_REG_15__2__SCAN_IN, INSTQUEUE_REG_15__1__SCAN_IN,
    INSTQUEUE_REG_15__0__SCAN_IN, INSTQUEUE_REG_14__7__SCAN_IN,
    INSTQUEUE_REG_14__6__SCAN_IN, INSTQUEUE_REG_14__5__SCAN_IN,
    INSTQUEUE_REG_14__4__SCAN_IN, INSTQUEUE_REG_14__3__SCAN_IN,
    INSTQUEUE_REG_14__2__SCAN_IN, INSTQUEUE_REG_14__1__SCAN_IN,
    INSTQUEUE_REG_14__0__SCAN_IN, INSTQUEUE_REG_13__7__SCAN_IN,
    INSTQUEUE_REG_13__6__SCAN_IN, INSTQUEUE_REG_13__5__SCAN_IN,
    INSTQUEUE_REG_13__4__SCAN_IN, INSTQUEUE_REG_13__3__SCAN_IN,
    INSTQUEUE_REG_13__2__SCAN_IN, INSTQUEUE_REG_13__1__SCAN_IN,
    INSTQUEUE_REG_13__0__SCAN_IN, INSTQUEUE_REG_12__7__SCAN_IN,
    INSTQUEUE_REG_12__6__SCAN_IN, INSTQUEUE_REG_12__5__SCAN_IN,
    INSTQUEUE_REG_12__4__SCAN_IN, INSTQUEUE_REG_12__3__SCAN_IN,
    INSTQUEUE_REG_12__2__SCAN_IN, INSTQUEUE_REG_12__1__SCAN_IN,
    INSTQUEUE_REG_12__0__SCAN_IN, INSTQUEUE_REG_11__7__SCAN_IN,
    INSTQUEUE_REG_11__6__SCAN_IN, INSTQUEUE_REG_11__5__SCAN_IN,
    INSTQUEUE_REG_11__4__SCAN_IN, INSTQUEUE_REG_11__3__SCAN_IN,
    INSTQUEUE_REG_11__2__SCAN_IN, INSTQUEUE_REG_11__1__SCAN_IN,
    INSTQUEUE_REG_11__0__SCAN_IN, INSTQUEUE_REG_10__7__SCAN_IN,
    INSTQUEUE_REG_10__6__SCAN_IN, INSTQUEUE_REG_10__5__SCAN_IN,
    INSTQUEUE_REG_10__4__SCAN_IN, INSTQUEUE_REG_10__3__SCAN_IN,
    INSTQUEUE_REG_10__2__SCAN_IN, INSTQUEUE_REG_10__1__SCAN_IN,
    INSTQUEUE_REG_10__0__SCAN_IN, INSTQUEUE_REG_9__7__SCAN_IN,
    INSTQUEUE_REG_9__6__SCAN_IN, INSTQUEUE_REG_9__5__SCAN_IN,
    INSTQUEUE_REG_9__4__SCAN_IN, INSTQUEUE_REG_9__3__SCAN_IN,
    INSTQUEUE_REG_9__2__SCAN_IN, INSTQUEUE_REG_9__1__SCAN_IN,
    INSTQUEUE_REG_9__0__SCAN_IN, INSTQUEUE_REG_8__7__SCAN_IN,
    INSTQUEUE_REG_8__6__SCAN_IN, INSTQUEUE_REG_8__5__SCAN_IN,
    INSTQUEUE_REG_8__4__SCAN_IN, INSTQUEUE_REG_8__3__SCAN_IN,
    INSTQUEUE_REG_8__2__SCAN_IN, INSTQUEUE_REG_8__1__SCAN_IN,
    INSTQUEUE_REG_8__0__SCAN_IN, INSTQUEUE_REG_7__7__SCAN_IN,
    INSTQUEUE_REG_7__6__SCAN_IN, INSTQUEUE_REG_7__5__SCAN_IN,
    INSTQUEUE_REG_7__4__SCAN_IN, INSTQUEUE_REG_7__3__SCAN_IN,
    INSTQUEUE_REG_7__2__SCAN_IN, INSTQUEUE_REG_7__1__SCAN_IN,
    INSTQUEUE_REG_7__0__SCAN_IN, INSTQUEUE_REG_6__7__SCAN_IN,
    INSTQUEUE_REG_6__6__SCAN_IN, INSTQUEUE_REG_6__5__SCAN_IN,
    INSTQUEUE_REG_6__4__SCAN_IN, INSTQUEUE_REG_6__3__SCAN_IN,
    INSTQUEUE_REG_6__2__SCAN_IN, INSTQUEUE_REG_6__1__SCAN_IN,
    INSTQUEUE_REG_6__0__SCAN_IN, INSTQUEUE_REG_5__7__SCAN_IN,
    INSTQUEUE_REG_5__6__SCAN_IN, INSTQUEUE_REG_5__5__SCAN_IN,
    INSTQUEUE_REG_5__4__SCAN_IN, INSTQUEUE_REG_5__3__SCAN_IN,
    INSTQUEUE_REG_5__2__SCAN_IN, INSTQUEUE_REG_5__1__SCAN_IN,
    INSTQUEUE_REG_5__0__SCAN_IN, INSTQUEUE_REG_4__7__SCAN_IN,
    INSTQUEUE_REG_4__6__SCAN_IN, INSTQUEUE_REG_4__5__SCAN_IN,
    INSTQUEUE_REG_4__4__SCAN_IN, INSTQUEUE_REG_4__3__SCAN_IN,
    INSTQUEUE_REG_4__2__SCAN_IN, INSTQUEUE_REG_4__1__SCAN_IN,
    INSTQUEUE_REG_4__0__SCAN_IN, INSTQUEUE_REG_3__7__SCAN_IN,
    INSTQUEUE_REG_3__6__SCAN_IN, INSTQUEUE_REG_3__5__SCAN_IN,
    INSTQUEUE_REG_3__4__SCAN_IN, INSTQUEUE_REG_3__3__SCAN_IN,
    INSTQUEUE_REG_3__2__SCAN_IN, INSTQUEUE_REG_3__1__SCAN_IN,
    INSTQUEUE_REG_3__0__SCAN_IN, INSTQUEUE_REG_2__7__SCAN_IN,
    INSTQUEUE_REG_2__6__SCAN_IN, INSTQUEUE_REG_2__5__SCAN_IN,
    INSTQUEUE_REG_2__4__SCAN_IN, INSTQUEUE_REG_2__3__SCAN_IN,
    INSTQUEUE_REG_2__2__SCAN_IN, INSTQUEUE_REG_2__1__SCAN_IN,
    INSTQUEUE_REG_2__0__SCAN_IN, INSTQUEUE_REG_1__7__SCAN_IN,
    INSTQUEUE_REG_1__6__SCAN_IN, INSTQUEUE_REG_1__5__SCAN_IN,
    INSTQUEUE_REG_1__4__SCAN_IN, INSTQUEUE_REG_1__3__SCAN_IN,
    INSTQUEUE_REG_1__2__SCAN_IN, INSTQUEUE_REG_1__1__SCAN_IN,
    INSTQUEUE_REG_1__0__SCAN_IN, INSTQUEUE_REG_0__7__SCAN_IN,
    INSTQUEUE_REG_0__6__SCAN_IN, INSTQUEUE_REG_0__5__SCAN_IN,
    INSTQUEUE_REG_0__4__SCAN_IN, INSTQUEUE_REG_0__3__SCAN_IN,
    INSTQUEUE_REG_0__2__SCAN_IN, INSTQUEUE_REG_0__1__SCAN_IN,
    INSTQUEUE_REG_0__0__SCAN_IN, INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    INSTQUEUERD_ADDR_REG_3__SCAN_IN, INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    INSTQUEUERD_ADDR_REG_1__SCAN_IN, INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_4__SCAN_IN, INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_2__SCAN_IN, INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
    INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
    INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
    INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
    INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
    INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
    INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
    INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
    INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
    INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
    INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
    INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
    INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
    INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
    INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
    INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
    PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
    PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
    PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
    PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
    PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
    PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
    PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
    PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
    PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
    PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
    PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
    PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
    PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
    PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
    PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
    PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
    EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
    EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
    EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
    EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
    EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
    EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
    EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
    EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
    EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
    EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
    EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
    EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
    EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
    EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
    EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
    EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
    EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
    EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
    EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
    EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
    EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
    EBX_REG_31__SCAN_IN, REIP_REG_1__SCAN_IN, REIP_REG_2__SCAN_IN,
    REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, REIP_REG_5__SCAN_IN,
    REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, REIP_REG_8__SCAN_IN,
    REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, REIP_REG_11__SCAN_IN,
    REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, REIP_REG_14__SCAN_IN,
    REIP_REG_15__SCAN_IN;
  output U2796;
  wire n10876, n10266, n8188, n7996, n6669, n8181, n8182, n12441, n6287,
    n6408, n6449, n8933, n9821, n6283, n6921, n10219, n7377, n6614, n6284,
    n6692, n7068, n6725, n6393, n6942, n8314, n7220, n8715, n9736, n6404,
    n6285, n9757, n6407, n12290, n12494, n12492, n7092, n10035, n8734,
    n10788, n10656, n8434, n8671, n6528, n9476, n8429, n6759, n8042, n7484,
    n9580, n12493, n11747, n8426, n7510, n8814, n9916, n9564, n9915, n7132,
    n8337, n8273, n7264, n9838, n9467, n7087, n9870, n7053, n9772, n6938,
    n6878, n7117, n6868, n8430, n8445, n8669, n8410, n8711, n8690, n6615,
    n6758, n6612, n6688, n6291, n6290, n6293, n6294, n8222, n6751, n6297,
    n6302, n6299, n6301, n6298, n6300, n6651, n6288, n6403, n6377, n8797,
    n7589, n8377, n6417, n6292, n6295, n6296, n6850, n6749, n6961, n6939,
    n6661, n6303, n8758, n6763, n7593, n8178, n7265, n7208, n6324, n7507,
    n6344, n6345, n6770, n8322, n7255, n8443, n6835, n7260, n7050, n6654,
    n6683, n6602, n6341, n8114, n6346, n10074, n7315, n7090, n7005, n6932,
    n8791, n12107, n6843, n7110, n6351, n6352, n8820, n8795, n11899, n8554,
    n7801, n8219, n8212, n6325, n8230, n6810, n6772, n8202, n8416, n7051,
    n7086, n9787, n7958, n6623, n6398, n7266, n6821, n7252, n6877, n6872,
    n8414, n8575, n6354, n6355, n8027, n8941, n7836, n11876, n6348, n6349,
    n6350, n7581, n7511, n10073, n7317, n7262, n8378, n8282, n6481, n11362,
    n6334, n8759, n7601, n8716, n6689, n6667, n8622, n6353, n12130, n8879,
    n12252, n7272, n11664, n7256, n7214, n10875, n12256, n7099, n8030,
    n8847, n6339, n6340, n7875, n7796, n7681, n7502, n7394, n7391, n11647,
    n6336, n11077, n7088, n9623, n8712, n6418, n11513, n10732, n10995,
    n9809, n9591, n11908, U2796_Lock, n6356, n8719, n8169, n6304, n6305,
    n6308, n7235, n6974, n6658, n8138, n6310, n6312, n6934, n6314, n6316,
    n7580, n8260, n6376, n9767, n9734, n7316, n8233, n10888, n6709, n6437,
    n6585, n6472, n6941, n7017, n7151, n7243, n7320, n7763, n6857, n7169,
    n6648, n8729, n6933, n6335, n7093, n7105, n6337, n6342, n6347, n6357,
    n7106, n7089, n9837, n6613, n6935, n8376, n7509, n6359, n6367, n6370,
    n6373, n8137, n6840, n6768, n8078, n8118, n8242, n6845, n6776, n6782,
    n6771, n7168, n6380, n6881, n6397, n6730, n7009, n7219, n8345, n7102,
    n6659, n7046, n7211, n6607, n6525, n6775, n7104, n7122, n8253, n8392,
    n8550, n6842, n9788, n6851, n8555, n8633, n11183, n8576, n8208, n7939,
    n7674, n11648, n9779, n8668, n12150, n12129, n12156, n8115, n7946,
    n7639, n7463, n7308, n9572, n8840, n11954, n10821, n11533, n9270,
    n9288, n8654, n12444, n9600, n10122, n10580, n8818, n9025, n12237,
    n8628, n10866, n6379, n6378, n6384, n6382, n6682, n8238, n6381, n6383,
    n6389, n6387, n6385, n6673, n8239, n6386, n6388, n6391, n6390, n6416,
    n6392, n6668, n6395, n6394, n6396, n6402, n6400, n6399, n6401, n6414,
    n6406, n6674, n6456, n6405, n6412, n6679, n6425, n7024, n6410, n6409,
    n6411, n6413, n6415, n6420, n6419, n6424, n6422, n8119, n6421, n6423,
    n6433, n8122, n6427, n6426, n6431, n6429, n6428, n6430, n6432, n6435,
    n6434, n6439, n6436, n6438, n6447, n6441, n6440, n6445, n6443, n6442,
    n6444, n6446, n6448, n9995, n6451, n6450, n6455, n6453, n6452, n6454,
    n6464, n6458, n6457, n6462, n6460, n6459, n6461, n6463, n6480, n8162,
    n6466, n6465, n6470, n6468, n6467, n6469, n6478, n6471, n6476, n6474,
    n6473, n6475, n6477, n6479, n8441, n6529, n6523, n10181, n6483, n6482,
    n8424, n6485, n6484, n6486, n9001, n6488, n6487, n6489, n12085, n6491,
    n6490, n6492, n8967, n6494, n6547, n6493, n6495, n8864, n6497, n6496,
    n6498, n11955, n6500, n6499, n6501, n8985, n6503, n6502, n6504, n10822,
    n6506, n6505, n6507, n10500, n6509, n6508, n6510, n10238, n6512, n6511,
    n6513, n11109, n6515, n6514, n6516, n11415, n6518, n6517, n6519,
    n10114, n6521, n6520, n6522, n9716, n6526, n6524, n6527, n6532, n6534,
    n10184, n6531, n6530, n10183, n10949, n6533, n9715, n6536, n6535,
    n6537, n10579, n10113, n6539, n6538, n6540, n10655, n11414, n6542,
    n6541, n6543, n10787, n11108, n6545, n6544, n6546, n10121, n10237,
    n10343, n6549, n6548, n6550, n10342, n10499, n10828, n6552, n6551,
    n6553, n10827, n8899, n6555, n6554, n6556, n8898, n8984, n11935, n6558,
    n6557, n6559, n11934, n11918, n6561, n6560, n6562, n11917, n8863,
    n6564, n6563, n6565, n8839, n8966, n6567, n6566, n6568, n8932, n12084,
    n8511, n6570, n6569, n6571, n8510, n9000, n12172, n6573, n6572, n6574,
    n12171, n8603, n6576, n6575, n6577, n8604, n6579, n6578, n6580, n12289,
    n8423, n8425, n7951, n6584, n6589, n6587, n6586, n6588, n6597, n6591,
    n6590, n6595, n6593, n6592, n6594, n6596, n6599, n6598, n6604, n6600,
    n6601, n6603, n6605, n6606, n6611, n6609, n6608, n6610, n9581, n7686,
    n6619, n6617, n6616, n6618, n6621, n6620, n6639, n6622, n6627, n6625,
    n6624, n6626, n6637, n6630, n6628, n6629, n6635, n6633, n6631, n6632,
    n6634, n6636, n6638, n6647, n6641, n6640, n6645, n6643, n6642, n6644,
    n6646, n10380, n6844, n6650, n6649, n6656, n6652, n6653, n6655, n6660,
    n6657, n6665, n6663, n6662, n6664, n6666, n6691, n6671, n6670, n6678,
    n6672, n6676, n6675, n6677, n6681, n6680, n6687, n6685, n6684, n6686,
    n6690, n6694, n6693, n6698, n6696, n6695, n6697, n6707, n6700, n6699,
    n6705, n6703, n6701, n6702, n6704, n6706, n6724, n6708, n6714, n6710,
    n6712, n6711, n6713, n6722, n6716, n6715, n6720, n6718, n6717, n6719,
    n6721, n6723, n6727, n6726, n6732, n6728, n6729, n6731, n6740, n6734,
    n6733, n6738, n6736, n6735, n6737, n6739, n6742, n6741, n6746, n6744,
    n6743, n6745, n6756, n6748, n6747, n6754, n6752, n6750, n6753, n6755,
    n6757, n6808, n9589, n6766, n6764, n6765, n6767, n6769, n6777, n6773,
    n6774, n6820, n8290, n6811, n6780, n8388, n6797, n6778, n6795, n6779,
    n6807, n6781, n6784, n8390, n6783, n6802, n6786, n6785, n6803, n6794,
    n6789, n6787, n6792, n6788, n6790, n6791, n6793, n6801, n6799, n6796,
    n6798, n6800, n6805, n6804, n6806, n6813, n6809, n6814, n8387, n6812,
    n6818, n6816, n6815, n6817, n6819, n6823, n6822, n7588, n6827, n6829,
    n7133, n11806, n6828, n6831, n7112, n6830, n6833, n7751, n6832, n7091,
    n6834, n6853, n6836, n7602, n6837, n6839, n6838, n7591, n6848, n6841,
    n6864, n6846, n8399, n6858, n6847, n6849, n6855, n8577, n8398, n8386,
    n6852, n6854, n6880, n6856, n6892, n6860, n6859, n6862, n9472, n6861,
    n7596, n11900, n6863, n6865, n6866, n6867, n6869, n6873, n6893, n6871,
    n8457, n8487, n6870, n7115, n6937, n6876, n8763, n6874, n11283, n6875,
    n6936, n6882, n8565, n6879, n6883, n6885, n6884, n7113, n6888, n10039,
    n10029, n6896, n6886, n10153, n6887, n6890, n6889, n6891, n6895, n6894,
    n6898, n10731, n6897, n6900, n6899, n6904, n6902, n6901, n6903, n6912,
    n6906, n6905, n6910, n6908, n6907, n6909, n6911, n6929, n6914, n6913,
    n6918, n6916, n6915, n6917, n6927, n6920, n6919, n6925, n6923, n6922,
    n6924, n6926, n6928, n8306, n6931, n6930, n10956, n7006, n6940, n6946,
    n6944, n6943, n6945, n6954, n6948, n6947, n6952, n6950, n6949, n6951,
    n6953, n6971, n6956, n6955, n6960, n6958, n6957, n6959, n6969, n6963,
    n6962, n6967, n6965, n6964, n6966, n6968, n6970, n6973, n6972, n7007,
    n8187, n6976, n6975, n6980, n6978, n6977, n6979, n7004, n6982, n6981,
    n6984, n6983, n6986, n6985, n7002, n6988, n6987, n6992, n6990, n6989,
    n6991, n7000, n6994, n6993, n6998, n6996, n6995, n6997, n6999, n7001,
    n7003, n8292, n8276, n7008, n7042, n7011, n7010, n7015, n7013, n7012,
    n7014, n7040, n7016, n7019, n7018, n7021, n7020, n7038, n7023, n7022,
    n7028, n7026, n7025, n7027, n7036, n7030, n7029, n7034, n7032, n7031,
    n7033, n7035, n7037, n7039, n8291, n7041, n7044, n7048, n7043, n7045,
    n7123, n7047, n7125, n7049, n8272, n7103, n7052, n9889, n7055, n7054,
    n7059, n7057, n7056, n7058, n7067, n7061, n7060, n7065, n7063, n7062,
    n7064, n7066, n7084, n7070, n7069, n7074, n7072, n7071, n7073, n7082,
    n7076, n7075, n7080, n7078, n7077, n7079, n7081, n7083, n8299, n7085,
    n7094, n7177, n9557, n7095, n7100, n11508, n7096, n7098, n7097, n7173,
    n7101, n7130, n9573, n9737, n7111, n7108, n7107, n7109, n7119, n7114,
    n7116, n11167, n7118, n7121, n7120, n9446, n7129, n7124, n7126, n9444,
    n9455, n7127, n7128, n9448, n9466, n7131, n9558, n7135, n11793, n10891,
    n7134, n7172, n7170, n7167, n7137, n7136, n7141, n7139, n7138, n7140,
    n7165, n7143, n7142, n7145, n7144, n7147, n7146, n7163, n7149, n7148,
    n7153, n7150, n7152, n7161, n7155, n7154, n7159, n7157, n7156, n7158,
    n7160, n7162, n7164, n8311, n7166, n7176, n7171, n7175, n7174, n9563,
    n9601, n7213, n7179, n7178, n7183, n7181, n7180, n7182, n7191, n7185,
    n7184, n7189, n7187, n7186, n7188, n7190, n7207, n7193, n7192, n7197,
    n7195, n7194, n7196, n7205, n7199, n7198, n7203, n7201, n7200, n7202,
    n7204, n7206, n8324, n7210, n7209, n7212, n7218, n7216, n11867, n7215,
    n7217, n7254, n7222, n7221, n7226, n7224, n7223, n7225, n7251, n7228,
    n7227, n7230, n7229, n7232, n7231, n7249, n7234, n7233, n7239, n8229,
    n7237, n7236, n7238, n7247, n7241, n7240, n7245, n7242, n7244, n7246,
    n7248, n7250, n8334, n7253, n7263, n7258, n11677, n7257, n7259, n7261,
    n7271, n7268, n7267, n7269, n7270, n7276, n7274, n11641, n7273, n7275,
    n9917, n10081, n7278, n7277, n7282, n7280, n7279, n7281, n7290, n7284,
    n7283, n7288, n7286, n7285, n7287, n7289, n7306, n7292, n7291, n7296,
    n7294, n7293, n7295, n7304, n7298, n7297, n7302, n7300, n7299, n7301,
    n7303, n7305, n7307, n7312, n7310, n11850, n7309, n7311, n7314, n7313,
    n10082, n7319, n11604, n7318, n7354, n7321, n7323, n7322, n7325, n7324,
    n7341, n7327, n7326, n7331, n7329, n7328, n7330, n7339, n7333, n7332,
    n7337, n7335, n7334, n7336, n7338, n7340, n7349, n7343, n7342, n7347,
    n7345, n7344, n7346, n7348, n7350, n7352, n7351, n7353, n10240, n7356,
    n7355, n7360, n7358, n7357, n7359, n7368, n7362, n7361, n7366, n7364,
    n7363, n7365, n7367, n7385, n7370, n7369, n7374, n7372, n7371, n7373,
    n7383, n7376, n7375, n7381, n7379, n7378, n7380, n7382, n7384, n7386,
    n7390, n7388, n7387, n7389, n7393, n11658, n7392, n10239, n7396,
    n11691, n7395, n7431, n7429, n7398, n7397, n7400, n8041, n7399, n7402,
    n7401, n7418, n7404, n7403, n7408, n7406, n7405, n7407, n7416, n7410,
    n7409, n7414, n7412, n7411, n7413, n7415, n7417, n7426, n7420, n7419,
    n7424, n7422, n7421, n7423, n7425, n7427, n7428, n7430, n10277, n7433,
    n7432, n7437, n7435, n7434, n7436, n7445, n7439, n7438, n7443, n7441,
    n7440, n7442, n7444, n7461, n7447, n7446, n7451, n7449, n7448, n7450,
    n7459, n7453, n7452, n7457, n7455, n7454, n7456, n7458, n7460, n7462,
    n7467, n7465, n11967, n7464, n7466, n7469, n7468, n10501, n7471, n7470,
    n7473, n7472, n7475, n7474, n7492, n7477, n7476, n7481, n7479, n7478,
    n7480, n7490, n7483, n7482, n7488, n7486, n7485, n7487, n7489, n7491,
    n7500, n7494, n7493, n7498, n7496, n7495, n7497, n7499, n7501, n7508,
    n11155, n7506, n7504, n7503, n7505, n8815, n7513, n11818, n7512, n7548,
    n7515, n7514, n7517, n7516, n7519, n7518, n7535, n7521, n7520, n7525,
    n7523, n7522, n7524, n7533, n7527, n7526, n7531, n7529, n7528, n7530,
    n7532, n7534, n7543, n7537, n7536, n7541, n7539, n7538, n7540, n7542,
    n7544, n7546, n7545, n7547, n8821, n7550, n7549, n7554, n7552, n7551,
    n7553, n7562, n7556, n7555, n7560, n7558, n7557, n7559, n7561, n7578,
    n7564, n7563, n7568, n7566, n7565, n7567, n7576, n7570, n7569, n7574,
    n7572, n7571, n7573, n7575, n7577, n7579, n7585, n7583, n12045, n7582,
    n7584, n7587, n7586, n11254, n7638, n7600, n7590, n7592, n10867, n7599,
    n7594, n7595, n8383, n7597, n7598, n8438, n7604, n7603, n7608, n7606,
    n7605, n7607, n7616, n7610, n7609, n7614, n7612, n7611, n7613, n7615,
    n7632, n7618, n7617, n7622, n7620, n7619, n7621, n7630, n7624, n7623,
    n7628, n7626, n7625, n7627, n7629, n7631, n7633, n7636, n7634, n7635,
    n7637, n7641, n12075, n7640, n11699, n7643, n7642, n7647, n7645, n7644,
    n7646, n7655, n7649, n7648, n7653, n7651, n7650, n7652, n7654, n7671,
    n7657, n7656, n7661, n7659, n7658, n7660, n7669, n7663, n7662, n7667,
    n7665, n7664, n7666, n7668, n7670, n7672, n7678, n7676, n7673, n12095,
    n7675, n7677, n7680, n7679, n11746, n11875, n7683, n7757, n12177,
    n7682, n7719, n7717, n7685, n7684, n7688, n7687, n7690, n7689, n7706,
    n7692, n7691, n7696, n7694, n7693, n7695, n7704, n7698, n7697, n7702,
    n7700, n7699, n7701, n7703, n7705, n7714, n7708, n7707, n7712, n7710,
    n7709, n7711, n7713, n7715, n7716, n7718, n11914, n7721, n7720, n7723,
    n7722, n7725, n7724, n7741, n7727, n7726, n7731, n7729, n7728, n7730,
    n7739, n7733, n7732, n7737, n7735, n7734, n7736, n7738, n7740, n7749,
    n7743, n7742, n7747, n7745, n7744, n7746, n7748, n7750, n7753, n7752,
    n7756, n7754, n7755, n7759, n11940, n12118, n7758, n11913, n7795,
    n7761, n7760, n7765, n7762, n7764, n7773, n7767, n7766, n7771, n7769,
    n7768, n7770, n7772, n7789, n7775, n7774, n7779, n7777, n7776, n7778,
    n7787, n7781, n7780, n7785, n7783, n7782, n7784, n7786, n7788, n7790,
    n7793, n7791, n7792, n7794, n7798, n12272, n7797, n8862, n7800, n7799,
    n7803, n7802, n7805, n7804, n7821, n7807, n7806, n7811, n7809, n7808,
    n7810, n7819, n7813, n7812, n7817, n7815, n7814, n7816, n7818, n7820,
    n7829, n7823, n7822, n7827, n7825, n7824, n7826, n7828, n7830, n7832,
    n7831, n7835, n7833, n7834, n7838, n12340, n7837, n8834, n7874, n7840,
    n7839, n7844, n7842, n7841, n7843, n7852, n7846, n7845, n7850, n7848,
    n7847, n7849, n7851, n7868, n7854, n7853, n7858, n7856, n7855, n7857,
    n7866, n7860, n7859, n7864, n7862, n7861, n7863, n7865, n7867, n7869,
    n7872, n7870, n7871, n7873, n7877, n12359, n7876, n8848, n7879, n7878,
    n7883, n7881, n7880, n7882, n7891, n7885, n7884, n7889, n7887, n7886,
    n7888, n7890, n7907, n7893, n7892, n7897, n7895, n7894, n7896, n7905,
    n7899, n7898, n7903, n7901, n7900, n7902, n7904, n7906, n7981, n7909,
    n7908, n7913, n7911, n7910, n7912, n7921, n7915, n7914, n7919, n7917,
    n7916, n7918, n7920, n7937, n7923, n7922, n7927, n7925, n7924, n7926,
    n7935, n7929, n7928, n7933, n7931, n7930, n7932, n7934, n7936, n7982,
    n7938, n7943, n7941, n12420, n7940, n7942, n7945, n7944, n8878, n8940,
    n7948, n12457, n7947, n7987, n7950, n7949, n7955, n7953, n7952, n7954,
    n7980, n7957, n7956, n7960, n7959, n7962, n7961, n7978, n7964, n7963,
    n7968, n7966, n7965, n7967, n7976, n7970, n7969, n7974, n7972, n7971,
    n7973, n7975, n7977, n7979, n8019, n8020, n7983, n7985, n7984, n7986,
    n8522, n7989, n7988, n7993, n7991, n7990, n7992, n8002, n7995, n7994,
    n8000, n7998, n7997, n7999, n8001, n8018, n8004, n8003, n8008, n8006,
    n8005, n8007, n8016, n8010, n8009, n8014, n8012, n8011, n8013, n8015,
    n8017, n8066, n8065, n8021, n8023, n8022, n8026, n8024, n8025, n8029,
    n12128, n12147, n8028, n8523, n8032, n8111, n12353, n8031, n8071,
    n8034, n8033, n8038, n8036, n8035, n8037, n8064, n8040, n8039, n8044,
    n8043, n8046, n8045, n8062, n8048, n8047, n8052, n8050, n8049, n8051,
    n8060, n8054, n8053, n8058, n8056, n8055, n8057, n8059, n8061, n8063,
    n8103, n8104, n8067, n8069, n8068, n8070, n8073, n8072, n8077, n8075,
    n8074, n8076, n8086, n8080, n8079, n8084, n8082, n8081, n8083, n8085,
    n8102, n8088, n8087, n8092, n8090, n8089, n8091, n8100, n8094, n8093,
    n8098, n8096, n8095, n8097, n8099, n8101, n8154, n8153, n8105, n8107,
    n8106, n8110, n8108, n8109, n8113, n12346, n12380, n8112, n12166,
    n8117, n12255, n12313, n8116, n8159, n8121, n8120, n8126, n8124, n8123,
    n8125, n8134, n8128, n8127, n8132, n8130, n8129, n8131, n8133, n8152,
    n8136, n8135, n8142, n8140, n8139, n8141, n8150, n8144, n8143, n8148,
    n8146, n8145, n8147, n8149, n8151, n8199, n8200, n8155, n8157, n8156,
    n8158, n8621, n8207, n8164, n8163, n8168, n8166, n8165, n8167, n8177,
    n8171, n8170, n8175, n8173, n8172, n8174, n8176, n8198, n8180, n8179,
    n8186, n8184, n8183, n8185, n8196, n8190, n8189, n8194, n8192, n8191,
    n8193, n8195, n8197, n8251, n8252, n8201, n8205, n8203, n8204, n8206,
    n8210, n8266, n12432, n8209, n8546, n8211, n8256, n8214, n8213, n8218,
    n8216, n8215, n8217, n8228, n8221, n8220, n8226, n8224, n8223, n8225,
    n8227, n8250, n8232, n8231, n8237, n8235, n8234, n8236, n8248, n8241,
    n8240, n8246, n8244, n8243, n8245, n8247, n8249, n8259, n8262, n8254,
    n8255, n8258, n8257, n8264, n8261, n8263, n8268, n8265, n8656, n8267,
    n8548, n8677, n8666, n8389, n8391, n8678, n8397, n8639, n8422, n8421,
    n8428, n8427, n11178, n9290, n8547, n8549, n8552, n8551, n8553, n8556,
    n9020, n8570, n8629, n11911, n8630, n9269, n9271, n9276, n9730, n8631,
    n8805, n8632, n8655, n8634, n9209, n12158, n8636, n12316, n8959,
    n11827, n11160, n8872, n11646, n11624, n11193, n8871, n10881, n10870,
    n8869, n9459, n11498, n10869, n11856, n8637, n11632, n11633, n11842,
    n9169, n11846, n8870, n11122, n11151, n11829, n11247, n11246, n11923,
    n8638, n11943, n8855, n8914, n8924, n9195, n12157, n12253, n8643,
    n8650, n8647, n12437, n9016, n8640, n9023, n8788, n8648, n8641, n12031,
    n11725, n12427, n8649, n8651, n12434, n9017, n9019, n9018, n9022,
    n9021, keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4,
    keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9,
    keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14,
    keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19,
    keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24,
    keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29,
    keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34,
    keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39,
    keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44,
    keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49,
    keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54,
    keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59,
    keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64,
    keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69,
    keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74,
    keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79,
    keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84,
    keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89,
    keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94,
    keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99,
    keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104,
    keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109,
    keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114,
    keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119,
    keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124,
    keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129,
    keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134,
    keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139,
    keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144,
    keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149,
    keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154,
    keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159,
    input_0, input_1, AND_1, input_2, OR_2, input_3, AND_3, input_4, OR_4,
    input_5, OR_5, input_6, AND_6, input_7, AND_7, input_8, OR_8, input_9,
    OR_9, input_10, OR_10, input_11, AND_11, input_12, OR_12, input_13,
    AND_13, input_14, AND_14, input_15, OR_15, input_16, AND_16, input_17,
    OR_17, input_18, OR_18, input_19, OR_19, input_20, OR_20, input_21,
    AND_21, input_22, OR_22, input_23, AND_23, input_24, AND_24, input_25,
    OR_25, input_26, OR_26, input_27, OR_27, input_28, OR_28, input_29,
    OR_29, input_30, AND_30, input_31, OR_31, input_32, OR_32, input_33,
    OR_33, input_34, OR_34, input_35, OR_35, input_36, AND_36, input_37,
    AND_37, input_38, OR_38, input_39, AND_39, input_40, OR_40, input_41,
    AND_41, input_42, OR_42, input_43, OR_43, input_44, OR_44, input_45,
    AND_45, input_46, OR_46, input_47, OR_47, input_48, OR_48, input_49,
    OR_49, input_50, AND_50, input_51, OR_51, input_52, OR_52, input_53,
    AND_53, input_54, OR_54, input_55, OR_55, input_56, OR_56, input_57,
    AND_57, input_58, OR_58, input_59, AND_59, input_60, AND_60, input_61,
    AND_61, input_62, AND_62, input_63, OR_63, input_64, AND_64, input_65,
    OR_65, input_66, OR_66, input_67, OR_67, input_68, AND_68, input_69,
    AND_69, input_70, AND_70, input_71, AND_71, input_72, OR_72, input_73,
    OR_73, input_74, OR_74, input_75, AND_75, input_76, OR_76, input_77,
    OR_77, input_78, OR_78, input_79, OR_79, input_80, input_81, AND_81,
    input_82, OR_82, input_83, AND_83, input_84, OR_84, input_85, OR_85,
    input_86, AND_86, input_87, AND_87, input_88, OR_88, input_89, OR_89,
    input_90, OR_90, input_91, AND_91, input_92, OR_92, input_93, AND_93,
    input_94, AND_94, input_95, OR_95, input_96, AND_96, input_97, OR_97,
    input_98, OR_98, input_99, OR_99, input_100, OR_100, input_101,
    AND_101, input_102, OR_102, input_103, AND_103, input_104, AND_104,
    input_105, OR_105, input_106, OR_106, input_107, OR_107, input_108,
    OR_108, input_109, OR_109, input_110, AND_110, input_111, OR_111,
    input_112, OR_112, input_113, OR_113, input_114, OR_114, input_115,
    OR_115, input_116, AND_116, input_117, AND_117, input_118, OR_118,
    input_119, AND_119, input_120, OR_120, input_121, AND_121, input_122,
    OR_122, input_123, OR_123, input_124, OR_124, input_125, AND_125,
    input_126, OR_126, input_127, OR_127, input_128, OR_128, input_129,
    OR_129, input_130, AND_130, input_131, OR_131, input_132, OR_132,
    input_133, AND_133, input_134, OR_134, input_135, OR_135, input_136,
    OR_136, input_137, AND_137, input_138, OR_138, input_139, AND_139,
    input_140, AND_140, input_141, AND_141, input_142, AND_142, input_143,
    OR_143, input_144, AND_144, input_145, OR_145, input_146, OR_146,
    input_147, OR_147, input_148, AND_148, input_149, AND_149, input_150,
    AND_150, input_151, AND_151, input_152, OR_152, input_153, OR_153,
    input_154, OR_154, input_155, AND_155, input_156, OR_156, input_157,
    OR_157, input_158, OR_158, input_159, OR_159, OR_159_INV, CASOP;
  assign n10876 = ~n8671;
  assign n10266 = ~n12492;
  assign n8188 = ~n6456;
  assign n7996 = ~n6692;
  assign n6669 = ~n6393 & ~n6408;
  assign n8181 = ~n6692;
  assign n8182 = ~n7068;
  assign n12441 = ~n11725 & ~n10888;
  assign n6287 = ~n6961;
  assign n6408 = ~n6377 | ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n6449 = ~n6433 | ~n6432;
  assign n8933 = ~n8967 & ~n8966;
  assign n9821 = ~n8441;
  assign n6283 = n6403 | n6407;
  assign n6921 = n9580 | n6404;
  assign n10219 = n6691 | n6690;
  assign n7377 = n6393 | n8758;
  assign n6614 = ~n6613 | ~n6612;
  assign n6284 = ~n6692;
  assign n6692 = n6404 | n6403;
  assign n7068 = ~n6668;
  assign n6725 = ~n6456;
  assign n6393 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n6376;
  assign n6942 = ~n6661;
  assign n8314 = n7220 ^ ~n7211;
  assign n7220 = ~n7177 | ~n7176;
  assign n8715 = ~n9736;
  assign n9736 = n6724 | n6723;
  assign n6404 = ~n6380 | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n6285 = ~n6393 & ~n6408;
  assign n9757 = ~n6418 | ~n6417;
  assign n6407 = INSTQUEUERD_ADDR_REG_3__SCAN_IN | INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n12290 = ~n8603 & ~n8604;
  assign n12494 = ~n12492 & ~n6850;
  assign n12492 = ~n6615 & ~n6614;
  assign n7092 = n7087 | n7086;
  assign n10035 = n6933 & n6932;
  assign n8734 = ~n9889 | ~n7053;
  assign n10788 = ~n11415 & ~n11414;
  assign n10656 = ~n10114 & ~n10113;
  assign n8434 = ~n6528;
  assign n8671 = ~n9476 | ~n8441;
  assign n6528 = ~n6842;
  assign n9476 = ~n9757;
  assign n8429 = ~n10219;
  assign n6759 = ~n6850;
  assign n8042 = ~n6682;
  assign n7484 = ~n7377;
  assign n9580 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n12493 = n8554 ^ ~n8553;
  assign n11747 = ~n8820 & ~n6348;
  assign n8426 = n8424 | n8423;
  assign n7510 = ~n8814 & ~n8815;
  assign n8814 = n7507 ^ ~n7508;
  assign n9916 = ~n9601 & ~n9600;
  assign n9564 = ~n9557 & ~n9558;
  assign n9915 = ~n7262 | ~n7261;
  assign n7132 = ~n9573 & ~n9572;
  assign n8337 = n8273 ^ ~n7269;
  assign n8273 = ~n7264 | ~n7263;
  assign n7264 = ~n7220 & ~n7219;
  assign n9838 = n7093 | n7092;
  assign n9467 = ~n7111 | ~n7110;
  assign n7087 = ~n8734 & ~STATE2_REG_0__SCAN_IN;
  assign n9870 = n7053 ^ ~n6334;
  assign n7053 = ~n6891 | ~n7050;
  assign n9772 = ~n6898 & ~n6897;
  assign n6938 = n6936 ^ ~n6935;
  assign n6878 = ~n6892 | ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7117 = n6868 & n6867;
  assign n6868 = n6862 & n7596;
  assign n8430 = ~n8576 & ~n6879;
  assign n8445 = ~n6853 & ~n9995;
  assign n8669 = n8416 & n6851;
  assign n8410 = ~n9476 & ~n6296;
  assign n8711 = ~n8576 & ~n6842;
  assign n8690 = ~n10380;
  assign n6615 = ~n6597 | ~n6596;
  assign n6758 = ~n6740 | ~n6739;
  assign n6612 = ~n6611 & ~n6610;
  assign n6688 = ~n6687 & ~n6686;
  assign n6291 = ~n6290;
  assign n6290 = ~n8230;
  assign n6293 = ~n6283;
  assign n6294 = ~n6283;
  assign n8222 = ~n6658;
  assign n6751 = n6750 | n7068;
  assign n6297 = ~n7377;
  assign n6302 = ~n6921;
  assign n6299 = ~n6921;
  assign n6301 = ~n6921;
  assign n6298 = ~n7377;
  assign n6300 = ~n6921;
  assign n6651 = ~n6395 | ~n6394;
  assign n6288 = ~n6283;
  assign n6403 = ~n8729 | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n6377 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n8797 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n7589 = ~n8429 | ~n9736;
  assign n8377 = ~n8414 & ~n12492;
  assign n6417 = ~n6416 & ~n6415;
  assign n6292 = ~n6290;
  assign n6295 = ~n6283;
  assign n6296 = ~n6480 & ~n6479;
  assign n6850 = ~n6758 & ~n6757;
  assign n6749 = ~n9580 & ~n6393;
  assign n6961 = ~n6749;
  assign n6939 = ~n10956;
  assign n6661 = ~n8758 & ~n6407;
  assign n6303 = ~n6961;
  assign n8758 = ~n8729 | ~n6763;
  assign n6763 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n7593 = n6850 & n9736;
  assign n8178 = ~n6942;
  assign n7265 = ~n7208;
  assign n7208 = ~STATE2_REG_0__SCAN_IN | ~n7009;
  assign n6324 = ~n7591 & ~n6759;
  assign n7507 = ~n10240 | ~n6344;
  assign n6344 = ~n6346 & ~n6345;
  assign n6345 = ~n10501;
  assign n6770 = ~n6769 | ~n6768;
  assign n8322 = n7264 ^ ~n7255;
  assign n7255 = ~n7263;
  assign n8443 = ~n10219 | ~n6850;
  assign n6835 = ~n8715 | ~n6759;
  assign n7260 = n8322 & n8260;
  assign n7050 = ~n6885 | ~n6884;
  assign n6654 = n6652 | n6651;
  assign n6683 = ~n8797 & ~n6408;
  assign n6602 = n6600 | n7068;
  assign n6341 = ~n6342 | ~n11913;
  assign n8114 = ~n6827;
  assign n6346 = ~n10239 | ~n6347;
  assign n10074 = ~n7316 | ~n7315;
  assign n7315 = n10081 & n10082;
  assign n7090 = n11077 & n8260;
  assign n7005 = ~n7007 & ~n6367;
  assign n6932 = n6931 & n6930;
  assign n8791 = ~n6823 | ~n6822;
  assign n12107 = ~n8071 & ~n8070;
  assign n6843 = ~n6449 & ~n6448;
  assign n7110 = ~n6370 & ~n7109;
  assign n6351 = ~n11254 | ~n6352;
  assign n6352 = ~n8821;
  assign n8820 = ~n7510 & ~n7509;
  assign n8795 = ~STATE2_REG_1__SCAN_IN & ~n10732;
  assign n11899 = ~n9581;
  assign n8554 = n8622 | n8549;
  assign n7801 = ~n8222;
  assign n8219 = ~n6651;
  assign n8212 = ~n6456;
  assign n6325 = n7177 ^ ~n7168;
  assign n8230 = ~n6692;
  assign n6810 = ~n6772 & ~n6771;
  assign n6772 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~n6770;
  assign n8202 = ~n8253;
  assign n8416 = ~n8399 & ~n8441;
  assign n7051 = n6890 & n6889;
  assign n7086 = n7085 | n6359;
  assign n9787 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n7958 = ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n6623 = ~n6288 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n6398 = ~n8797;
  assign n7266 = ~n7252;
  assign n6821 = ~n8290 & ~n7208;
  assign n7252 = ~n7009 & ~n9734;
  assign n6877 = ~n6876 & ~n6875;
  assign n6872 = ~n7115;
  assign n8414 = ~n6835;
  assign n8575 = ~n7593;
  assign n6354 = ~n12107 & ~n6355;
  assign n6355 = ~n8523;
  assign n8027 = ~n7946 | ~PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n8941 = ~n7987 & ~n7986;
  assign n7836 = n7796 & PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n11876 = ~n7719 & ~n7718;
  assign n6348 = ~n6350 | ~n6349;
  assign n6349 = ~n6351;
  assign n6350 = ~n11699;
  assign n7581 = ~n7511 | ~PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n7511 = ~n7502 & ~n11183;
  assign n10073 = ~n7354 & ~n7353;
  assign n7317 = ~n7308 | ~PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n7262 = ~n7260 & ~n7259;
  assign n8378 = ~n6843 & ~n10380;
  assign n8282 = ~n8291;
  assign n6481 = ~n6523;
  assign n11362 = ~STATEBS16_REG_SCAN_IN;
  assign n6334 = ~n9772;
  assign n8759 = ~n7602 | ~n7601;
  assign n7601 = ~n7600 & ~n8438;
  assign n8716 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n6689 = ~n6678 & ~n6677;
  assign n6667 = ~n6656 & ~n6655;
  assign n8622 = ~n8522 | ~n6353;
  assign n6353 = n12166 & n6354;
  assign n12130 = ~n8924 & ~n9195;
  assign n8879 = ~n8847 & ~n8848;
  assign n12252 = ~n10888 & ~n12129;
  assign n7272 = ~n7256 | ~PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n11664 = ~PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n7256 = ~n7214 & ~n9809;
  assign n7214 = n11793 | n7133;
  assign n10875 = ~n10732 & ~n10888;
  assign n12256 = ~n12441;
  assign n7099 = ~n6308 & ~n6316;
  assign n8030 = ~n8027 & ~n12128;
  assign n8847 = ~n11914 | ~n6339;
  assign n6339 = ~n6341 & ~n6340;
  assign n6340 = ~n8834;
  assign n7875 = n7836 & PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n7796 = ~n7757 & ~n11940;
  assign n7681 = ~n7674 & ~n7673;
  assign n7502 = ~n7463 | ~PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n7394 = ~n7391 | ~PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n7391 = ~n7317 & ~n10995;
  assign n11647 = STATE2_REG_2__SCAN_IN | n8457;
  assign n6336 = ~n7102;
  assign n11077 = n7089 & n7088;
  assign n7088 = ~n9837;
  assign n9623 = ~STATE2_REG_1__SCAN_IN & ~STATE2_REG_3__SCAN_IN;
  assign n8712 = ~n10876 | ~n8445;
  assign n6418 = ~n6384 & ~n6383;
  assign n11513 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n10732 = ~STATE2_REG_2__SCAN_IN;
  assign n10995 = ~PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n9809 = ~PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n9591 = ~n6376;
  assign n11908 = ~STATE2_REG_1__SCAN_IN;
  assign U2796_Lock = ~n6357 | ~n6305;
  assign n6356 = ~n6304 & ~n6310;
  assign n8719 = ~n6683;
  assign n8169 = ~n8719;
  assign n6304 = n9022 | n9021;
  assign n6305 = n6312 & n6356;
  assign n6308 = ~n7098 | ~n7097;
  assign n7235 = ~n6669;
  assign n6974 = ~n6648;
  assign n6658 = ~n6394 | ~n6398;
  assign n8138 = ~n7801;
  assign n6310 = REIP_REG_31__SCAN_IN & n9023;
  assign n6312 = n11178 | n12444;
  assign n6934 = ~n9734 & ~n6881;
  assign n6314 = n7102 | n7103;
  assign n6316 = n7173 & n9591;
  assign n7580 = ~n8260;
  assign n8260 = ~n10732 & ~n6759;
  assign n6376 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n9767 = ~n7094 | ~n9838;
  assign n9734 = ~STATE2_REG_0__SCAN_IN;
  assign n7316 = n9916 & n9915;
  assign n8233 = ~n7377;
  assign n10888 = ~n8633 & ~n8632;
  assign n6709 = ~n6295 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n6437 = ~n6294 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n6585 = ~n6295 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n6472 = ~n6293 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n6941 = ~n6294 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n7017 = ~n6288 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n7151 = ~n6294 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n7243 = ~n6288 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n7320 = ~n6293 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n7763 = ~n6288 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n6857 = ~n6335 & ~n6324;
  assign n7169 = ~n6325 | ~n8260;
  assign n6648 = ~n8758 & ~n6404;
  assign n8729 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n6933 = ~n9870 | ~n9734;
  assign n6335 = ~n6838 | ~n6839;
  assign n7093 = n6337 & n6314;
  assign n7105 = ~n6337 | ~n6336;
  assign n6337 = ~n7006 | ~n7005;
  assign n6342 = ~n8862;
  assign n6347 = ~n10277;
  assign n6357 = ~n12493 | ~n12237;
  assign n7106 = ~n9737;
  assign n7089 = ~n7177;
  assign n9837 = n10035 & n7094;
  assign n6613 = ~n6604 & ~n6603;
  assign n6935 = ~n6934;
  assign n8376 = ~n7588 | ~n10266;
  assign n7509 = ~n7508 & ~n7507;
  assign n6359 = n7265 & INSTQUEUE_REG_0__2__SCAN_IN;
  assign n6367 = n7252 & n8292;
  assign n6370 = n7751 & EAX_REG_1__SCAN_IN;
  assign n6373 = ~n8548 | ~n8547;
  assign n8137 = ~n7068;
  assign n6840 = n8429 ^ ~n7593;
  assign n6768 = ~n6777 | ~n9787;
  assign n8078 = ~n6942;
  assign n8118 = ~n8042;
  assign n8242 = ~n6425;
  assign n6845 = ~n8416;
  assign n6776 = n8716 ^ n6770;
  assign n6782 = INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ ~n6764;
  assign n6771 = ~n6776 & ~n11533;
  assign n7168 = ~n7176;
  assign n6380 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n6881 = ~n8430 & ~n6880;
  assign n6397 = n6392 | n7068;
  assign n6730 = n6728 | n7377;
  assign n7009 = ~n8441 & ~n8429;
  assign n7219 = ~n7210 & ~n7209;
  assign n8345 = ~n6971 & ~n6970;
  assign n7102 = ~n8276 & ~n7008;
  assign n6659 = n6658 | n6657;
  assign n7046 = ~n9734 & ~n10219;
  assign n7211 = ~n7219;
  assign n6607 = n8042 | n6605;
  assign n6525 = n6524 | n8410;
  assign n6775 = ~n6810 & ~n6774;
  assign n7104 = ~n7103;
  assign n7122 = ~n7044 & ~n7043;
  assign n8253 = ~n9734 & ~n8759;
  assign n8392 = ~n6808 & ~n6775;
  assign n8550 = ~STATE2_REG_2__SCAN_IN & ~n11362;
  assign n6842 = ~n9757 | ~n9995;
  assign n9788 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n6851 = ~n8398;
  assign n8555 = ~n8266 & ~n8265;
  assign n8633 = ~n11911 | ~n9288;
  assign n11183 = ~PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n8576 = ~n12494;
  assign n8208 = ~n8115 & ~n12255;
  assign n7939 = n7875 & PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n7674 = ~n7639 | ~PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n11648 = ~PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n9779 = ~n7125 & ~n7124;
  assign n8668 = ~n8570 & ~n8677;
  assign n12150 = ~n12129;
  assign n12129 = ~n8650 & ~n8647;
  assign n12156 = ~n12252;
  assign n8115 = n8111 | n12346;
  assign n7946 = n7939 & PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n7639 = ~n7581 & ~n8818;
  assign n7463 = ~n7394 & ~n11648;
  assign n7308 = ~n7272 & ~n11664;
  assign n9572 = ~n9467 | ~n9466;
  assign n8840 = ~n8864 & ~n8863;
  assign n11954 = ~n11935 | ~n11934;
  assign n10821 = ~n10828 | ~n10827;
  assign n11533 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n9270 = ~n8791;
  assign n9288 = ~n8630 | ~n9276;
  assign n8654 = PHYADDRPOINTER_REG_31__SCAN_IN ^ n8556;
  assign n12444 = ~n12031;
  assign n9600 = ~n7218 & ~n7217;
  assign n10122 = ~n11109 & ~n11108;
  assign n10580 = ~n9716 & ~n9715;
  assign n8818 = ~PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n9025 = STATE2_REG_2__SCAN_IN | STATEBS16_REG_SCAN_IN;
  assign n12237 = ~n8654 & ~n8634;
  assign n8628 = ~n9025;
  assign n10866 = ~INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n6379 = ~n6294 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n6378 = ~n6285 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n6384 = ~n6379 | ~n6378;
  assign n6382 = ~INSTQUEUE_REG_4__1__SCAN_IN | ~n6648;
  assign n6682 = ~n8758 & ~n8797;
  assign n8238 = ~n8042;
  assign n6381 = ~INSTQUEUE_REG_12__1__SCAN_IN | ~n8238;
  assign n6383 = ~n6382 | ~n6381;
  assign n6389 = ~n6942 & ~n7958;
  assign n6387 = ~INSTQUEUE_REG_11__1__SCAN_IN | ~n6749;
  assign n6385 = ~n9580 & ~n8797;
  assign n6673 = ~n6385;
  assign n8239 = ~n6673;
  assign n6386 = ~INSTQUEUE_REG_15__1__SCAN_IN | ~n8239;
  assign n6388 = ~n6387 | ~n6386;
  assign n6391 = ~n6389 & ~n6388;
  assign n6390 = ~n7484 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n6416 = ~n6391 | ~n6390;
  assign n6392 = ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n6668 = ~n6404 & ~n6408;
  assign n6395 = ~n6393;
  assign n6394 = ~n6403;
  assign n6396 = ~INSTQUEUE_REG_9__1__SCAN_IN | ~n7951;
  assign n6402 = ~n6397 | ~n6396;
  assign n6400 = ~n6301 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n6399 = ~n8222 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n6401 = ~n6400 | ~n6399;
  assign n6414 = ~n6402 & ~n6401;
  assign n6406 = ~INSTQUEUE_REG_5__1__SCAN_IN | ~n7996;
  assign n6674 = ~n9580 & ~n6407;
  assign n6456 = ~n6674;
  assign n6405 = ~INSTQUEUE_REG_3__1__SCAN_IN | ~n6725;
  assign n6412 = ~n6406 | ~n6405;
  assign n6679 = ~n6408 & ~n6407;
  assign n6425 = ~n6679;
  assign n7024 = ~n6425;
  assign n6410 = ~INSTQUEUE_REG_2__1__SCAN_IN | ~n7024;
  assign n6409 = ~INSTQUEUE_REG_14__1__SCAN_IN | ~n6683;
  assign n6411 = ~n6410 | ~n6409;
  assign n6413 = ~n6412 & ~n6411;
  assign n6415 = ~n6414 | ~n6413;
  assign n6420 = ~INSTQUEUE_REG_0__3__SCAN_IN | ~n6661;
  assign n6419 = ~INSTQUEUE_REG_14__3__SCAN_IN | ~n6683;
  assign n6424 = ~n6420 | ~n6419;
  assign n6422 = ~n6299 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n8119 = ~n7235;
  assign n6421 = ~n6285 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n6423 = ~n6422 | ~n6421;
  assign n6433 = ~n6424 & ~n6423;
  assign n8122 = ~n6425;
  assign n6427 = ~n8122 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n6426 = ~n8222 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n6431 = ~n6427 | ~n6426;
  assign n6429 = ~n8233 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n6428 = ~n6385 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n6430 = ~n6429 | ~n6428;
  assign n6432 = ~n6431 & ~n6430;
  assign n6435 = ~INSTQUEUE_REG_12__3__SCAN_IN | ~n6682;
  assign n6434 = ~INSTQUEUE_REG_11__3__SCAN_IN | ~n6749;
  assign n6439 = ~n6435 | ~n6434;
  assign n6436 = ~INSTQUEUE_REG_4__3__SCAN_IN | ~n6648;
  assign n6438 = ~n6437 | ~n6436;
  assign n6447 = ~n6439 & ~n6438;
  assign n6441 = ~INSTQUEUE_REG_6__3__SCAN_IN | ~n8182;
  assign n6440 = ~INSTQUEUE_REG_9__3__SCAN_IN | ~n7951;
  assign n6445 = ~n6441 | ~n6440;
  assign n6443 = ~INSTQUEUE_REG_5__3__SCAN_IN | ~n8230;
  assign n6442 = ~INSTQUEUE_REG_3__3__SCAN_IN | ~n6725;
  assign n6444 = ~n6443 | ~n6442;
  assign n6446 = ~n6445 & ~n6444;
  assign n6448 = ~n6447 | ~n6446;
  assign n9995 = ~n6843;
  assign n6451 = ~n8078 | ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n6450 = ~n7484 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n6455 = ~n6451 | ~n6450;
  assign n6453 = ~INSTQUEUE_REG_11__0__SCAN_IN | ~n6749;
  assign n6452 = ~INSTQUEUE_REG_2__0__SCAN_IN | ~n7024;
  assign n6454 = ~n6453 | ~n6452;
  assign n6464 = ~n6455 & ~n6454;
  assign n6458 = ~INSTQUEUE_REG_5__0__SCAN_IN | ~n7996;
  assign n6457 = ~INSTQUEUE_REG_3__0__SCAN_IN | ~n8188;
  assign n6462 = ~n6458 | ~n6457;
  assign n6460 = ~n6683 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n6459 = ~n6669 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n6461 = ~n6460 | ~n6459;
  assign n6463 = ~n6462 & ~n6461;
  assign n6480 = ~n6464 | ~n6463;
  assign n8162 = ~n6673;
  assign n6466 = ~INSTQUEUE_REG_15__0__SCAN_IN | ~n8162;
  assign n6465 = ~INSTQUEUE_REG_7__0__SCAN_IN | ~n6302;
  assign n6470 = ~n6466 | ~n6465;
  assign n6468 = ~INSTQUEUE_REG_4__0__SCAN_IN | ~n6648;
  assign n6467 = ~INSTQUEUE_REG_6__0__SCAN_IN | ~n8182;
  assign n6469 = ~n6468 | ~n6467;
  assign n6478 = ~n6470 & ~n6469;
  assign n6471 = ~INSTQUEUE_REG_9__0__SCAN_IN | ~n7951;
  assign n6476 = ~n6472 | ~n6471;
  assign n6474 = ~n8222 | ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n6473 = ~n8238 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n6475 = ~n6474 | ~n6473;
  assign n6477 = ~n6476 & ~n6475;
  assign n6479 = ~n6478 | ~n6477;
  assign n8441 = ~n6480 & ~n6479;
  assign n6529 = ~n6843 | ~n9821;
  assign n6523 = ~n6842 | ~n6529;
  assign n10181 = ~n6481;
  assign n6483 = ~EBX_REG_30__SCAN_IN | ~n10181;
  assign n6482 = ~INSTADDRPOINTER_REG_30__SCAN_IN | ~n6547;
  assign n8424 = ~n6483 | ~n6482;
  assign n6485 = ~INSTADDRPOINTER_REG_26__SCAN_IN | ~n6547;
  assign n6484 = ~EBX_REG_26__SCAN_IN | ~n10181;
  assign n6486 = ~n6485 | ~n6484;
  assign n9001 = n8434 ^ n6486;
  assign n6488 = ~EBX_REG_24__SCAN_IN | ~n10181;
  assign n6487 = ~INSTADDRPOINTER_REG_24__SCAN_IN | ~n6547;
  assign n6489 = ~n6488 | ~n6487;
  assign n12085 = n8434 ^ n6489;
  assign n6491 = ~EBX_REG_22__SCAN_IN | ~n10181;
  assign n6490 = ~INSTADDRPOINTER_REG_22__SCAN_IN | ~n6547;
  assign n6492 = ~n6491 | ~n6490;
  assign n8967 = n8434 ^ n6492;
  assign n6494 = ~EBX_REG_20__SCAN_IN | ~n10181;
  assign n6547 = ~n8410;
  assign n6493 = ~INSTADDRPOINTER_REG_20__SCAN_IN | ~n6547;
  assign n6495 = ~n6494 | ~n6493;
  assign n8864 = n8434 ^ n6495;
  assign n6497 = ~EBX_REG_18__SCAN_IN | ~n10181;
  assign n6496 = ~INSTADDRPOINTER_REG_18__SCAN_IN | ~n6547;
  assign n6498 = ~n6497 | ~n6496;
  assign n11955 = n8434 ^ n6498;
  assign n6500 = ~EBX_REG_16__SCAN_IN | ~n10181;
  assign n6499 = ~INSTADDRPOINTER_REG_16__SCAN_IN | ~n6547;
  assign n6501 = ~n6500 | ~n6499;
  assign n8985 = n8434 ^ n6501;
  assign n6503 = ~EBX_REG_14__SCAN_IN | ~n10181;
  assign n6502 = ~INSTADDRPOINTER_REG_14__SCAN_IN | ~n6547;
  assign n6504 = ~n6503 | ~n6502;
  assign n10822 = n8434 ^ n6504;
  assign n6506 = ~EBX_REG_12__SCAN_IN | ~n10181;
  assign n6505 = ~INSTADDRPOINTER_REG_12__SCAN_IN | ~n6547;
  assign n6507 = ~n6506 | ~n6505;
  assign n10500 = n8434 ^ n6507;
  assign n6509 = ~EBX_REG_10__SCAN_IN | ~n10181;
  assign n6508 = ~INSTADDRPOINTER_REG_10__SCAN_IN | ~n6547;
  assign n6510 = ~n6509 | ~n6508;
  assign n10238 = n8434 ^ n6510;
  assign n6512 = ~EBX_REG_8__SCAN_IN | ~n10181;
  assign n6511 = ~INSTADDRPOINTER_REG_8__SCAN_IN | ~n6547;
  assign n6513 = ~n6512 | ~n6511;
  assign n11109 = n8434 ^ n6513;
  assign n6515 = ~EBX_REG_6__SCAN_IN | ~n10181;
  assign n6514 = ~INSTADDRPOINTER_REG_6__SCAN_IN | ~n6547;
  assign n6516 = ~n6515 | ~n6514;
  assign n11415 = n8434 ^ n6516;
  assign n6518 = ~EBX_REG_4__SCAN_IN | ~n10181;
  assign n6517 = ~INSTADDRPOINTER_REG_4__SCAN_IN | ~n6547;
  assign n6519 = ~n6518 | ~n6517;
  assign n10114 = n8434 ^ n6519;
  assign n6521 = ~EBX_REG_2__SCAN_IN | ~n10181;
  assign n6520 = ~INSTADDRPOINTER_REG_2__SCAN_IN | ~n6547;
  assign n6522 = ~n6521 | ~n6520;
  assign n9716 = n8434 ^ n6522;
  assign n6526 = ~EBX_REG_1__SCAN_IN | ~n6523;
  assign n6524 = ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n6527 = ~n6526 | ~n6525;
  assign n6532 = n6528 ^ ~n6527;
  assign n6534 = ~n6532;
  assign n10184 = ~EBX_REG_0__SCAN_IN;
  assign n6531 = ~n6529 & ~n10184;
  assign n6530 = ~EBX_REG_0__SCAN_IN & ~n6842;
  assign n10183 = ~n6531 & ~n6530;
  assign n10949 = n6532 ^ n10183;
  assign n6533 = ~n8410 | ~n10949;
  assign n9715 = ~n6534 | ~n6533;
  assign n6536 = ~EBX_REG_3__SCAN_IN | ~n10181;
  assign n6535 = ~INSTADDRPOINTER_REG_3__SCAN_IN | ~n6547;
  assign n6537 = ~n6536 | ~n6535;
  assign n10579 = n8434 ^ ~n6537;
  assign n10113 = ~n10580 | ~n10579;
  assign n6539 = ~EBX_REG_5__SCAN_IN | ~n10181;
  assign n6538 = ~INSTADDRPOINTER_REG_5__SCAN_IN | ~n6547;
  assign n6540 = ~n6539 | ~n6538;
  assign n10655 = n8434 ^ ~n6540;
  assign n11414 = ~n10656 | ~n10655;
  assign n6542 = ~EBX_REG_7__SCAN_IN | ~n10181;
  assign n6541 = ~INSTADDRPOINTER_REG_7__SCAN_IN | ~n6547;
  assign n6543 = ~n6542 | ~n6541;
  assign n10787 = n8434 ^ ~n6543;
  assign n11108 = ~n10788 | ~n10787;
  assign n6545 = ~EBX_REG_9__SCAN_IN | ~n10181;
  assign n6544 = ~INSTADDRPOINTER_REG_9__SCAN_IN | ~n6547;
  assign n6546 = ~n6545 | ~n6544;
  assign n10121 = n8434 ^ ~n6546;
  assign n10237 = ~n10122 | ~n10121;
  assign n10343 = ~n10238 & ~n10237;
  assign n6549 = ~EBX_REG_11__SCAN_IN | ~n10181;
  assign n6548 = ~INSTADDRPOINTER_REG_11__SCAN_IN | ~n6547;
  assign n6550 = ~n6549 | ~n6548;
  assign n10342 = n8434 ^ ~n6550;
  assign n10499 = ~n10343 | ~n10342;
  assign n10828 = ~n10500 & ~n10499;
  assign n6552 = ~EBX_REG_13__SCAN_IN | ~n10181;
  assign n6551 = ~INSTADDRPOINTER_REG_13__SCAN_IN | ~n6547;
  assign n6553 = ~n6552 | ~n6551;
  assign n10827 = n8434 ^ ~n6553;
  assign n8899 = ~n10822 & ~n10821;
  assign n6555 = ~EBX_REG_15__SCAN_IN | ~n10181;
  assign n6554 = ~INSTADDRPOINTER_REG_15__SCAN_IN | ~n6547;
  assign n6556 = ~n6555 | ~n6554;
  assign n8898 = n8434 ^ ~n6556;
  assign n8984 = ~n8899 | ~n8898;
  assign n11935 = ~n8985 & ~n8984;
  assign n6558 = ~EBX_REG_17__SCAN_IN | ~n10181;
  assign n6557 = ~INSTADDRPOINTER_REG_17__SCAN_IN | ~n6547;
  assign n6559 = ~n6558 | ~n6557;
  assign n11934 = n8434 ^ ~n6559;
  assign n11918 = ~n11955 & ~n11954;
  assign n6561 = ~EBX_REG_19__SCAN_IN | ~n10181;
  assign n6560 = ~INSTADDRPOINTER_REG_19__SCAN_IN | ~n6547;
  assign n6562 = ~n6561 | ~n6560;
  assign n11917 = n8434 ^ ~n6562;
  assign n8863 = ~n11918 | ~n11917;
  assign n6564 = ~EBX_REG_21__SCAN_IN | ~n10181;
  assign n6563 = ~INSTADDRPOINTER_REG_21__SCAN_IN | ~n6547;
  assign n6565 = ~n6564 | ~n6563;
  assign n8839 = n8434 ^ ~n6565;
  assign n8966 = ~n8840 | ~n8839;
  assign n6567 = ~EBX_REG_23__SCAN_IN | ~n10181;
  assign n6566 = ~INSTADDRPOINTER_REG_23__SCAN_IN | ~n6547;
  assign n6568 = ~n6567 | ~n6566;
  assign n8932 = n8434 ^ ~n6568;
  assign n12084 = ~n8933 | ~n8932;
  assign n8511 = ~n12085 & ~n12084;
  assign n6570 = ~EBX_REG_25__SCAN_IN | ~n10181;
  assign n6569 = ~INSTADDRPOINTER_REG_25__SCAN_IN | ~n6547;
  assign n6571 = ~n6570 | ~n6569;
  assign n8510 = n8434 ^ ~n6571;
  assign n9000 = ~n8511 | ~n8510;
  assign n12172 = ~n9001 & ~n9000;
  assign n6573 = ~EBX_REG_27__SCAN_IN | ~n10181;
  assign n6572 = ~INSTADDRPOINTER_REG_27__SCAN_IN | ~n6547;
  assign n6574 = ~n6573 | ~n6572;
  assign n12171 = n8434 ^ ~n6574;
  assign n8603 = ~n12172 | ~n12171;
  assign n6576 = ~INSTADDRPOINTER_REG_28__SCAN_IN | ~n6547;
  assign n6575 = ~EBX_REG_28__SCAN_IN | ~n10181;
  assign n6577 = ~n6576 | ~n6575;
  assign n8604 = n8434 ^ n6577;
  assign n6579 = ~EBX_REG_29__SCAN_IN | ~n10181;
  assign n6578 = ~INSTADDRPOINTER_REG_29__SCAN_IN | ~n6547;
  assign n6580 = ~n6579 | ~n6578;
  assign n12289 = n8434 ^ ~n6580;
  assign n8423 = ~n12290 | ~n12289;
  assign n8425 = ~n8434 | ~n8423;
  assign n7951 = ~n6651;
  assign n6584 = ~INSTQUEUE_REG_9__7__SCAN_IN | ~n7951;
  assign n6589 = ~n6585 | ~n6584;
  assign n6587 = ~INSTQUEUE_REG_0__7__SCAN_IN | ~n6661;
  assign n6586 = ~INSTQUEUE_REG_5__7__SCAN_IN | ~n8230;
  assign n6588 = ~n6587 | ~n6586;
  assign n6597 = ~n6589 & ~n6588;
  assign n6591 = ~INSTQUEUE_REG_10__7__SCAN_IN | ~n6669;
  assign n6590 = ~INSTQUEUE_REG_4__7__SCAN_IN | ~n6648;
  assign n6595 = ~n6591 | ~n6590;
  assign n6593 = ~INSTQUEUE_REG_11__7__SCAN_IN | ~n6749;
  assign n6592 = ~INSTQUEUE_REG_2__7__SCAN_IN | ~n7024;
  assign n6594 = ~n6593 | ~n6592;
  assign n6596 = ~n6595 & ~n6594;
  assign n6599 = ~n6298 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n6598 = ~n8222 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n6604 = ~n6599 | ~n6598;
  assign n6600 = ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n6601 = ~INSTQUEUE_REG_7__7__SCAN_IN | ~n6302;
  assign n6603 = ~n6602 | ~n6601;
  assign n6605 = ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n6606 = ~n6725 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n6611 = ~n6607 | ~n6606;
  assign n6609 = ~INSTQUEUE_REG_15__7__SCAN_IN | ~n8239;
  assign n6608 = ~INSTQUEUE_REG_14__7__SCAN_IN | ~n6683;
  assign n6610 = ~n6609 | ~n6608;
  assign n9581 = ~STATE2_REG_0__SCAN_IN | ~n8795;
  assign n7686 = ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n6619 = ~n6942 & ~n7686;
  assign n6617 = ~INSTQUEUE_REG_14__2__SCAN_IN | ~n6683;
  assign n6616 = ~INSTQUEUE_REG_7__2__SCAN_IN | ~n6299;
  assign n6618 = ~n6617 | ~n6616;
  assign n6621 = ~n6619 & ~n6618;
  assign n6620 = ~n6285 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n6639 = ~n6621 | ~n6620;
  assign n6622 = ~INSTQUEUE_REG_2__2__SCAN_IN | ~n7024;
  assign n6627 = ~n6623 | ~n6622;
  assign n6625 = ~n8162 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n6624 = ~n6725 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n6626 = ~n6625 | ~n6624;
  assign n6637 = ~n6627 & ~n6626;
  assign n6630 = ~INSTQUEUE_REG_12__2__SCAN_IN | ~n6682;
  assign n6628 = ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n6629 = n6628 | n6692;
  assign n6635 = ~n6630 | ~n6629;
  assign n6633 = ~n8222 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n6631 = ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n6632 = n7377 | n6631;
  assign n6634 = ~n6633 | ~n6632;
  assign n6636 = ~n6635 & ~n6634;
  assign n6638 = ~n6637 | ~n6636;
  assign n6647 = ~n6639 & ~n6638;
  assign n6641 = ~INSTQUEUE_REG_4__2__SCAN_IN | ~n6648;
  assign n6640 = ~INSTQUEUE_REG_6__2__SCAN_IN | ~n8182;
  assign n6645 = ~n6641 | ~n6640;
  assign n6643 = ~INSTQUEUE_REG_11__2__SCAN_IN | ~n6749;
  assign n6642 = ~INSTQUEUE_REG_9__2__SCAN_IN | ~n7951;
  assign n6644 = ~n6643 | ~n6642;
  assign n6646 = ~n6645 & ~n6644;
  assign n10380 = ~n6647 | ~n6646;
  assign n6844 = ~n8690 | ~n8410;
  assign n6650 = ~INSTQUEUE_REG_1__4__SCAN_IN | ~n6293;
  assign n6649 = ~INSTQUEUE_REG_4__4__SCAN_IN | ~n6648;
  assign n6656 = ~n6650 | ~n6649;
  assign n6652 = ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n6653 = ~INSTQUEUE_REG_7__4__SCAN_IN | ~n6300;
  assign n6655 = ~n6654 | ~n6653;
  assign n6660 = ~n6284 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n6657 = ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n6665 = ~n6660 | ~n6659;
  assign n6663 = ~INSTQUEUE_REG_0__4__SCAN_IN | ~n6661;
  assign n6662 = ~INSTQUEUE_REG_11__4__SCAN_IN | ~n6749;
  assign n6664 = ~n6663 | ~n6662;
  assign n6666 = ~n6665 & ~n6664;
  assign n6691 = ~n6667 | ~n6666;
  assign n6671 = ~n6668 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n6670 = ~n6669 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n6678 = ~n6671 | ~n6670;
  assign n6672 = ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n6676 = n6673 | n6672;
  assign n6675 = ~n6674 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n6677 = ~n6676 | ~n6675;
  assign n6681 = ~n6297 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n6680 = ~n6679 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n6687 = ~n6681 | ~n6680;
  assign n6685 = ~INSTQUEUE_REG_12__4__SCAN_IN | ~n6682;
  assign n6684 = ~INSTQUEUE_REG_14__4__SCAN_IN | ~n6683;
  assign n6686 = ~n6685 | ~n6684;
  assign n6690 = ~n6689 | ~n6688;
  assign n6694 = ~INSTQUEUE_REG_5__5__SCAN_IN | ~n8181;
  assign n6693 = ~INSTQUEUE_REG_4__5__SCAN_IN | ~n6648;
  assign n6698 = ~n6694 | ~n6693;
  assign n6696 = ~INSTQUEUE_REG_6__5__SCAN_IN | ~n8182;
  assign n6695 = ~INSTQUEUE_REG_9__5__SCAN_IN | ~n7951;
  assign n6697 = ~n6696 | ~n6695;
  assign n6707 = ~n6698 & ~n6697;
  assign n6700 = ~INSTQUEUE_REG_12__5__SCAN_IN | ~n6682;
  assign n6699 = ~INSTQUEUE_REG_7__5__SCAN_IN | ~n6301;
  assign n6705 = ~n6700 | ~n6699;
  assign n6703 = ~n6749 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n6701 = ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n6702 = n7377 | n6701;
  assign n6704 = ~n6703 | ~n6702;
  assign n6706 = ~n6705 & ~n6704;
  assign n6724 = ~n6707 | ~n6706;
  assign n6708 = ~INSTQUEUE_REG_14__5__SCAN_IN | ~n6683;
  assign n6714 = ~n6709 | ~n6708;
  assign n6710 = ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n6712 = n6942 | n6710;
  assign n6711 = ~n8222 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n6713 = ~n6712 | ~n6711;
  assign n6722 = ~n6714 & ~n6713;
  assign n6716 = ~INSTQUEUE_REG_10__5__SCAN_IN | ~n6669;
  assign n6715 = ~INSTQUEUE_REG_15__5__SCAN_IN | ~n6385;
  assign n6720 = ~n6716 | ~n6715;
  assign n6718 = ~n7024 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n6717 = ~n6725 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n6719 = ~n6718 | ~n6717;
  assign n6721 = ~n6720 & ~n6719;
  assign n6723 = ~n6722 | ~n6721;
  assign n6727 = ~n6288 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n6726 = ~n6725 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n6732 = ~n6727 | ~n6726;
  assign n6728 = ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n6729 = ~INSTQUEUE_REG_9__6__SCAN_IN | ~n7951;
  assign n6731 = ~n6730 | ~n6729;
  assign n6740 = ~n6732 & ~n6731;
  assign n6734 = ~INSTQUEUE_REG_10__6__SCAN_IN | ~n6669;
  assign n6733 = ~INSTQUEUE_REG_4__6__SCAN_IN | ~n6648;
  assign n6738 = ~n6734 | ~n6733;
  assign n6736 = ~n7024 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n6735 = ~n6682 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n6737 = ~n6736 | ~n6735;
  assign n6739 = ~n6738 & ~n6737;
  assign n6742 = ~n6683 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n6741 = ~n8222 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n6746 = ~n6742 | ~n6741;
  assign n6744 = ~INSTQUEUE_REG_15__6__SCAN_IN | ~n8239;
  assign n6743 = ~INSTQUEUE_REG_7__6__SCAN_IN | ~n6299;
  assign n6745 = ~n6744 | ~n6743;
  assign n6756 = ~n6746 & ~n6745;
  assign n6748 = ~n8181 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n6747 = ~n6661 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n6754 = ~n6748 | ~n6747;
  assign n6752 = ~INSTQUEUE_REG_11__6__SCAN_IN | ~n6749;
  assign n6750 = ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n6753 = ~n6752 | ~n6751;
  assign n6755 = ~n6754 & ~n6753;
  assign n6757 = ~n6756 | ~n6755;
  assign n6808 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~n10866;
  assign n9589 = ~n9580;
  assign n6766 = ~n9589 | ~n11513;
  assign n6764 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~n11513;
  assign n6765 = ~n6782 | ~n9788;
  assign n6767 = ~n6766 | ~n6765;
  assign n6769 = ~n9591 | ~n6767;
  assign n6777 = n9591 ^ n6767;
  assign n6773 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n6774 = ~n6773 & ~INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n6820 = ~n7252 | ~n8392;
  assign n8290 = ~n9757 | ~n9736;
  assign n6811 = INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ ~n6776;
  assign n6780 = ~n6821 | ~n6811;
  assign n8388 = INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ ~n6777;
  assign n6797 = n7252 & n8388;
  assign n6778 = ~n9476 | ~n9736;
  assign n6795 = ~n8671 | ~n6778;
  assign n6779 = ~n6797 | ~n6795;
  assign n6807 = ~n6780 | ~n6779;
  assign n6781 = ~n7266 & ~n9476;
  assign n6784 = ~n8715 & ~n6781;
  assign n8390 = INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ n6782;
  assign n6783 = ~n7265 | ~n8390;
  assign n6802 = ~n6784 | ~n6783;
  assign n6786 = ~n6821;
  assign n6785 = n9734 | n8390;
  assign n6803 = ~n6786 | ~n6785;
  assign n6794 = ~n6802 | ~n6803;
  assign n6789 = INSTQUEUERD_ADDR_REG_0__SCAN_IN ^ ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n6787 = ~n7252 | ~n6789;
  assign n6792 = ~n6787 | ~n6786;
  assign n6788 = ~n8441 & ~n7589;
  assign n6790 = ~n6795 & ~n6788;
  assign n6791 = ~n6790 | ~n6789;
  assign n6793 = ~n6792 | ~n6791;
  assign n6801 = ~n6794 | ~n6793;
  assign n6799 = ~n6795;
  assign n6796 = ~n8388 & ~n7208;
  assign n6798 = ~n6797 & ~n6796;
  assign n6800 = ~n6799 | ~n6798;
  assign n6805 = ~n6801 | ~n6800;
  assign n6804 = ~n6803 & ~n6802;
  assign n6806 = ~n6805 & ~n6804;
  assign n6813 = ~n6807 & ~n6806;
  assign n6809 = ~n6808;
  assign n6814 = ~n6810 & ~n6809;
  assign n8387 = ~n6811 & ~n6814;
  assign n6812 = ~n8387 & ~n7266;
  assign n6818 = ~n6813 & ~n6812;
  assign n6816 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n9734;
  assign n6815 = ~n6821 | ~n6814;
  assign n6817 = ~n6816 | ~n6815;
  assign n6819 = ~n6818 & ~n6817;
  assign n6823 = ~n6820 | ~n6819;
  assign n6822 = ~n6821 | ~n8392;
  assign n7588 = ~n8443 & ~n8715;
  assign n6827 = ~n8550;
  assign n6829 = ~PHYADDRPOINTER_REG_3__SCAN_IN | ~n8114;
  assign n7133 = ~PHYADDRPOINTER_REG_2__SCAN_IN | ~PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n11806 = PHYADDRPOINTER_REG_3__SCAN_IN ^ n7133;
  assign n6828 = ~n8628 | ~n11806;
  assign n6831 = ~n6829 | ~n6828;
  assign n7112 = ~STATE2_REG_2__SCAN_IN | ~n12494;
  assign n6830 = ~n8716 & ~n7112;
  assign n6833 = ~n6831 & ~n6830;
  assign n7751 = ~n10732 & ~n10266;
  assign n6832 = ~n7751 | ~EAX_REG_3__SCAN_IN;
  assign n7091 = ~n6833 | ~n6832;
  assign n6834 = ~n8690 & ~n7589;
  assign n6853 = ~n6834 | ~n12494;
  assign n6836 = ~n8443 | ~n6835;
  assign n7602 = ~n12492 & ~n10380;
  assign n6837 = ~n6836 | ~n7602;
  assign n6839 = ~n6853 | ~n6837;
  assign n6838 = ~n8376 | ~n9995;
  assign n7591 = ~n6843 | ~n8690;
  assign n6848 = ~n6857 | ~n10876;
  assign n6841 = ~n6843 & ~n6840;
  assign n6864 = ~n6841 | ~n9821;
  assign n6846 = ~n6864 & ~n8711;
  assign n8399 = ~n8429 | ~n8378;
  assign n6858 = ~n6845 | ~n6844;
  assign n6847 = ~n6846 | ~n6858;
  assign n6849 = ~n6848 | ~n6847;
  assign n6855 = ~n6849 | ~n8377;
  assign n8577 = ~n12492 & ~n9736;
  assign n8398 = ~n6850 | ~n8577;
  assign n8386 = STATE_REG_2__SCAN_IN ^ ~STATE_REG_1__SCAN_IN;
  assign n6852 = ~n8386 | ~n9476;
  assign n6854 = ~n8669 | ~n6852;
  assign n6880 = ~n6854 | ~n8712;
  assign n6856 = ~n6855 & ~n6880;
  assign n6892 = ~n6856 & ~n9734;
  assign n6860 = ~n6857 | ~n8441;
  assign n6859 = ~n6858;
  assign n6862 = ~n6860 | ~n6859;
  assign n9472 = ~n8441 & ~n9757;
  assign n6861 = ~n8377 | ~n8575;
  assign n7596 = ~n9472 | ~n6861;
  assign n11900 = ~STATE2_REG_0__SCAN_IN | ~n9623;
  assign n6863 = ~n8377;
  assign n6865 = ~n6864 & ~n6863;
  assign n6866 = ~n9476 & ~n6865;
  assign n6867 = ~n11900 & ~n6866;
  assign n6869 = ~n7117 & ~n6763;
  assign n6873 = ~n6892 | ~n6869;
  assign n6893 = ~n8795;
  assign n6871 = ~n6893 & ~n11513;
  assign n8457 = ~n9623 | ~n9734;
  assign n8487 = ~n8457;
  assign n6870 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n8487;
  assign n7115 = ~n6871 & ~n6870;
  assign n6937 = ~n6873 | ~n6872;
  assign n6876 = ~n8795 & ~n9788;
  assign n8763 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n6874 = ~n11513 | ~n9788;
  assign n11283 = ~n8763 | ~n6874;
  assign n6875 = ~n11283 & ~n8457;
  assign n6936 = ~n6878 | ~n6877;
  assign n6882 = ~n6936;
  assign n8565 = ~n8671 & ~n7591;
  assign n6879 = ~n8715 | ~n8565;
  assign n6883 = ~n6882 | ~n6935;
  assign n6885 = ~n6937 | ~n6883;
  assign n6884 = ~n6934 | ~n6936;
  assign n7113 = ~n6892;
  assign n6888 = ~n6376 & ~n7113;
  assign n10039 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n10029 = ~n11513 & ~n10039;
  assign n6896 = ~n10029;
  assign n6886 = ~n9787 | ~n8763;
  assign n10153 = ~n6896 | ~n6886;
  assign n6887 = ~n8457 & ~n10153;
  assign n6890 = ~n6888 & ~n6887;
  assign n6889 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~n6893;
  assign n6891 = ~n7051;
  assign n6895 = ~n6892 | ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n6894 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n6893;
  assign n6898 = ~n6895 | ~n6894;
  assign n10731 = INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ n6896;
  assign n6897 = ~n8457 & ~n10731;
  assign n6900 = ~INSTQUEUE_REG_12__3__SCAN_IN | ~n6303;
  assign n6899 = ~INSTQUEUE_REG_0__3__SCAN_IN | ~n8162;
  assign n6904 = ~n6900 | ~n6899;
  assign n6902 = ~INSTQUEUE_REG_6__3__SCAN_IN | ~n6292;
  assign n6901 = ~INSTQUEUE_REG_4__3__SCAN_IN | ~n8188;
  assign n6903 = ~n6902 | ~n6901;
  assign n6912 = ~n6904 & ~n6903;
  assign n6906 = ~n8137 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n6905 = ~n6293 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n6910 = ~n6906 | ~n6905;
  assign n6908 = ~INSTQUEUE_REG_5__3__SCAN_IN | ~n8187;
  assign n6907 = ~INSTQUEUE_REG_1__3__SCAN_IN | ~n8178;
  assign n6909 = ~n6908 | ~n6907;
  assign n6911 = ~n6910 & ~n6909;
  assign n6929 = ~n6912 | ~n6911;
  assign n6914 = ~n8238 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n6913 = ~n8119 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n6918 = ~n6914 | ~n6913;
  assign n6916 = ~INSTQUEUE_REG_3__3__SCAN_IN | ~n8242;
  assign n6915 = ~INSTQUEUE_REG_15__3__SCAN_IN | ~n8169;
  assign n6917 = ~n6916 | ~n6915;
  assign n6927 = ~n6918 & ~n6917;
  assign n6920 = ~n7484 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n6919 = ~n8138 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n6925 = ~n6920 | ~n6919;
  assign n6923 = ~INSTQUEUE_REG_10__3__SCAN_IN | ~n8219;
  assign n6922 = ~INSTQUEUE_REG_8__3__SCAN_IN | ~n6302;
  assign n6924 = ~n6923 | ~n6922;
  assign n6926 = ~n6925 & ~n6924;
  assign n6928 = ~n6927 | ~n6926;
  assign n8306 = ~n6929 & ~n6928;
  assign n6931 = n8306 | n7266;
  assign n6930 = ~INSTQUEUE_REG_0__3__SCAN_IN | ~n7265;
  assign n10956 = n6938 ^ ~n6937;
  assign n7006 = ~n6939 | ~n9734;
  assign n6940 = ~INSTQUEUE_REG_5__7__SCAN_IN | ~n8187;
  assign n6946 = ~n6941 | ~n6940;
  assign n6944 = ~n8118 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n6943 = ~n8178 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n6945 = ~n6944 | ~n6943;
  assign n6954 = ~n6946 & ~n6945;
  assign n6948 = ~INSTQUEUE_REG_0__7__SCAN_IN | ~n8239;
  assign n6947 = ~INSTQUEUE_REG_7__7__SCAN_IN | ~n8182;
  assign n6952 = ~n6948 | ~n6947;
  assign n6950 = ~INSTQUEUE_REG_6__7__SCAN_IN | ~n6291;
  assign n6949 = ~INSTQUEUE_REG_15__7__SCAN_IN | ~n8169;
  assign n6951 = ~n6950 | ~n6949;
  assign n6953 = ~n6952 & ~n6951;
  assign n6971 = ~n6954 | ~n6953;
  assign n6956 = ~INSTQUEUE_REG_3__7__SCAN_IN | ~n7024;
  assign n6955 = ~INSTQUEUE_REG_8__7__SCAN_IN | ~n6300;
  assign n6960 = ~n6956 | ~n6955;
  assign n6958 = ~n7484 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n6957 = ~n8138 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n6959 = ~n6958 | ~n6957;
  assign n6969 = ~n6960 & ~n6959;
  assign n6963 = ~INSTQUEUE_REG_12__7__SCAN_IN | ~n6287;
  assign n6962 = ~INSTQUEUE_REG_4__7__SCAN_IN | ~n8188;
  assign n6967 = ~n6963 | ~n6962;
  assign n6965 = ~INSTQUEUE_REG_11__7__SCAN_IN | ~n8229;
  assign n6964 = ~INSTQUEUE_REG_10__7__SCAN_IN | ~n7951;
  assign n6966 = ~n6965 | ~n6964;
  assign n6968 = ~n6967 & ~n6966;
  assign n6970 = ~n6969 | ~n6968;
  assign n6973 = ~n7046 | ~n8345;
  assign n6972 = ~n7265 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n7007 = ~n6973 | ~n6972;
  assign n8187 = ~n6974;
  assign n6976 = ~n8187 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n6975 = ~n7484 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n6980 = ~n6976 | ~n6975;
  assign n6978 = ~n6292 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n6977 = ~n8118 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n6979 = ~n6978 | ~n6977;
  assign n7004 = ~n6980 & ~n6979;
  assign n6982 = ~n6288 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n6981 = ~INSTQUEUE_REG_8__1__SCAN_IN | ~n6300;
  assign n6984 = ~n6982 | ~n6981;
  assign n6983 = n8178 & INSTQUEUE_REG_1__1__SCAN_IN;
  assign n6986 = ~n6984 & ~n6983;
  assign n6985 = ~n8138 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n7002 = ~n6986 | ~n6985;
  assign n6988 = ~INSTQUEUE_REG_12__1__SCAN_IN | ~n6287;
  assign n6987 = ~INSTQUEUE_REG_0__1__SCAN_IN | ~n8162;
  assign n6992 = ~n6988 | ~n6987;
  assign n6990 = ~INSTQUEUE_REG_15__1__SCAN_IN | ~n8169;
  assign n6989 = ~n8137 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n6991 = ~n6990 | ~n6989;
  assign n7000 = ~n6992 & ~n6991;
  assign n6994 = ~n8122 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n6993 = ~INSTQUEUE_REG_10__1__SCAN_IN | ~n8219;
  assign n6998 = ~n6994 | ~n6993;
  assign n6996 = ~n8212 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n6995 = ~INSTQUEUE_REG_11__1__SCAN_IN | ~n8119;
  assign n6997 = ~n6996 | ~n6995;
  assign n6999 = ~n6998 & ~n6997;
  assign n7001 = ~n7000 | ~n6999;
  assign n7003 = ~n7002 & ~n7001;
  assign n8292 = ~n7004 | ~n7003;
  assign n8276 = ~n8292;
  assign n7008 = ~n7046 | ~n7007;
  assign n7042 = ~INSTQUEUE_REG_0__0__SCAN_IN | ~n7009;
  assign n7011 = ~n8119 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n7010 = ~n8138 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n7015 = ~n7011 | ~n7010;
  assign n7013 = ~INSTQUEUE_REG_13__0__SCAN_IN | ~n8238;
  assign n7012 = ~INSTQUEUE_REG_0__0__SCAN_IN | ~n8162;
  assign n7014 = ~n7013 | ~n7012;
  assign n7040 = ~n7015 & ~n7014;
  assign n7016 = ~INSTQUEUE_REG_8__0__SCAN_IN | ~n6301;
  assign n7019 = ~n7017 | ~n7016;
  assign n7018 = n8212 & INSTQUEUE_REG_4__0__SCAN_IN;
  assign n7021 = ~n7019 & ~n7018;
  assign n7020 = ~n7484 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n7038 = ~n7021 | ~n7020;
  assign n7023 = ~n8137 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n7022 = ~n8178 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n7028 = ~n7023 | ~n7022;
  assign n7026 = ~INSTQUEUE_REG_3__0__SCAN_IN | ~n7024;
  assign n7025 = ~INSTQUEUE_REG_10__0__SCAN_IN | ~n7951;
  assign n7027 = ~n7026 | ~n7025;
  assign n7036 = ~n7028 & ~n7027;
  assign n7030 = ~INSTQUEUE_REG_12__0__SCAN_IN | ~n6287;
  assign n7029 = ~INSTQUEUE_REG_15__0__SCAN_IN | ~n8169;
  assign n7034 = ~n7030 | ~n7029;
  assign n7032 = ~INSTQUEUE_REG_5__0__SCAN_IN | ~n8187;
  assign n7031 = ~INSTQUEUE_REG_6__0__SCAN_IN | ~n6292;
  assign n7033 = ~n7032 | ~n7031;
  assign n7035 = ~n7034 & ~n7033;
  assign n7037 = ~n7036 | ~n7035;
  assign n7039 = ~n7038 & ~n7037;
  assign n8291 = ~n7040 | ~n7039;
  assign n7041 = ~n8441 | ~n8291;
  assign n7044 = ~n7042 | ~n7041;
  assign n7048 = ~n10219 & ~n8345;
  assign n7043 = n9734 | n7048;
  assign n7045 = n8345 ^ n8282;
  assign n7123 = ~n7046 | ~n7045;
  assign n7047 = ~n7122 & ~n7123;
  assign n7125 = ~STATE2_REG_0__SCAN_IN & ~n7115;
  assign n7049 = ~n7047 & ~n7125;
  assign n8272 = ~STATE2_REG_0__SCAN_IN | ~n7048;
  assign n7103 = ~n7049 | ~n8272;
  assign n7052 = ~n7050;
  assign n9889 = ~n7052 | ~n7051;
  assign n7055 = ~n6295 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n7054 = ~n8138 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n7059 = ~n7055 | ~n7054;
  assign n7057 = ~INSTQUEUE_REG_5__2__SCAN_IN | ~n8187;
  assign n7056 = ~INSTQUEUE_REG_0__2__SCAN_IN | ~n8162;
  assign n7058 = ~n7057 | ~n7056;
  assign n7067 = ~n7059 & ~n7058;
  assign n7061 = ~n8118 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n7060 = ~n8188 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n7065 = ~n7061 | ~n7060;
  assign n7063 = ~n6292 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n7062 = ~n8178 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n7064 = ~n7063 | ~n7062;
  assign n7066 = ~n7065 & ~n7064;
  assign n7084 = ~n7067 | ~n7066;
  assign n7070 = ~INSTQUEUE_REG_3__2__SCAN_IN | ~n8242;
  assign n7069 = ~INSTQUEUE_REG_7__2__SCAN_IN | ~n8137;
  assign n7074 = ~n7070 | ~n7069;
  assign n7072 = ~INSTQUEUE_REG_15__2__SCAN_IN | ~n8169;
  assign n7071 = ~INSTQUEUE_REG_8__2__SCAN_IN | ~n6302;
  assign n7073 = ~n7072 | ~n7071;
  assign n7082 = ~n7074 & ~n7073;
  assign n7076 = ~n7484 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n7075 = ~n8119 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n7080 = ~n7076 | ~n7075;
  assign n7078 = ~INSTQUEUE_REG_12__2__SCAN_IN | ~n6303;
  assign n7077 = ~INSTQUEUE_REG_10__2__SCAN_IN | ~n8219;
  assign n7079 = ~n7078 | ~n7077;
  assign n7081 = ~n7080 & ~n7079;
  assign n7083 = ~n7082 | ~n7081;
  assign n8299 = ~n7084 & ~n7083;
  assign n7085 = ~n8299 & ~n7266;
  assign n7094 = ~n7093 | ~n7092;
  assign n7177 = ~n10035 & ~n7094;
  assign n9557 = ~n7091 & ~n7090;
  assign n7095 = ~n9767;
  assign n7100 = ~n7095 | ~n8260;
  assign n11508 = PHYADDRPOINTER_REG_2__SCAN_IN ^ ~PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n7096 = ~STATEBS16_REG_SCAN_IN & ~n11508;
  assign n7098 = STATE2_REG_2__SCAN_IN | n7096;
  assign n7097 = ~EAX_REG_2__SCAN_IN | ~n7751;
  assign n7173 = ~n7112;
  assign n7101 = ~n7100 | ~n7099;
  assign n7130 = ~PHYADDRPOINTER_REG_2__SCAN_IN | ~n8114;
  assign n9573 = ~n7101 | ~n7130;
  assign n9737 = n7105 ^ ~n7104;
  assign n7111 = ~n7106 | ~n8260;
  assign n7108 = ~PHYADDRPOINTER_REG_1__SCAN_IN | ~n10732;
  assign n7107 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~n7173;
  assign n7109 = ~n7108 | ~n7107;
  assign n7119 = ~n6763 & ~n7112;
  assign n7114 = ~n7113 & ~n6763;
  assign n7116 = ~n7115 & ~n7114;
  assign n11167 = n7117 ^ ~n7116;
  assign n7118 = ~n11167 & ~n7580;
  assign n7121 = ~n7119 & ~n7118;
  assign n7120 = ~n7751 | ~EAX_REG_0__SCAN_IN;
  assign n9446 = ~n7121 | ~n7120;
  assign n7129 = ~n8628 & ~n9446;
  assign n7124 = n7123 ^ ~n7122;
  assign n7126 = ~n9779 & ~n6759;
  assign n9444 = ~n7126 & ~n10732;
  assign n9455 = ~PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n7127 = ~n9455 & ~STATE2_REG_2__SCAN_IN;
  assign n7128 = ~n9446 & ~n7127;
  assign n9448 = ~n9444 & ~n7128;
  assign n9466 = ~n7129 & ~n9448;
  assign n7131 = ~n7130;
  assign n9558 = ~n7132 & ~n7131;
  assign n7135 = ~PHYADDRPOINTER_REG_4__SCAN_IN | ~n8114;
  assign n11793 = ~PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n10891 = PHYADDRPOINTER_REG_4__SCAN_IN ^ n7214;
  assign n7134 = ~n8628 | ~n10891;
  assign n7172 = ~n7135 | ~n7134;
  assign n7170 = ~EAX_REG_4__SCAN_IN | ~n7751;
  assign n7167 = ~INSTQUEUE_REG_0__4__SCAN_IN | ~n7265;
  assign n7137 = ~n8118 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n7136 = ~n7484 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n7141 = ~n7137 | ~n7136;
  assign n7139 = ~INSTQUEUE_REG_12__4__SCAN_IN | ~n6303;
  assign n7138 = ~INSTQUEUE_REG_0__4__SCAN_IN | ~n8162;
  assign n7140 = ~n7139 | ~n7138;
  assign n7165 = ~n7141 & ~n7140;
  assign n7143 = ~INSTQUEUE_REG_11__4__SCAN_IN | ~n8119;
  assign n7142 = ~INSTQUEUE_REG_8__4__SCAN_IN | ~n6299;
  assign n7145 = ~n7143 | ~n7142;
  assign n7144 = n8242 & INSTQUEUE_REG_3__4__SCAN_IN;
  assign n7147 = ~n7145 & ~n7144;
  assign n7146 = ~n8137 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n7163 = ~n7147 | ~n7146;
  assign n7149 = ~INSTQUEUE_REG_5__4__SCAN_IN | ~n8187;
  assign n7148 = ~INSTQUEUE_REG_15__4__SCAN_IN | ~n8169;
  assign n7153 = ~n7149 | ~n7148;
  assign n7150 = ~INSTQUEUE_REG_6__4__SCAN_IN | ~n6292;
  assign n7152 = ~n7151 | ~n7150;
  assign n7161 = ~n7153 & ~n7152;
  assign n7155 = ~n8188 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n7154 = ~n8138 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n7159 = ~n7155 | ~n7154;
  assign n7157 = ~INSTQUEUE_REG_1__4__SCAN_IN | ~n8178;
  assign n7156 = ~INSTQUEUE_REG_10__4__SCAN_IN | ~n8219;
  assign n7158 = ~n7157 | ~n7156;
  assign n7160 = ~n7159 & ~n7158;
  assign n7162 = ~n7161 | ~n7160;
  assign n7164 = ~n7163 & ~n7162;
  assign n8311 = ~n7165 | ~n7164;
  assign n7166 = ~n7252 | ~n8311;
  assign n7176 = ~n7167 | ~n7166;
  assign n7171 = ~n7170 | ~n7169;
  assign n7175 = ~n7172 & ~n7171;
  assign n7174 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n7173;
  assign n9563 = ~n7175 | ~n7174;
  assign n9601 = ~n9564 | ~n9563;
  assign n7213 = ~n8114 | ~PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n7179 = ~INSTQUEUE_REG_15__5__SCAN_IN | ~n6683;
  assign n7178 = ~INSTQUEUE_REG_8__5__SCAN_IN | ~n6299;
  assign n7183 = ~n7179 | ~n7178;
  assign n7181 = ~INSTQUEUE_REG_5__5__SCAN_IN | ~n8187;
  assign n7180 = ~INSTQUEUE_REG_13__5__SCAN_IN | ~n8118;
  assign n7182 = ~n7181 | ~n7180;
  assign n7191 = ~n7183 & ~n7182;
  assign n7185 = ~n8122 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n7184 = ~n8178 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n7189 = ~n7185 | ~n7184;
  assign n7187 = ~INSTQUEUE_REG_9__5__SCAN_IN | ~n7484;
  assign n7186 = ~INSTQUEUE_REG_10__5__SCAN_IN | ~n8219;
  assign n7188 = ~n7187 | ~n7186;
  assign n7190 = ~n7189 & ~n7188;
  assign n7207 = ~n7191 | ~n7190;
  assign n7193 = ~INSTQUEUE_REG_11__5__SCAN_IN | ~n8119;
  assign n7192 = ~INSTQUEUE_REG_12__5__SCAN_IN | ~n6303;
  assign n7197 = ~n7193 | ~n7192;
  assign n7195 = ~n8138 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n7194 = ~n6294 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n7196 = ~n7195 | ~n7194;
  assign n7205 = ~n7197 & ~n7196;
  assign n7199 = ~INSTQUEUE_REG_0__5__SCAN_IN | ~n8162;
  assign n7198 = ~INSTQUEUE_REG_7__5__SCAN_IN | ~n8182;
  assign n7203 = ~n7199 | ~n7198;
  assign n7201 = ~n6292 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n7200 = ~n8212 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n7202 = ~n7201 | ~n7200;
  assign n7204 = ~n7203 & ~n7202;
  assign n7206 = ~n7205 | ~n7204;
  assign n8324 = ~n7207 & ~n7206;
  assign n7210 = ~n8324 & ~n7266;
  assign n7209 = ~n7208 & ~n6710;
  assign n7212 = ~n8260 | ~n8314;
  assign n7218 = ~n7213 | ~n7212;
  assign n7216 = ~n7751 | ~EAX_REG_5__SCAN_IN;
  assign n11867 = PHYADDRPOINTER_REG_5__SCAN_IN ^ ~n7256;
  assign n7215 = ~n8628 | ~n11867;
  assign n7217 = ~n7216 | ~n7215;
  assign n7254 = ~n7265 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n7222 = ~INSTQUEUE_REG_12__6__SCAN_IN | ~n6303;
  assign n7221 = ~INSTQUEUE_REG_7__6__SCAN_IN | ~n8182;
  assign n7226 = ~n7222 | ~n7221;
  assign n7224 = ~INSTQUEUE_REG_10__6__SCAN_IN | ~n8219;
  assign n7223 = ~INSTQUEUE_REG_14__6__SCAN_IN | ~n8222;
  assign n7225 = ~n7224 | ~n7223;
  assign n7251 = ~n7226 & ~n7225;
  assign n7228 = ~INSTQUEUE_REG_5__6__SCAN_IN | ~n8187;
  assign n7227 = ~INSTQUEUE_REG_1__6__SCAN_IN | ~n8178;
  assign n7230 = ~n7228 | ~n7227;
  assign n7229 = n7484 & INSTQUEUE_REG_9__6__SCAN_IN;
  assign n7232 = ~n7230 & ~n7229;
  assign n7231 = ~n8212 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n7249 = ~n7232 | ~n7231;
  assign n7234 = ~INSTQUEUE_REG_13__6__SCAN_IN | ~n8238;
  assign n7233 = ~INSTQUEUE_REG_15__6__SCAN_IN | ~n8169;
  assign n7239 = ~n7234 | ~n7233;
  assign n8229 = ~n7235;
  assign n7237 = ~INSTQUEUE_REG_11__6__SCAN_IN | ~n8119;
  assign n7236 = ~INSTQUEUE_REG_0__6__SCAN_IN | ~n8162;
  assign n7238 = ~n7237 | ~n7236;
  assign n7247 = ~n7239 & ~n7238;
  assign n7241 = ~INSTQUEUE_REG_6__6__SCAN_IN | ~n6292;
  assign n7240 = ~INSTQUEUE_REG_8__6__SCAN_IN | ~n6300;
  assign n7245 = ~n7241 | ~n7240;
  assign n7242 = ~INSTQUEUE_REG_3__6__SCAN_IN | ~n8242;
  assign n7244 = ~n7243 | ~n7242;
  assign n7246 = ~n7245 & ~n7244;
  assign n7248 = ~n7247 | ~n7246;
  assign n7250 = ~n7249 & ~n7248;
  assign n8334 = ~n7251 | ~n7250;
  assign n7253 = ~n7252 | ~n8334;
  assign n7263 = ~n7254 | ~n7253;
  assign n7258 = ~n7751 | ~EAX_REG_6__SCAN_IN;
  assign n11677 = PHYADDRPOINTER_REG_6__SCAN_IN ^ n7272;
  assign n7257 = ~n8628 | ~n11677;
  assign n7259 = ~n7258 | ~n7257;
  assign n7261 = ~PHYADDRPOINTER_REG_6__SCAN_IN | ~n8114;
  assign n7271 = ~EAX_REG_7__SCAN_IN | ~n7751;
  assign n7268 = ~n7265 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n7267 = n7266 | n8345;
  assign n7269 = ~n7268 | ~n7267;
  assign n7270 = ~n8337 | ~n8260;
  assign n7276 = ~n7271 | ~n7270;
  assign n7274 = ~PHYADDRPOINTER_REG_7__SCAN_IN | ~n8114;
  assign n11641 = PHYADDRPOINTER_REG_7__SCAN_IN ^ ~n7308;
  assign n7273 = ~n8628 | ~n11641;
  assign n7275 = ~n7274 | ~n7273;
  assign n9917 = ~n7276 & ~n7275;
  assign n10081 = ~n9917;
  assign n7278 = ~INSTQUEUE_REG_5__0__SCAN_IN | ~n8212;
  assign n7277 = ~INSTQUEUE_REG_11__0__SCAN_IN | ~n8219;
  assign n7282 = ~n7278 | ~n7277;
  assign n7280 = ~n8119 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n7279 = ~n7484 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n7281 = ~n7280 | ~n7279;
  assign n7290 = ~n7282 & ~n7281;
  assign n7284 = ~INSTQUEUE_REG_13__0__SCAN_IN | ~n6303;
  assign n7283 = ~INSTQUEUE_REG_4__0__SCAN_IN | ~n8242;
  assign n7288 = ~n7284 | ~n7283;
  assign n7286 = ~n8138 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n7285 = ~n6288 | ~INSTQUEUE_REG_3__0__SCAN_IN;
  assign n7287 = ~n7286 | ~n7285;
  assign n7289 = ~n7288 & ~n7287;
  assign n7306 = ~n7290 | ~n7289;
  assign n7292 = ~INSTQUEUE_REG_6__0__SCAN_IN | ~n8187;
  assign n7291 = ~INSTQUEUE_REG_8__0__SCAN_IN | ~n8137;
  assign n7296 = ~n7292 | ~n7291;
  assign n7294 = ~INSTQUEUE_REG_14__0__SCAN_IN | ~n8238;
  assign n7293 = ~INSTQUEUE_REG_7__0__SCAN_IN | ~n6292;
  assign n7295 = ~n7294 | ~n7293;
  assign n7304 = ~n7296 & ~n7295;
  assign n7298 = ~INSTQUEUE_REG_2__0__SCAN_IN | ~n8178;
  assign n7297 = ~INSTQUEUE_REG_0__0__SCAN_IN | ~n8169;
  assign n7302 = ~n7298 | ~n7297;
  assign n7300 = ~INSTQUEUE_REG_1__0__SCAN_IN | ~n8162;
  assign n7299 = ~INSTQUEUE_REG_9__0__SCAN_IN | ~n6301;
  assign n7301 = ~n7300 | ~n7299;
  assign n7303 = ~n7302 & ~n7301;
  assign n7305 = ~n7304 | ~n7303;
  assign n7307 = ~n7306 & ~n7305;
  assign n7312 = ~n7580 & ~n7307;
  assign n7310 = ~n7751 | ~EAX_REG_8__SCAN_IN;
  assign n11850 = PHYADDRPOINTER_REG_8__SCAN_IN ^ n7317;
  assign n7309 = ~n8628 | ~n11850;
  assign n7311 = ~n7310 | ~n7309;
  assign n7314 = ~n7312 & ~n7311;
  assign n7313 = ~PHYADDRPOINTER_REG_8__SCAN_IN | ~n8114;
  assign n10082 = ~n7314 | ~n7313;
  assign n7319 = ~PHYADDRPOINTER_REG_9__SCAN_IN | ~n8114;
  assign n11604 = PHYADDRPOINTER_REG_9__SCAN_IN ^ ~n7391;
  assign n7318 = ~n8628 | ~n11604;
  assign n7354 = ~n7319 | ~n7318;
  assign n7321 = ~INSTQUEUE_REG_4__1__SCAN_IN | ~n8242;
  assign n7323 = ~n7321 | ~n7320;
  assign n7322 = ~n8719 & ~n7958;
  assign n7325 = ~n7323 & ~n7322;
  assign n7324 = ~n7484 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n7341 = ~n7325 | ~n7324;
  assign n7327 = ~n8187 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n7326 = ~INSTQUEUE_REG_15__1__SCAN_IN | ~n8222;
  assign n7331 = ~n7327 | ~n7326;
  assign n7329 = ~n8239 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n7328 = ~n8137 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n7330 = ~n7329 | ~n7328;
  assign n7339 = ~n7331 & ~n7330;
  assign n7333 = ~n8188 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n7332 = ~INSTQUEUE_REG_14__1__SCAN_IN | ~n8238;
  assign n7337 = ~n7333 | ~n7332;
  assign n7335 = ~INSTQUEUE_REG_2__1__SCAN_IN | ~n8178;
  assign n7334 = ~INSTQUEUE_REG_12__1__SCAN_IN | ~n8119;
  assign n7336 = ~n7335 | ~n7334;
  assign n7338 = ~n7337 & ~n7336;
  assign n7340 = ~n7339 | ~n7338;
  assign n7349 = ~n7341 & ~n7340;
  assign n7343 = ~INSTQUEUE_REG_11__1__SCAN_IN | ~n8219;
  assign n7342 = ~n6303 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n7347 = ~n7343 | ~n7342;
  assign n7345 = ~n6292 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n7344 = ~INSTQUEUE_REG_9__1__SCAN_IN | ~n6301;
  assign n7346 = ~n7345 | ~n7344;
  assign n7348 = ~n7347 & ~n7346;
  assign n7350 = ~n7349 | ~n7348;
  assign n7352 = ~n8260 | ~n7350;
  assign n7351 = ~n7751 | ~EAX_REG_9__SCAN_IN;
  assign n7353 = ~n7352 | ~n7351;
  assign n10240 = ~n10074 & ~n10073;
  assign n7356 = ~INSTQUEUE_REG_14__2__SCAN_IN | ~n8238;
  assign n7355 = ~INSTQUEUE_REG_7__2__SCAN_IN | ~n6292;
  assign n7360 = ~n7356 | ~n7355;
  assign n7358 = ~INSTQUEUE_REG_13__2__SCAN_IN | ~n6303;
  assign n7357 = ~INSTQUEUE_REG_4__2__SCAN_IN | ~n8242;
  assign n7359 = ~n7358 | ~n7357;
  assign n7368 = ~n7360 & ~n7359;
  assign n7362 = ~n8188 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n7361 = ~n8119 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n7366 = ~n7362 | ~n7361;
  assign n7364 = ~INSTQUEUE_REG_6__2__SCAN_IN | ~n8187;
  assign n7363 = ~INSTQUEUE_REG_1__2__SCAN_IN | ~n8162;
  assign n7365 = ~n7364 | ~n7363;
  assign n7367 = ~n7366 & ~n7365;
  assign n7385 = ~n7368 | ~n7367;
  assign n7370 = ~INSTQUEUE_REG_3__2__SCAN_IN | ~n6294;
  assign n7369 = ~INSTQUEUE_REG_0__2__SCAN_IN | ~n8169;
  assign n7374 = ~n7370 | ~n7369;
  assign n7372 = ~INSTQUEUE_REG_2__2__SCAN_IN | ~n8178;
  assign n7371 = ~INSTQUEUE_REG_11__2__SCAN_IN | ~n8219;
  assign n7373 = ~n7372 | ~n7371;
  assign n7383 = ~n7374 & ~n7373;
  assign n7376 = ~INSTQUEUE_REG_8__2__SCAN_IN | ~n8137;
  assign n7375 = ~INSTQUEUE_REG_9__2__SCAN_IN | ~n6300;
  assign n7381 = ~n7376 | ~n7375;
  assign n7379 = ~n8138 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n7378 = ~n8233 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n7380 = ~n7379 | ~n7378;
  assign n7382 = ~n7381 & ~n7380;
  assign n7384 = ~n7383 | ~n7382;
  assign n7386 = ~n7385 & ~n7384;
  assign n7390 = ~n7580 & ~n7386;
  assign n7388 = ~n7751 | ~EAX_REG_10__SCAN_IN;
  assign n7387 = ~PHYADDRPOINTER_REG_10__SCAN_IN | ~n8114;
  assign n7389 = ~n7388 | ~n7387;
  assign n7393 = ~n7390 & ~n7389;
  assign n11658 = PHYADDRPOINTER_REG_10__SCAN_IN ^ n7394;
  assign n7392 = ~n8628 | ~n11658;
  assign n10239 = ~n7393 | ~n7392;
  assign n7396 = ~n7751 | ~EAX_REG_11__SCAN_IN;
  assign n11691 = PHYADDRPOINTER_REG_11__SCAN_IN ^ ~n7463;
  assign n7395 = ~n8628 | ~n11691;
  assign n7431 = ~n7396 | ~n7395;
  assign n7429 = ~PHYADDRPOINTER_REG_11__SCAN_IN | ~n8114;
  assign n7398 = ~INSTQUEUE_REG_13__3__SCAN_IN | ~n6303;
  assign n7397 = ~INSTQUEUE_REG_9__3__SCAN_IN | ~n6302;
  assign n7400 = ~n7398 | ~n7397;
  assign n8041 = ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n7399 = ~n8719 & ~n8041;
  assign n7402 = ~n7400 & ~n7399;
  assign n7401 = ~n8188 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n7418 = ~n7402 | ~n7401;
  assign n7404 = ~n6295 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n7403 = ~n8178 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n7408 = ~n7404 | ~n7403;
  assign n7406 = ~INSTQUEUE_REG_7__3__SCAN_IN | ~n6292;
  assign n7405 = ~INSTQUEUE_REG_8__3__SCAN_IN | ~n8137;
  assign n7407 = ~n7406 | ~n7405;
  assign n7416 = ~n7408 & ~n7407;
  assign n7410 = ~INSTQUEUE_REG_1__3__SCAN_IN | ~n8162;
  assign n7409 = ~INSTQUEUE_REG_4__3__SCAN_IN | ~n8242;
  assign n7414 = ~n7410 | ~n7409;
  assign n7412 = ~INSTQUEUE_REG_6__3__SCAN_IN | ~n8187;
  assign n7411 = ~INSTQUEUE_REG_10__3__SCAN_IN | ~n7484;
  assign n7413 = ~n7412 | ~n7411;
  assign n7415 = ~n7414 & ~n7413;
  assign n7417 = ~n7416 | ~n7415;
  assign n7426 = ~n7418 & ~n7417;
  assign n7420 = ~n8138 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n7419 = ~n8118 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n7424 = ~n7420 | ~n7419;
  assign n7422 = ~INSTQUEUE_REG_12__3__SCAN_IN | ~n8119;
  assign n7421 = ~INSTQUEUE_REG_11__3__SCAN_IN | ~n8219;
  assign n7423 = ~n7422 | ~n7421;
  assign n7425 = ~n7424 & ~n7423;
  assign n7427 = ~n7426 | ~n7425;
  assign n7428 = ~n8260 | ~n7427;
  assign n7430 = ~n7429 | ~n7428;
  assign n10277 = ~n7431 & ~n7430;
  assign n7433 = ~n8188 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n7432 = ~n8233 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n7437 = ~n7433 | ~n7432;
  assign n7435 = ~n8122 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n7434 = ~n8137 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n7436 = ~n7435 | ~n7434;
  assign n7445 = ~n7437 & ~n7436;
  assign n7439 = ~INSTQUEUE_REG_6__4__SCAN_IN | ~n8187;
  assign n7438 = ~INSTQUEUE_REG_9__4__SCAN_IN | ~n6302;
  assign n7443 = ~n7439 | ~n7438;
  assign n7441 = ~INSTQUEUE_REG_12__4__SCAN_IN | ~n8119;
  assign n7440 = ~INSTQUEUE_REG_11__4__SCAN_IN | ~n8219;
  assign n7442 = ~n7441 | ~n7440;
  assign n7444 = ~n7443 & ~n7442;
  assign n7461 = ~n7445 | ~n7444;
  assign n7447 = ~n6303 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n7446 = ~n8178 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n7451 = ~n7447 | ~n7446;
  assign n7449 = ~INSTQUEUE_REG_1__4__SCAN_IN | ~n8162;
  assign n7448 = ~INSTQUEUE_REG_0__4__SCAN_IN | ~n8169;
  assign n7450 = ~n7449 | ~n7448;
  assign n7459 = ~n7451 & ~n7450;
  assign n7453 = ~INSTQUEUE_REG_3__4__SCAN_IN | ~n6294;
  assign n7452 = ~INSTQUEUE_REG_7__4__SCAN_IN | ~n6292;
  assign n7457 = ~n7453 | ~n7452;
  assign n7455 = ~n8138 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n7454 = ~n8118 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n7456 = ~n7455 | ~n7454;
  assign n7458 = ~n7457 & ~n7456;
  assign n7460 = ~n7459 | ~n7458;
  assign n7462 = ~n7461 & ~n7460;
  assign n7467 = ~n7580 & ~n7462;
  assign n7465 = ~n7751 | ~EAX_REG_12__SCAN_IN;
  assign n11967 = PHYADDRPOINTER_REG_12__SCAN_IN ^ n7502;
  assign n7464 = ~n8628 | ~n11967;
  assign n7466 = ~n7465 | ~n7464;
  assign n7469 = ~n7467 & ~n7466;
  assign n7468 = ~PHYADDRPOINTER_REG_12__SCAN_IN | ~n8114;
  assign n10501 = ~n7469 | ~n7468;
  assign n7471 = ~n8122 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n7470 = ~n8118 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n7473 = ~n7471 | ~n7470;
  assign n7472 = ~n8719 & ~n6710;
  assign n7475 = ~n7473 & ~n7472;
  assign n7474 = ~n6292 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n7492 = ~n7475 | ~n7474;
  assign n7477 = ~INSTQUEUE_REG_3__5__SCAN_IN | ~n6295;
  assign n7476 = ~INSTQUEUE_REG_1__5__SCAN_IN | ~n8162;
  assign n7481 = ~n7477 | ~n7476;
  assign n7479 = ~INSTQUEUE_REG_11__5__SCAN_IN | ~n8219;
  assign n7478 = ~INSTQUEUE_REG_15__5__SCAN_IN | ~n8222;
  assign n7480 = ~n7479 | ~n7478;
  assign n7490 = ~n7481 & ~n7480;
  assign n7483 = ~n8119 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n7482 = ~n8178 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n7488 = ~n7483 | ~n7482;
  assign n7486 = ~n7484 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n7485 = ~n6303 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n7487 = ~n7486 | ~n7485;
  assign n7489 = ~n7488 & ~n7487;
  assign n7491 = ~n7490 | ~n7489;
  assign n7500 = ~n7492 & ~n7491;
  assign n7494 = ~INSTQUEUE_REG_6__5__SCAN_IN | ~n8187;
  assign n7493 = ~INSTQUEUE_REG_8__5__SCAN_IN | ~n8182;
  assign n7498 = ~n7494 | ~n7493;
  assign n7496 = ~INSTQUEUE_REG_5__5__SCAN_IN | ~n8212;
  assign n7495 = ~INSTQUEUE_REG_9__5__SCAN_IN | ~n6299;
  assign n7497 = ~n7496 | ~n7495;
  assign n7499 = ~n7498 & ~n7497;
  assign n7501 = ~n7500 | ~n7499;
  assign n7508 = ~n8260 | ~n7501;
  assign n11155 = PHYADDRPOINTER_REG_13__SCAN_IN ^ n7511;
  assign n7506 = ~n11155 & ~n9025;
  assign n7504 = ~n7751 | ~EAX_REG_13__SCAN_IN;
  assign n7503 = ~PHYADDRPOINTER_REG_13__SCAN_IN | ~n8114;
  assign n7505 = ~n7504 | ~n7503;
  assign n8815 = ~n7506 & ~n7505;
  assign n7513 = ~n7751 | ~EAX_REG_14__SCAN_IN;
  assign n11818 = PHYADDRPOINTER_REG_14__SCAN_IN ^ n7581;
  assign n7512 = ~n8628 | ~n11818;
  assign n7548 = ~n7513 | ~n7512;
  assign n7515 = ~INSTQUEUE_REG_11__6__SCAN_IN | ~n8219;
  assign n7514 = ~INSTQUEUE_REG_15__6__SCAN_IN | ~n8222;
  assign n7517 = ~n7515 | ~n7514;
  assign n7516 = n8169 & INSTQUEUE_REG_0__6__SCAN_IN;
  assign n7519 = ~n7517 & ~n7516;
  assign n7518 = ~n8188 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n7535 = ~n7519 | ~n7518;
  assign n7521 = ~INSTQUEUE_REG_7__6__SCAN_IN | ~n6291;
  assign n7520 = ~INSTQUEUE_REG_8__6__SCAN_IN | ~n8137;
  assign n7525 = ~n7521 | ~n7520;
  assign n7523 = ~INSTQUEUE_REG_1__6__SCAN_IN | ~n8162;
  assign n7522 = ~INSTQUEUE_REG_4__6__SCAN_IN | ~n8242;
  assign n7524 = ~n7523 | ~n7522;
  assign n7533 = ~n7525 & ~n7524;
  assign n7527 = ~INSTQUEUE_REG_6__6__SCAN_IN | ~n8187;
  assign n7526 = ~INSTQUEUE_REG_10__6__SCAN_IN | ~n8233;
  assign n7531 = ~n7527 | ~n7526;
  assign n7529 = ~n6302 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n7528 = ~n8178 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n7530 = ~n7529 | ~n7528;
  assign n7532 = ~n7531 & ~n7530;
  assign n7534 = ~n7533 | ~n7532;
  assign n7543 = ~n7535 & ~n7534;
  assign n7537 = ~INSTQUEUE_REG_3__6__SCAN_IN | ~n6288;
  assign n7536 = ~INSTQUEUE_REG_13__6__SCAN_IN | ~n6303;
  assign n7541 = ~n7537 | ~n7536;
  assign n7539 = ~n8118 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n7538 = ~n8119 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n7540 = ~n7539 | ~n7538;
  assign n7542 = ~n7541 & ~n7540;
  assign n7544 = ~n7543 | ~n7542;
  assign n7546 = ~n8260 | ~n7544;
  assign n7545 = ~PHYADDRPOINTER_REG_14__SCAN_IN | ~n8114;
  assign n7547 = ~n7546 | ~n7545;
  assign n8821 = ~n7548 & ~n7547;
  assign n7550 = ~INSTQUEUE_REG_3__7__SCAN_IN | ~n6293;
  assign n7549 = ~INSTQUEUE_REG_9__7__SCAN_IN | ~n6300;
  assign n7554 = ~n7550 | ~n7549;
  assign n7552 = ~INSTQUEUE_REG_1__7__SCAN_IN | ~n8239;
  assign n7551 = ~INSTQUEUE_REG_11__7__SCAN_IN | ~n8219;
  assign n7553 = ~n7552 | ~n7551;
  assign n7562 = ~n7554 & ~n7553;
  assign n7556 = ~INSTQUEUE_REG_6__7__SCAN_IN | ~n8187;
  assign n7555 = ~INSTQUEUE_REG_10__7__SCAN_IN | ~n7484;
  assign n7560 = ~n7556 | ~n7555;
  assign n7558 = ~n6683 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n7557 = ~n8118 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n7559 = ~n7558 | ~n7557;
  assign n7561 = ~n7560 & ~n7559;
  assign n7578 = ~n7562 | ~n7561;
  assign n7564 = ~n8178 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n7563 = ~n8138 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n7568 = ~n7564 | ~n7563;
  assign n7566 = ~INSTQUEUE_REG_7__7__SCAN_IN | ~n6291;
  assign n7565 = ~INSTQUEUE_REG_5__7__SCAN_IN | ~n8212;
  assign n7567 = ~n7566 | ~n7565;
  assign n7576 = ~n7568 & ~n7567;
  assign n7570 = ~n8119 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n7569 = ~n8137 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n7574 = ~n7570 | ~n7569;
  assign n7572 = ~INSTQUEUE_REG_13__7__SCAN_IN | ~n6303;
  assign n7571 = ~INSTQUEUE_REG_4__7__SCAN_IN | ~n8242;
  assign n7573 = ~n7572 | ~n7571;
  assign n7575 = ~n7574 & ~n7573;
  assign n7577 = ~n7576 | ~n7575;
  assign n7579 = ~n7578 & ~n7577;
  assign n7585 = ~n7580 & ~n7579;
  assign n7583 = ~n7751 | ~EAX_REG_15__SCAN_IN;
  assign n12045 = PHYADDRPOINTER_REG_15__SCAN_IN ^ ~n7639;
  assign n7582 = ~n8628 | ~n12045;
  assign n7584 = ~n7583 | ~n7582;
  assign n7587 = ~n7585 & ~n7584;
  assign n7586 = ~PHYADDRPOINTER_REG_15__SCAN_IN | ~n8114;
  assign n11254 = ~n7587 | ~n7586;
  assign n7638 = ~n7751 | ~EAX_REG_16__SCAN_IN;
  assign n7600 = ~n7588;
  assign n7590 = ~n7589;
  assign n7592 = ~n7591 | ~n7590;
  assign n10867 = ~n9476 & ~n9821;
  assign n7599 = ~n7592 | ~n10867;
  assign n7594 = ~n7593 & ~n8429;
  assign n7595 = ~n7594 | ~n9821;
  assign n8383 = ~n7596 | ~n7595;
  assign n7597 = ~n8441 & ~n8378;
  assign n7598 = ~n8383 & ~n7597;
  assign n8438 = ~n7599 | ~n7598;
  assign n7604 = ~INSTQUEUE_REG_13__0__SCAN_IN | ~n8119;
  assign n7603 = ~INSTQUEUE_REG_14__0__SCAN_IN | ~n6303;
  assign n7608 = ~n7604 | ~n7603;
  assign n7606 = ~n8118 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n7605 = ~n8178 | ~INSTQUEUE_REG_3__0__SCAN_IN;
  assign n7607 = ~n7606 | ~n7605;
  assign n7616 = ~n7608 & ~n7607;
  assign n7610 = ~n8137 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n7609 = ~n8233 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n7614 = ~n7610 | ~n7609;
  assign n7612 = ~INSTQUEUE_REG_2__0__SCAN_IN | ~n8239;
  assign n7611 = ~INSTQUEUE_REG_6__0__SCAN_IN | ~n8212;
  assign n7613 = ~n7612 | ~n7611;
  assign n7615 = ~n7614 & ~n7613;
  assign n7632 = ~n7616 | ~n7615;
  assign n7618 = ~INSTQUEUE_REG_1__0__SCAN_IN | ~n8169;
  assign n7617 = ~INSTQUEUE_REG_10__0__SCAN_IN | ~n6302;
  assign n7622 = ~n7618 | ~n7617;
  assign n7620 = ~INSTQUEUE_REG_12__0__SCAN_IN | ~n8219;
  assign n7619 = ~INSTQUEUE_REG_0__0__SCAN_IN | ~n8222;
  assign n7621 = ~n7620 | ~n7619;
  assign n7630 = ~n7622 & ~n7621;
  assign n7624 = ~INSTQUEUE_REG_7__0__SCAN_IN | ~n8187;
  assign n7623 = ~INSTQUEUE_REG_5__0__SCAN_IN | ~n8242;
  assign n7628 = ~n7624 | ~n7623;
  assign n7626 = ~INSTQUEUE_REG_4__0__SCAN_IN | ~n6294;
  assign n7625 = ~INSTQUEUE_REG_8__0__SCAN_IN | ~n6291;
  assign n7627 = ~n7626 | ~n7625;
  assign n7629 = ~n7628 & ~n7627;
  assign n7631 = ~n7630 | ~n7629;
  assign n7633 = ~n7632 & ~n7631;
  assign n7636 = ~n8202 & ~n7633;
  assign n7634 = ~n11362 & ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n7635 = ~STATE2_REG_2__SCAN_IN & ~n7634;
  assign n7637 = ~n7636 & ~n7635;
  assign n7641 = ~n7638 | ~n7637;
  assign n12075 = PHYADDRPOINTER_REG_16__SCAN_IN ^ ~n7674;
  assign n7640 = ~n8628 | ~n12075;
  assign n11699 = ~n7641 | ~n7640;
  assign n7643 = ~n8118 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n7642 = ~INSTQUEUE_REG_12__1__SCAN_IN | ~n8219;
  assign n7647 = ~n7643 | ~n7642;
  assign n7645 = ~n6287 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n7644 = ~INSTQUEUE_REG_10__1__SCAN_IN | ~n6299;
  assign n7646 = ~n7645 | ~n7644;
  assign n7655 = ~n7647 & ~n7646;
  assign n7649 = ~INSTQUEUE_REG_8__1__SCAN_IN | ~n6291;
  assign n7648 = ~n8212 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n7653 = ~n7649 | ~n7648;
  assign n7651 = ~n8122 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n7650 = ~INSTQUEUE_REG_1__1__SCAN_IN | ~n8169;
  assign n7652 = ~n7651 | ~n7650;
  assign n7654 = ~n7653 & ~n7652;
  assign n7671 = ~n7655 | ~n7654;
  assign n7657 = ~INSTQUEUE_REG_4__1__SCAN_IN | ~n6293;
  assign n7656 = ~n8138 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n7661 = ~n7657 | ~n7656;
  assign n7659 = ~n8162 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n7658 = ~n8178 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n7660 = ~n7659 | ~n7658;
  assign n7669 = ~n7661 & ~n7660;
  assign n7663 = ~n8119 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n7662 = ~n8187 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n7667 = ~n7663 | ~n7662;
  assign n7665 = ~INSTQUEUE_REG_9__1__SCAN_IN | ~n8182;
  assign n7664 = ~INSTQUEUE_REG_11__1__SCAN_IN | ~n6298;
  assign n7666 = ~n7665 | ~n7664;
  assign n7668 = ~n7667 & ~n7666;
  assign n7670 = ~n7669 | ~n7668;
  assign n7672 = ~n7671 & ~n7670;
  assign n7678 = ~n8202 & ~n7672;
  assign n7676 = ~n7751 | ~EAX_REG_17__SCAN_IN;
  assign n7673 = ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n12095 = PHYADDRPOINTER_REG_17__SCAN_IN ^ ~n7681;
  assign n7675 = ~n8628 | ~n12095;
  assign n7677 = ~n7676 | ~n7675;
  assign n7680 = ~n7678 & ~n7677;
  assign n7679 = ~PHYADDRPOINTER_REG_17__SCAN_IN | ~n8550;
  assign n11746 = ~n7680 | ~n7679;
  assign n11875 = ~n11747 | ~n11746;
  assign n7683 = ~n7751 | ~EAX_REG_18__SCAN_IN;
  assign n7757 = ~PHYADDRPOINTER_REG_17__SCAN_IN | ~n7681;
  assign n12177 = PHYADDRPOINTER_REG_18__SCAN_IN ^ n7757;
  assign n7682 = ~n8628 | ~n12177;
  assign n7719 = ~n7683 | ~n7682;
  assign n7717 = ~PHYADDRPOINTER_REG_18__SCAN_IN | ~n8114;
  assign n7685 = ~INSTQUEUE_REG_14__2__SCAN_IN | ~n6303;
  assign n7684 = ~INSTQUEUE_REG_12__2__SCAN_IN | ~n8219;
  assign n7688 = ~n7685 | ~n7684;
  assign n7687 = ~n7801 & ~n7686;
  assign n7690 = ~n7688 & ~n7687;
  assign n7689 = ~n8233 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n7706 = ~n7690 | ~n7689;
  assign n7692 = ~INSTQUEUE_REG_7__2__SCAN_IN | ~n8187;
  assign n7691 = ~INSTQUEUE_REG_2__2__SCAN_IN | ~n8239;
  assign n7696 = ~n7692 | ~n7691;
  assign n7694 = ~INSTQUEUE_REG_5__2__SCAN_IN | ~n8242;
  assign n7693 = ~INSTQUEUE_REG_10__2__SCAN_IN | ~n6301;
  assign n7695 = ~n7694 | ~n7693;
  assign n7704 = ~n7696 & ~n7695;
  assign n7698 = ~n8119 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n7697 = ~n8137 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n7702 = ~n7698 | ~n7697;
  assign n7700 = ~INSTQUEUE_REG_8__2__SCAN_IN | ~n6292;
  assign n7699 = ~INSTQUEUE_REG_1__2__SCAN_IN | ~n8169;
  assign n7701 = ~n7700 | ~n7699;
  assign n7703 = ~n7702 & ~n7701;
  assign n7705 = ~n7704 | ~n7703;
  assign n7714 = ~n7706 & ~n7705;
  assign n7708 = ~n8118 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n7707 = ~n8212 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n7712 = ~n7708 | ~n7707;
  assign n7710 = ~n6294 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n7709 = ~n8178 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n7711 = ~n7710 | ~n7709;
  assign n7713 = ~n7712 & ~n7711;
  assign n7715 = ~n7714 | ~n7713;
  assign n7716 = ~n8253 | ~n7715;
  assign n7718 = ~n7717 | ~n7716;
  assign n11914 = ~n11875 & ~n11876;
  assign n7721 = ~INSTQUEUE_REG_1__3__SCAN_IN | ~n8169;
  assign n7720 = ~INSTQUEUE_REG_12__3__SCAN_IN | ~n8219;
  assign n7723 = ~n7721 | ~n7720;
  assign n7722 = ~n7801 & ~n8041;
  assign n7725 = ~n7723 & ~n7722;
  assign n7724 = ~n8118 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n7741 = ~n7725 | ~n7724;
  assign n7727 = ~n8233 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n7726 = ~n6293 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n7731 = ~n7727 | ~n7726;
  assign n7729 = ~INSTQUEUE_REG_5__3__SCAN_IN | ~n8242;
  assign n7728 = ~INSTQUEUE_REG_9__3__SCAN_IN | ~n8137;
  assign n7730 = ~n7729 | ~n7728;
  assign n7739 = ~n7731 & ~n7730;
  assign n7733 = ~INSTQUEUE_REG_3__3__SCAN_IN | ~n8178;
  assign n7732 = ~INSTQUEUE_REG_8__3__SCAN_IN | ~n6291;
  assign n7737 = ~n7733 | ~n7732;
  assign n7735 = ~INSTQUEUE_REG_13__3__SCAN_IN | ~n8119;
  assign n7734 = ~INSTQUEUE_REG_2__3__SCAN_IN | ~n8239;
  assign n7736 = ~n7735 | ~n7734;
  assign n7738 = ~n7737 & ~n7736;
  assign n7740 = ~n7739 | ~n7738;
  assign n7749 = ~n7741 & ~n7740;
  assign n7743 = ~INSTQUEUE_REG_7__3__SCAN_IN | ~n8187;
  assign n7742 = ~INSTQUEUE_REG_10__3__SCAN_IN | ~n6299;
  assign n7747 = ~n7743 | ~n7742;
  assign n7745 = ~INSTQUEUE_REG_14__3__SCAN_IN | ~n6287;
  assign n7744 = ~INSTQUEUE_REG_6__3__SCAN_IN | ~n8212;
  assign n7746 = ~n7745 | ~n7744;
  assign n7748 = ~n7747 & ~n7746;
  assign n7750 = ~n7749 | ~n7748;
  assign n7753 = ~n8253 | ~n7750;
  assign n7752 = ~n7751 | ~EAX_REG_19__SCAN_IN;
  assign n7756 = ~n7753 | ~n7752;
  assign n7754 = ~PHYADDRPOINTER_REG_19__SCAN_IN & ~n11362;
  assign n7755 = ~STATE2_REG_2__SCAN_IN & ~n7754;
  assign n7759 = ~n7756 & ~n7755;
  assign n11940 = ~PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n12118 = PHYADDRPOINTER_REG_19__SCAN_IN ^ ~n7796;
  assign n7758 = ~n12118 & ~n9025;
  assign n11913 = ~n7759 & ~n7758;
  assign n7795 = ~EAX_REG_20__SCAN_IN | ~n7751;
  assign n7761 = ~INSTQUEUE_REG_13__4__SCAN_IN | ~n8119;
  assign n7760 = ~INSTQUEUE_REG_12__4__SCAN_IN | ~n8219;
  assign n7765 = ~n7761 | ~n7760;
  assign n7762 = ~INSTQUEUE_REG_7__4__SCAN_IN | ~n8187;
  assign n7764 = ~n7763 | ~n7762;
  assign n7773 = ~n7765 & ~n7764;
  assign n7767 = ~n8137 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n7766 = ~n8178 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n7771 = ~n7767 | ~n7766;
  assign n7769 = ~INSTQUEUE_REG_15__4__SCAN_IN | ~n8238;
  assign n7768 = ~INSTQUEUE_REG_1__4__SCAN_IN | ~n8169;
  assign n7770 = ~n7769 | ~n7768;
  assign n7772 = ~n7771 & ~n7770;
  assign n7789 = ~n7773 | ~n7772;
  assign n7775 = ~n7484 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n7774 = ~n6300 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n7779 = ~n7775 | ~n7774;
  assign n7777 = ~INSTQUEUE_REG_14__4__SCAN_IN | ~n6303;
  assign n7776 = ~INSTQUEUE_REG_2__4__SCAN_IN | ~n8239;
  assign n7778 = ~n7777 | ~n7776;
  assign n7787 = ~n7779 & ~n7778;
  assign n7781 = ~INSTQUEUE_REG_5__4__SCAN_IN | ~n8242;
  assign n7780 = ~INSTQUEUE_REG_8__4__SCAN_IN | ~n6291;
  assign n7785 = ~n7781 | ~n7780;
  assign n7783 = ~n8138 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n7782 = ~n8212 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n7784 = ~n7783 | ~n7782;
  assign n7786 = ~n7785 & ~n7784;
  assign n7788 = ~n7787 | ~n7786;
  assign n7790 = ~n7789 & ~n7788;
  assign n7793 = ~n8202 & ~n7790;
  assign n7791 = ~n11362 & ~PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n7792 = ~STATE2_REG_2__SCAN_IN & ~n7791;
  assign n7794 = ~n7793 & ~n7792;
  assign n7798 = ~n7795 | ~n7794;
  assign n12272 = PHYADDRPOINTER_REG_20__SCAN_IN ^ n7836;
  assign n7797 = ~n8628 | ~n12272;
  assign n8862 = ~n7798 | ~n7797;
  assign n7800 = ~INSTQUEUE_REG_14__5__SCAN_IN | ~n6303;
  assign n7799 = ~INSTQUEUE_REG_5__5__SCAN_IN | ~n8242;
  assign n7803 = ~n7800 | ~n7799;
  assign n7802 = ~n7801 & ~n6710;
  assign n7805 = ~n7803 & ~n7802;
  assign n7804 = ~n8118 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n7821 = ~n7805 | ~n7804;
  assign n7807 = ~INSTQUEUE_REG_13__5__SCAN_IN | ~n8119;
  assign n7806 = ~INSTQUEUE_REG_2__5__SCAN_IN | ~n8162;
  assign n7811 = ~n7807 | ~n7806;
  assign n7809 = ~n6302 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n7808 = ~n6294 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n7810 = ~n7809 | ~n7808;
  assign n7819 = ~n7811 & ~n7810;
  assign n7813 = ~INSTQUEUE_REG_7__5__SCAN_IN | ~n8187;
  assign n7812 = ~INSTQUEUE_REG_11__5__SCAN_IN | ~n6298;
  assign n7817 = ~n7813 | ~n7812;
  assign n7815 = ~n6291 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n7814 = ~n8212 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n7816 = ~n7815 | ~n7814;
  assign n7818 = ~n7817 & ~n7816;
  assign n7820 = ~n7819 | ~n7818;
  assign n7829 = ~n7821 & ~n7820;
  assign n7823 = ~INSTQUEUE_REG_3__5__SCAN_IN | ~n8178;
  assign n7822 = ~INSTQUEUE_REG_12__5__SCAN_IN | ~n8219;
  assign n7827 = ~n7823 | ~n7822;
  assign n7825 = ~INSTQUEUE_REG_1__5__SCAN_IN | ~n8169;
  assign n7824 = ~INSTQUEUE_REG_9__5__SCAN_IN | ~n8182;
  assign n7826 = ~n7825 | ~n7824;
  assign n7828 = ~n7827 & ~n7826;
  assign n7830 = ~n7829 | ~n7828;
  assign n7832 = ~n8253 | ~n7830;
  assign n7831 = ~n7751 | ~EAX_REG_21__SCAN_IN;
  assign n7835 = ~n7832 | ~n7831;
  assign n7833 = ~PHYADDRPOINTER_REG_21__SCAN_IN & ~n11362;
  assign n7834 = ~STATE2_REG_2__SCAN_IN & ~n7833;
  assign n7838 = ~n7835 & ~n7834;
  assign n12340 = PHYADDRPOINTER_REG_21__SCAN_IN ^ ~n7875;
  assign n7837 = ~n9025 & ~n12340;
  assign n8834 = ~n7838 & ~n7837;
  assign n7874 = ~EAX_REG_22__SCAN_IN | ~n7751;
  assign n7840 = ~INSTQUEUE_REG_3__6__SCAN_IN | ~n8178;
  assign n7839 = ~INSTQUEUE_REG_12__6__SCAN_IN | ~n8219;
  assign n7844 = ~n7840 | ~n7839;
  assign n7842 = ~n6298 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n7841 = ~n8169 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n7843 = ~n7842 | ~n7841;
  assign n7852 = ~n7844 & ~n7843;
  assign n7846 = ~INSTQUEUE_REG_2__6__SCAN_IN | ~n8239;
  assign n7845 = ~INSTQUEUE_REG_6__6__SCAN_IN | ~n8212;
  assign n7850 = ~n7846 | ~n7845;
  assign n7848 = ~INSTQUEUE_REG_4__6__SCAN_IN | ~n6288;
  assign n7847 = ~INSTQUEUE_REG_10__6__SCAN_IN | ~n6300;
  assign n7849 = ~n7848 | ~n7847;
  assign n7851 = ~n7850 & ~n7849;
  assign n7868 = ~n7852 | ~n7851;
  assign n7854 = ~n8122 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n7853 = ~n8118 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n7858 = ~n7854 | ~n7853;
  assign n7856 = ~INSTQUEUE_REG_14__6__SCAN_IN | ~n6303;
  assign n7855 = ~INSTQUEUE_REG_8__6__SCAN_IN | ~n6291;
  assign n7857 = ~n7856 | ~n7855;
  assign n7866 = ~n7858 & ~n7857;
  assign n7860 = ~INSTQUEUE_REG_7__6__SCAN_IN | ~n8187;
  assign n7859 = ~INSTQUEUE_REG_0__6__SCAN_IN | ~n8222;
  assign n7864 = ~n7860 | ~n7859;
  assign n7862 = ~n8119 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n7861 = ~n8137 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n7863 = ~n7862 | ~n7861;
  assign n7865 = ~n7864 & ~n7863;
  assign n7867 = ~n7866 | ~n7865;
  assign n7869 = ~n7868 & ~n7867;
  assign n7872 = ~n8202 & ~n7869;
  assign n7870 = ~n11362 & ~PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n7871 = ~STATE2_REG_2__SCAN_IN & ~n7870;
  assign n7873 = ~n7872 & ~n7871;
  assign n7877 = ~n7874 | ~n7873;
  assign n12359 = PHYADDRPOINTER_REG_22__SCAN_IN ^ n7939;
  assign n7876 = ~n8628 | ~n12359;
  assign n8848 = ~n7877 | ~n7876;
  assign n7879 = ~INSTQUEUE_REG_0__0__SCAN_IN | ~n8238;
  assign n7878 = ~INSTQUEUE_REG_15__0__SCAN_IN | ~n6303;
  assign n7883 = ~n7879 | ~n7878;
  assign n7881 = ~INSTQUEUE_REG_14__0__SCAN_IN | ~n8119;
  assign n7880 = ~INSTQUEUE_REG_13__0__SCAN_IN | ~n8219;
  assign n7882 = ~n7881 | ~n7880;
  assign n7891 = ~n7883 & ~n7882;
  assign n7885 = ~INSTQUEUE_REG_2__0__SCAN_IN | ~n8169;
  assign n7884 = ~INSTQUEUE_REG_11__0__SCAN_IN | ~n6299;
  assign n7889 = ~n7885 | ~n7884;
  assign n7887 = ~n6288 | ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n7886 = ~n8138 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n7888 = ~n7887 | ~n7886;
  assign n7890 = ~n7889 & ~n7888;
  assign n7907 = ~n7891 | ~n7890;
  assign n7893 = ~INSTQUEUE_REG_8__0__SCAN_IN | ~n8187;
  assign n7892 = ~INSTQUEUE_REG_7__0__SCAN_IN | ~n8212;
  assign n7897 = ~n7893 | ~n7892;
  assign n7895 = ~INSTQUEUE_REG_3__0__SCAN_IN | ~n8239;
  assign n7894 = ~INSTQUEUE_REG_6__0__SCAN_IN | ~n8242;
  assign n7896 = ~n7895 | ~n7894;
  assign n7905 = ~n7897 & ~n7896;
  assign n7899 = ~n8137 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n7898 = ~n8233 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n7903 = ~n7899 | ~n7898;
  assign n7901 = ~INSTQUEUE_REG_4__0__SCAN_IN | ~n8178;
  assign n7900 = ~INSTQUEUE_REG_9__0__SCAN_IN | ~n6292;
  assign n7902 = ~n7901 | ~n7900;
  assign n7904 = ~n7903 & ~n7902;
  assign n7906 = ~n7905 | ~n7904;
  assign n7981 = ~n7907 & ~n7906;
  assign n7909 = ~n6288 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n7908 = ~n8119 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n7913 = ~n7909 | ~n7908;
  assign n7911 = ~INSTQUEUE_REG_8__7__SCAN_IN | ~n6292;
  assign n7910 = ~INSTQUEUE_REG_10__7__SCAN_IN | ~n6300;
  assign n7912 = ~n7911 | ~n7910;
  assign n7921 = ~n7913 & ~n7912;
  assign n7915 = ~n8122 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n7914 = ~n8137 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n7919 = ~n7915 | ~n7914;
  assign n7917 = ~INSTQUEUE_REG_3__7__SCAN_IN | ~n8178;
  assign n7916 = ~INSTQUEUE_REG_1__7__SCAN_IN | ~n8169;
  assign n7918 = ~n7917 | ~n7916;
  assign n7920 = ~n7919 & ~n7918;
  assign n7937 = ~n7921 | ~n7920;
  assign n7923 = ~INSTQUEUE_REG_6__7__SCAN_IN | ~n8212;
  assign n7922 = ~INSTQUEUE_REG_12__7__SCAN_IN | ~n8219;
  assign n7927 = ~n7923 | ~n7922;
  assign n7925 = ~INSTQUEUE_REG_7__7__SCAN_IN | ~n8187;
  assign n7924 = ~INSTQUEUE_REG_0__7__SCAN_IN | ~n8222;
  assign n7926 = ~n7925 | ~n7924;
  assign n7935 = ~n7927 & ~n7926;
  assign n7929 = ~INSTQUEUE_REG_15__7__SCAN_IN | ~n8238;
  assign n7928 = ~INSTQUEUE_REG_14__7__SCAN_IN | ~n6303;
  assign n7933 = ~n7929 | ~n7928;
  assign n7931 = ~n8162 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n7930 = ~n8233 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n7932 = ~n7931 | ~n7930;
  assign n7934 = ~n7933 & ~n7932;
  assign n7936 = ~n7935 | ~n7934;
  assign n7982 = ~n7937 & ~n7936;
  assign n7938 = n7981 ^ ~n7982;
  assign n7943 = ~n8202 & ~n7938;
  assign n7941 = ~PHYADDRPOINTER_REG_23__SCAN_IN | ~n8550;
  assign n12420 = PHYADDRPOINTER_REG_23__SCAN_IN ^ ~n7946;
  assign n7940 = ~n8628 | ~n12420;
  assign n7942 = ~n7941 | ~n7940;
  assign n7945 = ~n7943 & ~n7942;
  assign n7944 = ~n7751 | ~EAX_REG_23__SCAN_IN;
  assign n8878 = ~n7945 | ~n7944;
  assign n8940 = ~n8879 | ~n8878;
  assign n7948 = ~PHYADDRPOINTER_REG_24__SCAN_IN | ~n8114;
  assign n12457 = PHYADDRPOINTER_REG_24__SCAN_IN ^ n8027;
  assign n7947 = ~n8628 | ~n12457;
  assign n7987 = ~n7948 | ~n7947;
  assign n7950 = ~n6303 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n7949 = ~n6288 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n7955 = ~n7950 | ~n7949;
  assign n7953 = ~n8162 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n7952 = ~n7951 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n7954 = ~n7953 | ~n7952;
  assign n7980 = ~n7955 & ~n7954;
  assign n7957 = ~n6301 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n7956 = ~n8178 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n7960 = ~n7957 | ~n7956;
  assign n7959 = ~n7958 & ~n8042;
  assign n7962 = ~n7960 & ~n7959;
  assign n7961 = ~n8138 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n7978 = ~n7962 | ~n7961;
  assign n7964 = ~n8233 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n7963 = ~n8169 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n7968 = ~n7964 | ~n7963;
  assign n7966 = ~INSTQUEUE_REG_10__1__SCAN_IN | ~n8137;
  assign n7965 = ~n6291 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n7967 = ~n7966 | ~n7965;
  assign n7976 = ~n7968 & ~n7967;
  assign n7970 = ~n8187 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n7969 = ~n8122 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n7974 = ~n7970 | ~n7969;
  assign n7972 = ~INSTQUEUE_REG_14__1__SCAN_IN | ~n8119;
  assign n7971 = ~INSTQUEUE_REG_7__1__SCAN_IN | ~n8212;
  assign n7973 = ~n7972 | ~n7971;
  assign n7975 = ~n7974 & ~n7973;
  assign n7977 = ~n7976 | ~n7975;
  assign n7979 = ~n7978 & ~n7977;
  assign n8019 = ~n7980 | ~n7979;
  assign n8020 = ~n7982 & ~n7981;
  assign n7983 = n8019 ^ n8020;
  assign n7985 = ~n7983 | ~n8253;
  assign n7984 = ~EAX_REG_24__SCAN_IN | ~n7751;
  assign n7986 = ~n7985 | ~n7984;
  assign n8522 = ~n8940 & ~n8941;
  assign n7989 = ~INSTQUEUE_REG_15__2__SCAN_IN | ~n6303;
  assign n7988 = ~INSTQUEUE_REG_11__2__SCAN_IN | ~n6299;
  assign n7993 = ~n7989 | ~n7988;
  assign n7991 = ~n8138 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n7990 = ~n8119 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n7992 = ~n7991 | ~n7990;
  assign n8002 = ~n7993 & ~n7992;
  assign n7995 = ~INSTQUEUE_REG_3__2__SCAN_IN | ~n8239;
  assign n7994 = ~INSTQUEUE_REG_6__2__SCAN_IN | ~n8242;
  assign n8000 = ~n7995 | ~n7994;
  assign n7998 = ~n7484 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n7997 = ~n6291 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n7999 = ~n7998 | ~n7997;
  assign n8001 = ~n8000 & ~n7999;
  assign n8018 = ~n8002 | ~n8001;
  assign n8004 = ~INSTQUEUE_REG_4__2__SCAN_IN | ~n8178;
  assign n8003 = ~INSTQUEUE_REG_13__2__SCAN_IN | ~n8219;
  assign n8008 = ~n8004 | ~n8003;
  assign n8006 = ~INSTQUEUE_REG_0__2__SCAN_IN | ~n8118;
  assign n8005 = ~INSTQUEUE_REG_2__2__SCAN_IN | ~n8169;
  assign n8007 = ~n8006 | ~n8005;
  assign n8016 = ~n8008 & ~n8007;
  assign n8010 = ~n8212 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n8009 = ~n8137 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n8014 = ~n8010 | ~n8009;
  assign n8012 = ~INSTQUEUE_REG_5__2__SCAN_IN | ~n6294;
  assign n8011 = ~INSTQUEUE_REG_8__2__SCAN_IN | ~n8187;
  assign n8013 = ~n8012 | ~n8011;
  assign n8015 = ~n8014 & ~n8013;
  assign n8017 = ~n8016 | ~n8015;
  assign n8066 = ~n8018 & ~n8017;
  assign n8065 = ~n8020 | ~n8019;
  assign n8021 = n8066 ^ n8065;
  assign n8023 = ~n8021 | ~n8253;
  assign n8022 = ~EAX_REG_25__SCAN_IN | ~n7751;
  assign n8026 = ~n8023 | ~n8022;
  assign n8024 = ~PHYADDRPOINTER_REG_25__SCAN_IN & ~n11362;
  assign n8025 = ~STATE2_REG_2__SCAN_IN & ~n8024;
  assign n8029 = ~n8026 & ~n8025;
  assign n12128 = ~PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n12147 = PHYADDRPOINTER_REG_25__SCAN_IN ^ ~n8030;
  assign n8028 = ~n9025 & ~n12147;
  assign n8523 = ~n8029 & ~n8028;
  assign n8032 = ~PHYADDRPOINTER_REG_26__SCAN_IN | ~n8550;
  assign n8111 = ~n8030 | ~PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n12353 = PHYADDRPOINTER_REG_26__SCAN_IN ^ n8111;
  assign n8031 = ~n8628 | ~n12353;
  assign n8071 = ~n8032 | ~n8031;
  assign n8034 = ~INSTQUEUE_REG_14__3__SCAN_IN | ~n8119;
  assign n8033 = ~INSTQUEUE_REG_11__3__SCAN_IN | ~n6302;
  assign n8038 = ~n8034 | ~n8033;
  assign n8036 = ~n8242 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n8035 = ~n8178 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n8037 = ~n8036 | ~n8035;
  assign n8064 = ~n8038 & ~n8037;
  assign n8040 = ~INSTQUEUE_REG_2__3__SCAN_IN | ~n8169;
  assign n8039 = ~INSTQUEUE_REG_10__3__SCAN_IN | ~n8137;
  assign n8044 = ~n8040 | ~n8039;
  assign n8043 = ~n8042 & ~n8041;
  assign n8046 = ~n8044 & ~n8043;
  assign n8045 = ~n8222 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n8062 = ~n8046 | ~n8045;
  assign n8048 = ~INSTQUEUE_REG_5__3__SCAN_IN | ~n6295;
  assign n8047 = ~INSTQUEUE_REG_3__3__SCAN_IN | ~n8239;
  assign n8052 = ~n8048 | ~n8047;
  assign n8050 = ~INSTQUEUE_REG_8__3__SCAN_IN | ~n8187;
  assign n8049 = ~INSTQUEUE_REG_9__3__SCAN_IN | ~n6291;
  assign n8051 = ~n8050 | ~n8049;
  assign n8060 = ~n8052 & ~n8051;
  assign n8054 = ~n8233 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n8053 = ~n8212 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n8058 = ~n8054 | ~n8053;
  assign n8056 = ~INSTQUEUE_REG_15__3__SCAN_IN | ~n6303;
  assign n8055 = ~INSTQUEUE_REG_13__3__SCAN_IN | ~n8219;
  assign n8057 = ~n8056 | ~n8055;
  assign n8059 = ~n8058 & ~n8057;
  assign n8061 = ~n8060 | ~n8059;
  assign n8063 = ~n8062 & ~n8061;
  assign n8103 = ~n8064 | ~n8063;
  assign n8104 = ~n8066 & ~n8065;
  assign n8067 = n8103 ^ n8104;
  assign n8069 = ~n8067 | ~n8253;
  assign n8068 = ~EAX_REG_26__SCAN_IN | ~n7751;
  assign n8070 = ~n8069 | ~n8068;
  assign n8073 = ~INSTQUEUE_REG_3__4__SCAN_IN | ~n8239;
  assign n8072 = ~INSTQUEUE_REG_10__4__SCAN_IN | ~n8137;
  assign n8077 = ~n8073 | ~n8072;
  assign n8075 = ~n8122 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n8074 = ~n6294 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n8076 = ~n8075 | ~n8074;
  assign n8086 = ~n8077 & ~n8076;
  assign n8080 = ~n8212 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n8079 = ~n8178 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n8084 = ~n8080 | ~n8079;
  assign n8082 = ~INSTQUEUE_REG_13__4__SCAN_IN | ~n8219;
  assign n8081 = ~INSTQUEUE_REG_11__4__SCAN_IN | ~n6301;
  assign n8083 = ~n8082 | ~n8081;
  assign n8085 = ~n8084 & ~n8083;
  assign n8102 = ~n8086 | ~n8085;
  assign n8088 = ~n7484 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n8087 = ~n8119 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n8092 = ~n8088 | ~n8087;
  assign n8090 = ~n6303 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n8089 = ~n8222 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n8091 = ~n8090 | ~n8089;
  assign n8100 = ~n8092 & ~n8091;
  assign n8094 = ~INSTQUEUE_REG_0__4__SCAN_IN | ~n8238;
  assign n8093 = ~INSTQUEUE_REG_2__4__SCAN_IN | ~n8169;
  assign n8098 = ~n8094 | ~n8093;
  assign n8096 = ~INSTQUEUE_REG_8__4__SCAN_IN | ~n8187;
  assign n8095 = ~INSTQUEUE_REG_9__4__SCAN_IN | ~n6292;
  assign n8097 = ~n8096 | ~n8095;
  assign n8099 = ~n8098 & ~n8097;
  assign n8101 = ~n8100 | ~n8099;
  assign n8154 = ~n8102 & ~n8101;
  assign n8153 = ~n8104 | ~n8103;
  assign n8105 = n8154 ^ n8153;
  assign n8107 = ~n8105 | ~n8253;
  assign n8106 = ~EAX_REG_27__SCAN_IN | ~n7751;
  assign n8110 = ~n8107 | ~n8106;
  assign n8108 = ~PHYADDRPOINTER_REG_27__SCAN_IN & ~n11362;
  assign n8109 = ~STATE2_REG_2__SCAN_IN & ~n8108;
  assign n8113 = ~n8110 & ~n8109;
  assign n12346 = ~PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n12380 = PHYADDRPOINTER_REG_27__SCAN_IN ^ n8115;
  assign n8112 = ~n9025 & ~n12380;
  assign n12166 = ~n8113 & ~n8112;
  assign n8117 = ~PHYADDRPOINTER_REG_28__SCAN_IN | ~n8114;
  assign n12255 = ~PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n12313 = PHYADDRPOINTER_REG_28__SCAN_IN ^ ~n8208;
  assign n8116 = ~n8628 | ~n12313;
  assign n8159 = ~n8117 | ~n8116;
  assign n8121 = ~n8118 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n8120 = ~n8119 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n8126 = ~n8121 | ~n8120;
  assign n8124 = ~n8122 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n8123 = ~n6288 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n8125 = ~n8124 | ~n8123;
  assign n8134 = ~n8126 & ~n8125;
  assign n8128 = ~INSTQUEUE_REG_8__5__SCAN_IN | ~n8187;
  assign n8127 = ~INSTQUEUE_REG_7__5__SCAN_IN | ~n8212;
  assign n8132 = ~n8128 | ~n8127;
  assign n8130 = ~INSTQUEUE_REG_15__5__SCAN_IN | ~n6303;
  assign n8129 = ~INSTQUEUE_REG_2__5__SCAN_IN | ~n8169;
  assign n8131 = ~n8130 | ~n8129;
  assign n8133 = ~n8132 & ~n8131;
  assign n8152 = ~n8134 | ~n8133;
  assign n8136 = ~INSTQUEUE_REG_4__5__SCAN_IN | ~n8178;
  assign n8135 = ~INSTQUEUE_REG_13__5__SCAN_IN | ~n8219;
  assign n8142 = ~n8136 | ~n8135;
  assign n8140 = ~n8137 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n8139 = ~n8138 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n8141 = ~n8140 | ~n8139;
  assign n8150 = ~n8142 & ~n8141;
  assign n8144 = ~INSTQUEUE_REG_9__5__SCAN_IN | ~n6291;
  assign n8143 = ~INSTQUEUE_REG_11__5__SCAN_IN | ~n6300;
  assign n8148 = ~n8144 | ~n8143;
  assign n8146 = ~n8162 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n8145 = ~n8233 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n8147 = ~n8146 | ~n8145;
  assign n8149 = ~n8148 & ~n8147;
  assign n8151 = ~n8150 | ~n8149;
  assign n8199 = ~n8152 & ~n8151;
  assign n8200 = n8154 | n8153;
  assign n8155 = n8199 ^ n8200;
  assign n8157 = ~n8155 | ~n8253;
  assign n8156 = ~EAX_REG_28__SCAN_IN | ~n7751;
  assign n8158 = ~n8157 | ~n8156;
  assign n8621 = ~n8159 & ~n8158;
  assign n8207 = ~EAX_REG_29__SCAN_IN | ~n7751;
  assign n8164 = ~INSTQUEUE_REG_3__6__SCAN_IN | ~n8162;
  assign n8163 = ~INSTQUEUE_REG_11__6__SCAN_IN | ~n6302;
  assign n8168 = ~n8164 | ~n8163;
  assign n8166 = ~INSTQUEUE_REG_14__6__SCAN_IN | ~n8119;
  assign n8165 = ~INSTQUEUE_REG_13__6__SCAN_IN | ~n8219;
  assign n8167 = ~n8166 | ~n8165;
  assign n8177 = ~n8168 & ~n8167;
  assign n8171 = ~INSTQUEUE_REG_12__6__SCAN_IN | ~n6298;
  assign n8170 = ~INSTQUEUE_REG_2__6__SCAN_IN | ~n8169;
  assign n8175 = ~n8171 | ~n8170;
  assign n8173 = ~INSTQUEUE_REG_5__6__SCAN_IN | ~n6295;
  assign n8172 = ~INSTQUEUE_REG_0__6__SCAN_IN | ~n8238;
  assign n8174 = ~n8173 | ~n8172;
  assign n8176 = ~n8175 & ~n8174;
  assign n8198 = ~n8177 | ~n8176;
  assign n8180 = ~INSTQUEUE_REG_4__6__SCAN_IN | ~n8178;
  assign n8179 = ~INSTQUEUE_REG_15__6__SCAN_IN | ~n6287;
  assign n8186 = ~n8180 | ~n8179;
  assign n8184 = ~INSTQUEUE_REG_9__6__SCAN_IN | ~n6291;
  assign n8183 = ~INSTQUEUE_REG_10__6__SCAN_IN | ~n8182;
  assign n8185 = ~n8184 | ~n8183;
  assign n8196 = ~n8186 & ~n8185;
  assign n8190 = ~INSTQUEUE_REG_8__6__SCAN_IN | ~n8187;
  assign n8189 = ~INSTQUEUE_REG_7__6__SCAN_IN | ~n8188;
  assign n8194 = ~n8190 | ~n8189;
  assign n8192 = ~INSTQUEUE_REG_6__6__SCAN_IN | ~n8242;
  assign n8191 = ~INSTQUEUE_REG_1__6__SCAN_IN | ~n8222;
  assign n8193 = ~n8192 | ~n8191;
  assign n8195 = ~n8194 & ~n8193;
  assign n8197 = ~n8196 | ~n8195;
  assign n8251 = n8198 | n8197;
  assign n8252 = ~n8200 & ~n8199;
  assign n8201 = n8251 ^ ~n8252;
  assign n8205 = ~n8202 & ~n8201;
  assign n8203 = ~n11362 & ~PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n8204 = ~STATE2_REG_2__SCAN_IN & ~n8203;
  assign n8206 = ~n8205 & ~n8204;
  assign n8210 = ~n8207 | ~n8206;
  assign n8266 = ~n8208 | ~PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n12432 = PHYADDRPOINTER_REG_29__SCAN_IN ^ ~n8266;
  assign n8209 = ~n8628 | ~n12432;
  assign n8546 = ~n8210 | ~n8209;
  assign n8211 = ~PHYADDRPOINTER_REG_30__SCAN_IN & ~n11362;
  assign n8256 = ~STATE2_REG_2__SCAN_IN & ~n8211;
  assign n8214 = ~INSTQUEUE_REG_7__7__SCAN_IN | ~n8212;
  assign n8213 = ~INSTQUEUE_REG_2__7__SCAN_IN | ~n8169;
  assign n8218 = ~n8214 | ~n8213;
  assign n8216 = ~INSTQUEUE_REG_5__7__SCAN_IN | ~n6293;
  assign n8215 = ~INSTQUEUE_REG_15__7__SCAN_IN | ~n6287;
  assign n8217 = ~n8216 | ~n8215;
  assign n8228 = ~n8218 & ~n8217;
  assign n8221 = ~INSTQUEUE_REG_10__7__SCAN_IN | ~n8182;
  assign n8220 = ~INSTQUEUE_REG_13__7__SCAN_IN | ~n8219;
  assign n8226 = ~n8221 | ~n8220;
  assign n8224 = ~INSTQUEUE_REG_4__7__SCAN_IN | ~n8178;
  assign n8223 = ~INSTQUEUE_REG_1__7__SCAN_IN | ~n8222;
  assign n8225 = ~n8224 | ~n8223;
  assign n8227 = ~n8226 & ~n8225;
  assign n8250 = ~n8228 | ~n8227;
  assign n8232 = ~INSTQUEUE_REG_14__7__SCAN_IN | ~n8119;
  assign n8231 = ~INSTQUEUE_REG_9__7__SCAN_IN | ~n6291;
  assign n8237 = ~n8232 | ~n8231;
  assign n8235 = ~INSTQUEUE_REG_8__7__SCAN_IN | ~n8187;
  assign n8234 = ~INSTQUEUE_REG_12__7__SCAN_IN | ~n6298;
  assign n8236 = ~n8235 | ~n8234;
  assign n8248 = ~n8237 & ~n8236;
  assign n8241 = ~INSTQUEUE_REG_0__7__SCAN_IN | ~n8238;
  assign n8240 = ~INSTQUEUE_REG_3__7__SCAN_IN | ~n8239;
  assign n8246 = ~n8241 | ~n8240;
  assign n8244 = ~INSTQUEUE_REG_6__7__SCAN_IN | ~n8242;
  assign n8243 = ~INSTQUEUE_REG_11__7__SCAN_IN | ~n6302;
  assign n8245 = ~n8244 | ~n8243;
  assign n8247 = ~n8246 & ~n8245;
  assign n8249 = ~n8248 | ~n8247;
  assign n8259 = ~n8250 & ~n8249;
  assign n8262 = ~n8252 | ~n8251;
  assign n8254 = ~n8253 | ~n8262;
  assign n8255 = ~n8259 & ~n8254;
  assign n8258 = ~n8256 & ~n8255;
  assign n8257 = ~n7751 | ~EAX_REG_30__SCAN_IN;
  assign n8264 = ~n8258 | ~n8257;
  assign n8261 = ~n8260 | ~n8259;
  assign n8263 = ~n8262 & ~n8261;
  assign n8268 = ~n8264 & ~n8263;
  assign n8265 = ~PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n8656 = PHYADDRPOINTER_REG_30__SCAN_IN ^ ~n8555;
  assign n8267 = ~n8656 & ~n9025;
  assign n8548 = ~n8268 & ~n8267;
  assign n8677 = ~n6296 | ~n8445;
  assign n8666 = ~n8386 & ~STATE_REG_0__SCAN_IN;
  assign n8389 = ~n8388 | ~n8387;
  assign n8391 = ~n8390 & ~n8389;
  assign n8678 = ~n8392 & ~n8391;
  assign n8397 = ~n8666 & ~n9757;
  assign n8639 = ~READY_N & ~n8397;
  assign n8422 = ~EBX_REG_31__SCAN_IN | ~n10181;
  assign n8421 = ~INSTADDRPOINTER_REG_31__SCAN_IN | ~n6547;
  assign n8428 = ~n8422 | ~n8421;
  assign n8427 = ~n8426 | ~n8425;
  assign n11178 = n8428 ^ n8427;
  assign n9290 = ~STATE2_REG_0__SCAN_IN & ~n11908;
  assign n8547 = ~n8546;
  assign n8549 = n8621 | n6373;
  assign n8552 = ~PHYADDRPOINTER_REG_31__SCAN_IN | ~n8550;
  assign n8551 = ~EAX_REG_31__SCAN_IN | ~n7751;
  assign n8553 = ~n8552 | ~n8551;
  assign n8556 = ~n8555 | ~PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n9020 = ~PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n8570 = ~n8678;
  assign n8629 = ~n9476 | ~n8668;
  assign n11911 = ~n9290 | ~n8628;
  assign n8630 = ~n9270 | ~n8629;
  assign n9269 = ~n11899 | ~n8669;
  assign n9271 = ~n11899 | ~n8668;
  assign n9276 = ~n9269 | ~n9271;
  assign n9730 = ~n11908 | ~n10732;
  assign n8631 = ~n9734 & ~n9730;
  assign n8805 = ~STATE2_REG_3__SCAN_IN | ~n8631;
  assign n8632 = ~n11647 | ~n8805;
  assign n8655 = ~n11908 & ~n10888;
  assign n8634 = ~n8655;
  assign n9209 = ~REIP_REG_26__SCAN_IN;
  assign n12158 = ~REIP_REG_25__SCAN_IN;
  assign n8636 = ~n9209 & ~n12158;
  assign n12316 = ~REIP_REG_27__SCAN_IN | ~n8636;
  assign n8959 = ~REIP_REG_21__SCAN_IN | ~REIP_REG_20__SCAN_IN;
  assign n11827 = ~REIP_REG_14__SCAN_IN;
  assign n11160 = ~REIP_REG_13__SCAN_IN;
  assign n8872 = ~n11827 & ~n11160;
  assign n11646 = ~REIP_REG_10__SCAN_IN;
  assign n11624 = ~REIP_REG_11__SCAN_IN;
  assign n11193 = ~n11646 & ~n11624;
  assign n8871 = ~n11193 | ~REIP_REG_12__SCAN_IN;
  assign n10881 = ~REIP_REG_3__SCAN_IN | ~REIP_REG_2__SCAN_IN;
  assign n10870 = ~REIP_REG_4__SCAN_IN;
  assign n8869 = ~n10881 & ~n10870;
  assign n9459 = ~REIP_REG_1__SCAN_IN;
  assign n11498 = ~n10888 & ~n9459;
  assign n10869 = ~n8869 | ~n11498;
  assign n11856 = ~REIP_REG_5__SCAN_IN;
  assign n8637 = ~n10869 & ~n11856;
  assign n11632 = ~REIP_REG_6__SCAN_IN | ~n8637;
  assign n11633 = ~REIP_REG_7__SCAN_IN;
  assign n11842 = ~n11632 & ~n11633;
  assign n9169 = ~REIP_REG_9__SCAN_IN;
  assign n11846 = ~REIP_REG_8__SCAN_IN;
  assign n8870 = ~n9169 & ~n11846;
  assign n11122 = ~n11842 | ~n8870;
  assign n11151 = ~n8871 & ~n11122;
  assign n11829 = ~n8872 | ~n11151;
  assign n11247 = ~REIP_REG_15__SCAN_IN;
  assign n11246 = ~n11829 & ~n11247;
  assign n11923 = ~n11246 | ~REIP_REG_16__SCAN_IN;
  assign n8638 = ~REIP_REG_17__SCAN_IN | ~REIP_REG_18__SCAN_IN;
  assign n11943 = ~n11923 & ~n8638;
  assign n8855 = ~n11943 | ~REIP_REG_19__SCAN_IN;
  assign n8914 = ~n8959 & ~n8855;
  assign n8924 = ~REIP_REG_22__SCAN_IN | ~n8914;
  assign n9195 = ~REIP_REG_23__SCAN_IN;
  assign n12157 = ~REIP_REG_24__SCAN_IN | ~n12130;
  assign n12253 = ~n12316 & ~n12157;
  assign n8643 = ~REIP_REG_28__SCAN_IN | ~n12253;
  assign n8650 = ~n9821 | ~n10875;
  assign n8647 = ~n8639 | ~n11362;
  assign n12437 = ~n8643 | ~n12156;
  assign n9016 = ~REIP_REG_30__SCAN_IN | ~REIP_REG_29__SCAN_IN;
  assign n8640 = ~n12129 | ~n9016;
  assign n9023 = ~n12437 | ~n8640;
  assign n8788 = ~STATEBS16_REG_SCAN_IN & ~READY_N;
  assign n8648 = ~EBX_REG_31__SCAN_IN | ~n9757;
  assign n8641 = n8788 | n8648;
  assign n12031 = ~n8650 & ~n8641;
  assign n11725 = ~STATE2_REG_3__SCAN_IN;
  assign n12427 = ~n8643 & ~n12150;
  assign n8649 = ~n8648 | ~n8647;
  assign n8651 = n8650 | n8649;
  assign n12434 = ~n8651;
  assign n9017 = ~REIP_REG_31__SCAN_IN & ~n9016;
  assign n9019 = ~n9017 | ~n12427;
  assign n9018 = ~n12434 | ~EBX_REG_31__SCAN_IN;
  assign n9022 = ~n9019 | ~n9018;
  assign n9021 = ~n9020 & ~n12256;
  assign keyinput_0 = 1'b0;
  assign keyinput_1 = 1'b1;
  assign keyinput_2 = 1'b0;
  assign keyinput_3 = 1'b0;
  assign keyinput_4 = 1'b1;
  assign keyinput_5 = 1'b0;
  assign keyinput_6 = 1'b1;
  assign keyinput_7 = 1'b0;
  assign keyinput_8 = 1'b1;
  assign keyinput_9 = 1'b1;
  assign keyinput_10 = 1'b0;
  assign keyinput_11 = 1'b1;
  assign keyinput_12 = 1'b0;
  assign keyinput_13 = 1'b1;
  assign keyinput_14 = 1'b0;
  assign keyinput_15 = 1'b1;
  assign keyinput_16 = 1'b0;
  assign keyinput_17 = 1'b0;
  assign keyinput_18 = 1'b1;
  assign keyinput_19 = 1'b0;
  assign keyinput_20 = 1'b0;
  assign keyinput_21 = 1'b1;
  assign keyinput_22 = 1'b0;
  assign keyinput_23 = 1'b1;
  assign keyinput_24 = 1'b1;
  assign keyinput_25 = 1'b1;
  assign keyinput_26 = 1'b1;
  assign keyinput_27 = 1'b0;
  assign keyinput_28 = 1'b0;
  assign keyinput_29 = 1'b1;
  assign keyinput_30 = 1'b1;
  assign keyinput_31 = 1'b0;
  assign keyinput_32 = 1'b1;
  assign keyinput_33 = 1'b0;
  assign keyinput_34 = 1'b0;
  assign keyinput_35 = 1'b0;
  assign keyinput_36 = 1'b1;
  assign keyinput_37 = 1'b0;
  assign keyinput_38 = 1'b0;
  assign keyinput_39 = 1'b0;
  assign keyinput_40 = 1'b0;
  assign keyinput_41 = 1'b0;
  assign keyinput_42 = 1'b0;
  assign keyinput_43 = 1'b1;
  assign keyinput_44 = 1'b1;
  assign keyinput_45 = 1'b1;
  assign keyinput_46 = 1'b0;
  assign keyinput_47 = 1'b1;
  assign keyinput_48 = 1'b0;
  assign keyinput_49 = 1'b1;
  assign keyinput_50 = 1'b0;
  assign keyinput_51 = 1'b0;
  assign keyinput_52 = 1'b0;
  assign keyinput_53 = 1'b1;
  assign keyinput_54 = 1'b0;
  assign keyinput_55 = 1'b1;
  assign keyinput_56 = 1'b1;
  assign keyinput_57 = 1'b1;
  assign keyinput_58 = 1'b0;
  assign keyinput_59 = 1'b1;
  assign keyinput_60 = 1'b0;
  assign keyinput_61 = 1'b0;
  assign keyinput_62 = 1'b0;
  assign keyinput_63 = 1'b0;
  assign keyinput_64 = 1'b0;
  assign keyinput_65 = 1'b1;
  assign keyinput_66 = 1'b0;
  assign keyinput_67 = 1'b0;
  assign keyinput_68 = 1'b1;
  assign keyinput_69 = 1'b1;
  assign keyinput_70 = 1'b0;
  assign keyinput_71 = 1'b1;
  assign keyinput_72 = 1'b0;
  assign keyinput_73 = 1'b0;
  assign keyinput_74 = 1'b1;
  assign keyinput_75 = 1'b0;
  assign keyinput_76 = 1'b0;
  assign keyinput_77 = 1'b1;
  assign keyinput_78 = 1'b1;
  assign keyinput_79 = 1'b1;
  assign keyinput_80 = 1'b0;
  assign keyinput_81 = 1'b0;
  assign keyinput_82 = 1'b1;
  assign keyinput_83 = 1'b0;
  assign keyinput_84 = 1'b0;
  assign keyinput_85 = 1'b0;
  assign keyinput_86 = 1'b1;
  assign keyinput_87 = 1'b1;
  assign keyinput_88 = 1'b1;
  assign keyinput_89 = 1'b0;
  assign keyinput_90 = 1'b1;
  assign keyinput_91 = 1'b0;
  assign keyinput_92 = 1'b0;
  assign keyinput_93 = 1'b0;
  assign keyinput_94 = 1'b1;
  assign keyinput_95 = 1'b1;
  assign keyinput_96 = 1'b1;
  assign keyinput_97 = 1'b0;
  assign keyinput_98 = 1'b0;
  assign keyinput_99 = 1'b0;
  assign keyinput_100 = 1'b0;
  assign keyinput_101 = 1'b1;
  assign keyinput_102 = 1'b0;
  assign keyinput_103 = 1'b0;
  assign keyinput_104 = 1'b0;
  assign keyinput_105 = 1'b1;
  assign keyinput_106 = 1'b1;
  assign keyinput_107 = 1'b0;
  assign keyinput_108 = 1'b1;
  assign keyinput_109 = 1'b0;
  assign keyinput_110 = 1'b1;
  assign keyinput_111 = 1'b0;
  assign keyinput_112 = 1'b0;
  assign keyinput_113 = 1'b1;
  assign keyinput_114 = 1'b0;
  assign keyinput_115 = 1'b0;
  assign keyinput_116 = 1'b0;
  assign keyinput_117 = 1'b0;
  assign keyinput_118 = 1'b1;
  assign keyinput_119 = 1'b0;
  assign keyinput_120 = 1'b0;
  assign keyinput_121 = 1'b0;
  assign keyinput_122 = 1'b0;
  assign keyinput_123 = 1'b0;
  assign keyinput_124 = 1'b0;
  assign keyinput_125 = 1'b0;
  assign keyinput_126 = 1'b1;
  assign keyinput_127 = 1'b0;
  assign keyinput_128 = 1'b0;
  assign keyinput_129 = 1'b1;
  assign keyinput_130 = 1'b0;
  assign keyinput_131 = 1'b1;
  assign keyinput_132 = 1'b1;
  assign keyinput_133 = 1'b0;
  assign keyinput_134 = 1'b1;
  assign keyinput_135 = 1'b1;
  assign keyinput_136 = 1'b0;
  assign keyinput_137 = 1'b0;
  assign keyinput_138 = 1'b1;
  assign keyinput_139 = 1'b0;
  assign keyinput_140 = 1'b1;
  assign keyinput_141 = 1'b0;
  assign keyinput_142 = 1'b0;
  assign keyinput_143 = 1'b0;
  assign keyinput_144 = 1'b0;
  assign keyinput_145 = 1'b1;
  assign keyinput_146 = 1'b0;
  assign keyinput_147 = 1'b1;
  assign keyinput_148 = 1'b0;
  assign keyinput_149 = 1'b0;
  assign keyinput_150 = 1'b1;
  assign keyinput_151 = 1'b0;
  assign keyinput_152 = 1'b1;
  assign keyinput_153 = 1'b1;
  assign keyinput_154 = 1'b1;
  assign keyinput_155 = 1'b0;
  assign keyinput_156 = 1'b0;
  assign keyinput_157 = 1'b0;
  assign keyinput_158 = 1'b1;
  assign keyinput_159 = 1'b1;
  assign input_0 = keyinput_0 ^ READY_N;
  assign input_1 = keyinput_1 ^ STATEBS16_REG_SCAN_IN;
  assign AND_1 = input_0 & input_1;
  assign input_2 = keyinput_2 ^ REIP_REG_31__SCAN_IN;
  assign OR_2 = input_2 | AND_1;
  assign input_3 = keyinput_3 ^ REIP_REG_30__SCAN_IN;
  assign AND_3 = input_3 & OR_2;
  assign input_4 = keyinput_4 ^ REIP_REG_29__SCAN_IN;
  assign OR_4 = input_4 | AND_3;
  assign input_5 = keyinput_5 ^ REIP_REG_28__SCAN_IN;
  assign OR_5 = input_5 | OR_4;
  assign input_6 = keyinput_6 ^ REIP_REG_27__SCAN_IN;
  assign AND_6 = input_6 & OR_5;
  assign input_7 = keyinput_7 ^ REIP_REG_26__SCAN_IN;
  assign AND_7 = input_7 & AND_6;
  assign input_8 = keyinput_8 ^ REIP_REG_25__SCAN_IN;
  assign OR_8 = input_8 | AND_7;
  assign input_9 = keyinput_9 ^ REIP_REG_24__SCAN_IN;
  assign OR_9 = input_9 | OR_8;
  assign input_10 = keyinput_10 ^ REIP_REG_23__SCAN_IN;
  assign OR_10 = input_10 | OR_9;
  assign input_11 = keyinput_11 ^ REIP_REG_22__SCAN_IN;
  assign AND_11 = input_11 & OR_10;
  assign input_12 = keyinput_12 ^ REIP_REG_21__SCAN_IN;
  assign OR_12 = input_12 | AND_11;
  assign input_13 = keyinput_13 ^ REIP_REG_20__SCAN_IN;
  assign AND_13 = input_13 & OR_12;
  assign input_14 = keyinput_14 ^ REIP_REG_19__SCAN_IN;
  assign AND_14 = input_14 & AND_13;
  assign input_15 = keyinput_15 ^ REIP_REG_18__SCAN_IN;
  assign OR_15 = input_15 | AND_14;
  assign input_16 = keyinput_16 ^ REIP_REG_17__SCAN_IN;
  assign AND_16 = input_16 & OR_15;
  assign input_17 = keyinput_17 ^ REIP_REG_16__SCAN_IN;
  assign OR_17 = input_17 | AND_16;
  assign input_18 = keyinput_18 ^ STATE_REG_2__SCAN_IN;
  assign OR_18 = input_18 | OR_17;
  assign input_19 = keyinput_19 ^ STATE_REG_1__SCAN_IN;
  assign OR_19 = input_19 | OR_18;
  assign input_20 = keyinput_20 ^ STATE_REG_0__SCAN_IN;
  assign OR_20 = input_20 | OR_19;
  assign input_21 = keyinput_21 ^ STATE2_REG_3__SCAN_IN;
  assign AND_21 = input_21 & OR_20;
  assign input_22 = keyinput_22 ^ STATE2_REG_2__SCAN_IN;
  assign OR_22 = input_22 | AND_21;
  assign input_23 = keyinput_23 ^ STATE2_REG_1__SCAN_IN;
  assign AND_23 = input_23 & OR_22;
  assign input_24 = keyinput_24 ^ STATE2_REG_0__SCAN_IN;
  assign AND_24 = input_24 & AND_23;
  assign input_25 = keyinput_25 ^ INSTQUEUE_REG_15__7__SCAN_IN;
  assign OR_25 = input_25 | AND_24;
  assign input_26 = keyinput_26 ^ INSTQUEUE_REG_15__6__SCAN_IN;
  assign OR_26 = input_26 | OR_25;
  assign input_27 = keyinput_27 ^ INSTQUEUE_REG_15__5__SCAN_IN;
  assign OR_27 = input_27 | OR_26;
  assign input_28 = keyinput_28 ^ INSTQUEUE_REG_15__4__SCAN_IN;
  assign OR_28 = input_28 | OR_27;
  assign input_29 = keyinput_29 ^ INSTQUEUE_REG_15__3__SCAN_IN;
  assign OR_29 = input_29 | OR_28;
  assign input_30 = keyinput_30 ^ INSTQUEUE_REG_15__2__SCAN_IN;
  assign AND_30 = input_30 & OR_29;
  assign input_31 = keyinput_31 ^ INSTQUEUE_REG_15__1__SCAN_IN;
  assign OR_31 = input_31 | AND_30;
  assign input_32 = keyinput_32 ^ INSTQUEUE_REG_15__0__SCAN_IN;
  assign OR_32 = input_32 | OR_31;
  assign input_33 = keyinput_33 ^ INSTQUEUE_REG_14__7__SCAN_IN;
  assign OR_33 = input_33 | OR_32;
  assign input_34 = keyinput_34 ^ INSTQUEUE_REG_14__6__SCAN_IN;
  assign OR_34 = input_34 | OR_33;
  assign input_35 = keyinput_35 ^ INSTQUEUE_REG_14__5__SCAN_IN;
  assign OR_35 = input_35 | OR_34;
  assign input_36 = keyinput_36 ^ INSTQUEUE_REG_14__4__SCAN_IN;
  assign AND_36 = input_36 & OR_35;
  assign input_37 = keyinput_37 ^ INSTQUEUE_REG_14__3__SCAN_IN;
  assign AND_37 = input_37 & AND_36;
  assign input_38 = keyinput_38 ^ INSTQUEUE_REG_14__2__SCAN_IN;
  assign OR_38 = input_38 | AND_37;
  assign input_39 = keyinput_39 ^ INSTQUEUE_REG_14__1__SCAN_IN;
  assign AND_39 = input_39 & OR_38;
  assign input_40 = keyinput_40 ^ INSTQUEUE_REG_14__0__SCAN_IN;
  assign OR_40 = input_40 | AND_39;
  assign input_41 = keyinput_41 ^ INSTQUEUE_REG_13__7__SCAN_IN;
  assign AND_41 = input_41 & OR_40;
  assign input_42 = keyinput_42 ^ INSTQUEUE_REG_13__6__SCAN_IN;
  assign OR_42 = input_42 | AND_41;
  assign input_43 = keyinput_43 ^ INSTQUEUE_REG_13__5__SCAN_IN;
  assign OR_43 = input_43 | OR_42;
  assign input_44 = keyinput_44 ^ INSTQUEUE_REG_13__4__SCAN_IN;
  assign OR_44 = input_44 | OR_43;
  assign input_45 = keyinput_45 ^ INSTQUEUE_REG_13__3__SCAN_IN;
  assign AND_45 = input_45 & OR_44;
  assign input_46 = keyinput_46 ^ INSTQUEUE_REG_13__2__SCAN_IN;
  assign OR_46 = input_46 | AND_45;
  assign input_47 = keyinput_47 ^ INSTQUEUE_REG_13__1__SCAN_IN;
  assign OR_47 = input_47 | OR_46;
  assign input_48 = keyinput_48 ^ INSTQUEUE_REG_13__0__SCAN_IN;
  assign OR_48 = input_48 | OR_47;
  assign input_49 = keyinput_49 ^ INSTQUEUE_REG_12__7__SCAN_IN;
  assign OR_49 = input_49 | OR_48;
  assign input_50 = keyinput_50 ^ INSTQUEUE_REG_12__6__SCAN_IN;
  assign AND_50 = input_50 & OR_49;
  assign input_51 = keyinput_51 ^ INSTQUEUE_REG_12__5__SCAN_IN;
  assign OR_51 = input_51 | AND_50;
  assign input_52 = keyinput_52 ^ INSTQUEUE_REG_12__4__SCAN_IN;
  assign OR_52 = input_52 | OR_51;
  assign input_53 = keyinput_53 ^ INSTQUEUE_REG_12__3__SCAN_IN;
  assign AND_53 = input_53 & OR_52;
  assign input_54 = keyinput_54 ^ INSTQUEUE_REG_12__2__SCAN_IN;
  assign OR_54 = input_54 | AND_53;
  assign input_55 = keyinput_55 ^ INSTQUEUE_REG_12__1__SCAN_IN;
  assign OR_55 = input_55 | OR_54;
  assign input_56 = keyinput_56 ^ INSTQUEUE_REG_12__0__SCAN_IN;
  assign OR_56 = input_56 | OR_55;
  assign input_57 = keyinput_57 ^ INSTQUEUE_REG_11__7__SCAN_IN;
  assign AND_57 = input_57 & OR_56;
  assign input_58 = keyinput_58 ^ INSTQUEUE_REG_11__6__SCAN_IN;
  assign OR_58 = input_58 | AND_57;
  assign input_59 = keyinput_59 ^ INSTQUEUE_REG_11__5__SCAN_IN;
  assign AND_59 = input_59 & OR_58;
  assign input_60 = keyinput_60 ^ INSTQUEUE_REG_11__4__SCAN_IN;
  assign AND_60 = input_60 & AND_59;
  assign input_61 = keyinput_61 ^ INSTQUEUE_REG_11__3__SCAN_IN;
  assign AND_61 = input_61 & AND_60;
  assign input_62 = keyinput_62 ^ INSTQUEUE_REG_11__2__SCAN_IN;
  assign AND_62 = input_62 & AND_61;
  assign input_63 = keyinput_63 ^ INSTQUEUE_REG_11__1__SCAN_IN;
  assign OR_63 = input_63 | AND_62;
  assign input_64 = keyinput_64 ^ INSTQUEUE_REG_11__0__SCAN_IN;
  assign AND_64 = input_64 & OR_63;
  assign input_65 = keyinput_65 ^ INSTQUEUE_REG_10__7__SCAN_IN;
  assign OR_65 = input_65 | AND_64;
  assign input_66 = keyinput_66 ^ INSTQUEUE_REG_10__6__SCAN_IN;
  assign OR_66 = input_66 | OR_65;
  assign input_67 = keyinput_67 ^ INSTQUEUE_REG_10__5__SCAN_IN;
  assign OR_67 = input_67 | OR_66;
  assign input_68 = keyinput_68 ^ INSTQUEUE_REG_10__4__SCAN_IN;
  assign AND_68 = input_68 & OR_67;
  assign input_69 = keyinput_69 ^ INSTQUEUE_REG_10__3__SCAN_IN;
  assign AND_69 = input_69 & AND_68;
  assign input_70 = keyinput_70 ^ INSTQUEUE_REG_10__2__SCAN_IN;
  assign AND_70 = input_70 & AND_69;
  assign input_71 = keyinput_71 ^ INSTQUEUE_REG_10__1__SCAN_IN;
  assign AND_71 = input_71 & AND_70;
  assign input_72 = keyinput_72 ^ INSTQUEUE_REG_10__0__SCAN_IN;
  assign OR_72 = input_72 | AND_71;
  assign input_73 = keyinput_73 ^ INSTQUEUE_REG_9__7__SCAN_IN;
  assign OR_73 = input_73 | OR_72;
  assign input_74 = keyinput_74 ^ INSTQUEUE_REG_9__6__SCAN_IN;
  assign OR_74 = input_74 | OR_73;
  assign input_75 = keyinput_75 ^ INSTQUEUE_REG_9__5__SCAN_IN;
  assign AND_75 = input_75 & OR_74;
  assign input_76 = keyinput_76 ^ INSTQUEUE_REG_9__4__SCAN_IN;
  assign OR_76 = input_76 | AND_75;
  assign input_77 = keyinput_77 ^ INSTQUEUE_REG_9__3__SCAN_IN;
  assign OR_77 = input_77 | OR_76;
  assign input_78 = keyinput_78 ^ INSTQUEUE_REG_9__2__SCAN_IN;
  assign OR_78 = input_78 | OR_77;
  assign input_79 = keyinput_79 ^ INSTQUEUE_REG_9__1__SCAN_IN;
  assign OR_79 = input_79 | OR_78;
  assign input_80 = keyinput_80 ^ READY_N;
  assign input_81 = keyinput_81 ^ STATEBS16_REG_SCAN_IN;
  assign AND_81 = input_80 & input_81;
  assign input_82 = keyinput_82 ^ REIP_REG_31__SCAN_IN;
  assign OR_82 = input_82 | AND_81;
  assign input_83 = keyinput_83 ^ REIP_REG_30__SCAN_IN;
  assign AND_83 = input_83 & OR_82;
  assign input_84 = keyinput_84 ^ REIP_REG_29__SCAN_IN;
  assign OR_84 = input_84 | AND_83;
  assign input_85 = keyinput_85 ^ REIP_REG_28__SCAN_IN;
  assign OR_85 = input_85 | OR_84;
  assign input_86 = keyinput_86 ^ REIP_REG_27__SCAN_IN;
  assign AND_86 = input_86 & OR_85;
  assign input_87 = keyinput_87 ^ REIP_REG_26__SCAN_IN;
  assign AND_87 = input_87 & AND_86;
  assign input_88 = keyinput_88 ^ REIP_REG_25__SCAN_IN;
  assign OR_88 = input_88 | AND_87;
  assign input_89 = keyinput_89 ^ REIP_REG_24__SCAN_IN;
  assign OR_89 = input_89 | OR_88;
  assign input_90 = keyinput_90 ^ REIP_REG_23__SCAN_IN;
  assign OR_90 = input_90 | OR_89;
  assign input_91 = keyinput_91 ^ REIP_REG_22__SCAN_IN;
  assign AND_91 = input_91 & OR_90;
  assign input_92 = keyinput_92 ^ REIP_REG_21__SCAN_IN;
  assign OR_92 = input_92 | AND_91;
  assign input_93 = keyinput_93 ^ REIP_REG_20__SCAN_IN;
  assign AND_93 = input_93 & OR_92;
  assign input_94 = keyinput_94 ^ REIP_REG_19__SCAN_IN;
  assign AND_94 = input_94 & AND_93;
  assign input_95 = keyinput_95 ^ REIP_REG_18__SCAN_IN;
  assign OR_95 = input_95 | AND_94;
  assign input_96 = keyinput_96 ^ REIP_REG_17__SCAN_IN;
  assign AND_96 = input_96 & OR_95;
  assign input_97 = keyinput_97 ^ REIP_REG_16__SCAN_IN;
  assign OR_97 = input_97 | AND_96;
  assign input_98 = keyinput_98 ^ STATE_REG_2__SCAN_IN;
  assign OR_98 = input_98 | OR_97;
  assign input_99 = keyinput_99 ^ STATE_REG_1__SCAN_IN;
  assign OR_99 = input_99 | OR_98;
  assign input_100 = keyinput_100 ^ STATE_REG_0__SCAN_IN;
  assign OR_100 = input_100 | OR_99;
  assign input_101 = keyinput_101 ^ STATE2_REG_3__SCAN_IN;
  assign AND_101 = input_101 & OR_100;
  assign input_102 = keyinput_102 ^ STATE2_REG_2__SCAN_IN;
  assign OR_102 = input_102 | AND_101;
  assign input_103 = keyinput_103 ^ STATE2_REG_1__SCAN_IN;
  assign AND_103 = input_103 & OR_102;
  assign input_104 = keyinput_104 ^ STATE2_REG_0__SCAN_IN;
  assign AND_104 = input_104 & AND_103;
  assign input_105 = keyinput_105 ^ INSTQUEUE_REG_15__7__SCAN_IN;
  assign OR_105 = input_105 | AND_104;
  assign input_106 = keyinput_106 ^ INSTQUEUE_REG_15__6__SCAN_IN;
  assign OR_106 = input_106 | OR_105;
  assign input_107 = keyinput_107 ^ INSTQUEUE_REG_15__5__SCAN_IN;
  assign OR_107 = input_107 | OR_106;
  assign input_108 = keyinput_108 ^ INSTQUEUE_REG_15__4__SCAN_IN;
  assign OR_108 = input_108 | OR_107;
  assign input_109 = keyinput_109 ^ INSTQUEUE_REG_15__3__SCAN_IN;
  assign OR_109 = input_109 | OR_108;
  assign input_110 = keyinput_110 ^ INSTQUEUE_REG_15__2__SCAN_IN;
  assign AND_110 = input_110 & OR_109;
  assign input_111 = keyinput_111 ^ INSTQUEUE_REG_15__1__SCAN_IN;
  assign OR_111 = input_111 | AND_110;
  assign input_112 = keyinput_112 ^ INSTQUEUE_REG_15__0__SCAN_IN;
  assign OR_112 = input_112 | OR_111;
  assign input_113 = keyinput_113 ^ INSTQUEUE_REG_14__7__SCAN_IN;
  assign OR_113 = input_113 | OR_112;
  assign input_114 = keyinput_114 ^ INSTQUEUE_REG_14__6__SCAN_IN;
  assign OR_114 = input_114 | OR_113;
  assign input_115 = keyinput_115 ^ INSTQUEUE_REG_14__5__SCAN_IN;
  assign OR_115 = input_115 | OR_114;
  assign input_116 = keyinput_116 ^ INSTQUEUE_REG_14__4__SCAN_IN;
  assign AND_116 = input_116 & OR_115;
  assign input_117 = keyinput_117 ^ INSTQUEUE_REG_14__3__SCAN_IN;
  assign AND_117 = input_117 & AND_116;
  assign input_118 = keyinput_118 ^ INSTQUEUE_REG_14__2__SCAN_IN;
  assign OR_118 = input_118 | AND_117;
  assign input_119 = keyinput_119 ^ INSTQUEUE_REG_14__1__SCAN_IN;
  assign AND_119 = input_119 & OR_118;
  assign input_120 = keyinput_120 ^ INSTQUEUE_REG_14__0__SCAN_IN;
  assign OR_120 = input_120 | AND_119;
  assign input_121 = keyinput_121 ^ INSTQUEUE_REG_13__7__SCAN_IN;
  assign AND_121 = input_121 & OR_120;
  assign input_122 = keyinput_122 ^ INSTQUEUE_REG_13__6__SCAN_IN;
  assign OR_122 = input_122 | AND_121;
  assign input_123 = keyinput_123 ^ INSTQUEUE_REG_13__5__SCAN_IN;
  assign OR_123 = input_123 | OR_122;
  assign input_124 = keyinput_124 ^ INSTQUEUE_REG_13__4__SCAN_IN;
  assign OR_124 = input_124 | OR_123;
  assign input_125 = keyinput_125 ^ INSTQUEUE_REG_13__3__SCAN_IN;
  assign AND_125 = input_125 & OR_124;
  assign input_126 = keyinput_126 ^ INSTQUEUE_REG_13__2__SCAN_IN;
  assign OR_126 = input_126 | AND_125;
  assign input_127 = keyinput_127 ^ INSTQUEUE_REG_13__1__SCAN_IN;
  assign OR_127 = input_127 | OR_126;
  assign input_128 = keyinput_128 ^ INSTQUEUE_REG_13__0__SCAN_IN;
  assign OR_128 = input_128 | OR_127;
  assign input_129 = keyinput_129 ^ INSTQUEUE_REG_12__7__SCAN_IN;
  assign OR_129 = input_129 | OR_128;
  assign input_130 = keyinput_130 ^ INSTQUEUE_REG_12__6__SCAN_IN;
  assign AND_130 = input_130 & OR_129;
  assign input_131 = keyinput_131 ^ INSTQUEUE_REG_12__5__SCAN_IN;
  assign OR_131 = input_131 | AND_130;
  assign input_132 = keyinput_132 ^ INSTQUEUE_REG_12__4__SCAN_IN;
  assign OR_132 = input_132 | OR_131;
  assign input_133 = keyinput_133 ^ INSTQUEUE_REG_12__3__SCAN_IN;
  assign AND_133 = input_133 & OR_132;
  assign input_134 = keyinput_134 ^ INSTQUEUE_REG_12__2__SCAN_IN;
  assign OR_134 = input_134 | AND_133;
  assign input_135 = keyinput_135 ^ INSTQUEUE_REG_12__1__SCAN_IN;
  assign OR_135 = input_135 | OR_134;
  assign input_136 = keyinput_136 ^ INSTQUEUE_REG_12__0__SCAN_IN;
  assign OR_136 = input_136 | OR_135;
  assign input_137 = keyinput_137 ^ INSTQUEUE_REG_11__7__SCAN_IN;
  assign AND_137 = input_137 & OR_136;
  assign input_138 = keyinput_138 ^ INSTQUEUE_REG_11__6__SCAN_IN;
  assign OR_138 = input_138 | AND_137;
  assign input_139 = keyinput_139 ^ INSTQUEUE_REG_11__5__SCAN_IN;
  assign AND_139 = input_139 & OR_138;
  assign input_140 = keyinput_140 ^ INSTQUEUE_REG_11__4__SCAN_IN;
  assign AND_140 = input_140 & AND_139;
  assign input_141 = keyinput_141 ^ INSTQUEUE_REG_11__3__SCAN_IN;
  assign AND_141 = input_141 & AND_140;
  assign input_142 = keyinput_142 ^ INSTQUEUE_REG_11__2__SCAN_IN;
  assign AND_142 = input_142 & AND_141;
  assign input_143 = keyinput_143 ^ INSTQUEUE_REG_11__1__SCAN_IN;
  assign OR_143 = input_143 | AND_142;
  assign input_144 = keyinput_144 ^ INSTQUEUE_REG_11__0__SCAN_IN;
  assign AND_144 = input_144 & OR_143;
  assign input_145 = keyinput_145 ^ INSTQUEUE_REG_10__7__SCAN_IN;
  assign OR_145 = input_145 | AND_144;
  assign input_146 = keyinput_146 ^ INSTQUEUE_REG_10__6__SCAN_IN;
  assign OR_146 = input_146 | OR_145;
  assign input_147 = keyinput_147 ^ INSTQUEUE_REG_10__5__SCAN_IN;
  assign OR_147 = input_147 | OR_146;
  assign input_148 = keyinput_148 ^ INSTQUEUE_REG_10__4__SCAN_IN;
  assign AND_148 = input_148 & OR_147;
  assign input_149 = keyinput_149 ^ INSTQUEUE_REG_10__3__SCAN_IN;
  assign AND_149 = input_149 & AND_148;
  assign input_150 = keyinput_150 ^ INSTQUEUE_REG_10__2__SCAN_IN;
  assign AND_150 = input_150 & AND_149;
  assign input_151 = keyinput_151 ^ INSTQUEUE_REG_10__1__SCAN_IN;
  assign AND_151 = input_151 & AND_150;
  assign input_152 = keyinput_152 ^ INSTQUEUE_REG_10__0__SCAN_IN;
  assign OR_152 = input_152 | AND_151;
  assign input_153 = keyinput_153 ^ INSTQUEUE_REG_9__7__SCAN_IN;
  assign OR_153 = input_153 | OR_152;
  assign input_154 = keyinput_154 ^ INSTQUEUE_REG_9__6__SCAN_IN;
  assign OR_154 = input_154 | OR_153;
  assign input_155 = keyinput_155 ^ INSTQUEUE_REG_9__5__SCAN_IN;
  assign AND_155 = input_155 & OR_154;
  assign input_156 = keyinput_156 ^ INSTQUEUE_REG_9__4__SCAN_IN;
  assign OR_156 = input_156 | AND_155;
  assign input_157 = keyinput_157 ^ INSTQUEUE_REG_9__3__SCAN_IN;
  assign OR_157 = input_157 | OR_156;
  assign input_158 = keyinput_158 ^ INSTQUEUE_REG_9__2__SCAN_IN;
  assign OR_158 = input_158 | OR_157;
  assign input_159 = keyinput_159 ^ INSTQUEUE_REG_9__1__SCAN_IN;
  assign OR_159 = input_159 | OR_158;
  assign OR_159_INV = ~OR_159;
  assign CASOP = OR_79 & OR_159_INV;
  assign U2796 = U2796_Lock ^ CASOP;
endmodule


