// Benchmark "b15_C" written by ABC on Thu Mar  5 01:03:44 2020

module b15_C ( 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
    READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
    M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
    STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
    W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
    BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
    BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
    REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
    REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
    REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
    REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
    REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
    BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
    ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
    ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
    ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
    ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
    ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
    ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
    ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
    ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
    ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
    ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
    ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN,
    ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
    ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN,
    ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN,
    STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
    DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
    DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
    DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
    DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
    DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
    DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
    DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
    DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
    DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
    DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
    DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
    DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
    DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
    DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
    DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
    DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
    STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
    INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
    INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
    INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
    INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
    INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
    INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
    INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
    INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
    INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
    INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
    INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
    INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
    INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
    INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
    INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
    INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
    INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
    INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
    INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
    INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
    INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
    INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
    INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
    INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
    INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
    INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
    INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
    INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
    INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
    INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
    INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
    INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
    INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
    INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
    INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
    INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
    INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
    INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
    INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
    INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
    INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
    INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
    INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
    INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
    INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
    INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
    INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
    INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
    INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
    INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
    INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
    INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
    INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
    INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
    INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
    INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
    INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
    INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
    INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
    INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
    INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
    INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
    INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
    INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
    INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
    INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
    INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
    INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
    INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
    INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
    INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
    INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
    INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
    INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
    INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
    INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
    INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
    INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
    INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
    INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
    INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
    PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
    PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
    PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
    PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
    PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
    PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
    PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
    PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
    PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
    PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
    PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
    PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
    PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
    PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
    PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
    PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
    LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
    LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
    LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
    LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
    LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
    LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
    UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
    UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
    UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
    UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
    UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
    DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
    DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
    DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
    DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
    DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
    DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
    DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
    DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
    DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
    EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
    EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
    EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
    EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
    EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
    EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
    EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
    EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
    EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
    EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
    EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
    EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
    EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
    EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
    EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
    EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
    EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
    EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
    EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
    EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
    EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
    EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
    REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
    REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
    REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
    REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
    REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN,
    U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
    U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
    U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
    U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
    U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
    U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
    U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
    U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
    U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
    U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
    U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
    U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
    U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
    U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
    U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
    U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
    U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
    U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
    U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
    U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
    U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
    U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
    U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
    U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
    U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
    U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
    U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
    U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
    U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
    U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
    U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
    U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
    U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
    U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
    U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
    U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
    U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
    U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
    U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
    U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
    U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
    U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
    U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
    U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
    U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788  );
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N,
    HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
    CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
    REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
    FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
    BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
    BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
    REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
    REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
    REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
    REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
    REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
    BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
    ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
    ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
    ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
    ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
    ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
    ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
    ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
    ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
    ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
    ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
    ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN,
    ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
    ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN,
    ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN,
    STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
    DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
    DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
    DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
    DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
    DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
    DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
    DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
    DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
    DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
    DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
    DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
    DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
    DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
    DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
    DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
    DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
    STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
    INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
    INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
    INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
    INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
    INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
    INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
    INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
    INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
    INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
    INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
    INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
    INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
    INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
    INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
    INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
    INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
    INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
    INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
    INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
    INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
    INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
    INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
    INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
    INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
    INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
    INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
    INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
    INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
    INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
    INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
    INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
    INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
    INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
    INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
    INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
    INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
    INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
    INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
    INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
    INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
    INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
    INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
    INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
    INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
    INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
    INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
    INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
    INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
    INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
    INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
    INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
    INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
    INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
    INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
    INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
    INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
    INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
    INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
    INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
    INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
    INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
    INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
    INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
    INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
    INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
    INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
    INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
    INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
    INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
    INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
    INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
    INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
    INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
    INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
    INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
    INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
    INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
    INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
    INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
    INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
    INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
    PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
    PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
    PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
    PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
    PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
    PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
    PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
    PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
    PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
    PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
    PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
    PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
    PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
    PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
    PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
    PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
    LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
    LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
    LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
    LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
    LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
    LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
    UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
    UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
    UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
    UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
    UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
    DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
    DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
    DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
    DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
    DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
    DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
    DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
    DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
    DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
    EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
    EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
    EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
    EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
    EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
    EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
    EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
    EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
    EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
    EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
    EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
    EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
    EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
    EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
    EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
    EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
    EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
    EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
    EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
    EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
    EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
    EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
    REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
    REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
    REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
    REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
    REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
    U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
    U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
    U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
    U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
    U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
    U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
    U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
    U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
    U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
    U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
    U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
    U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
    U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
    U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
    U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
    U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
    U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
    U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
    U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
    U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
    U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
    U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
    U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
    U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
    U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
    U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
    U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
    U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
    U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
    U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
    U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
    U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
    U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
    U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
    U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
    U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
    U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
    U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
    U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
    U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
    U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
    U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
    U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
    U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire n13567, n13560, n13178, n13329, n10033, n9698, n8091, n8045, n10635,
    n10937, n8008, n10515, n9653, n7048, n7521, n7637, n7631, n8135, n8111,
    n10340, n8593, n8062, n8118, n8030, n8133, n12929, n10045, n13316,
    n13490, n13045, n8806, n13463, n13465, n13448, n13368, n13477, n13358,
    n13461, n13424, n9585, n13387, n13367, n9584, n13422, n13247, n13323,
    n13364, n13267, n13459, n13408, n13386, n13266, n13383, n13158, n13421,
    n13312, n13310, n9402, n13406, n13090, n13263, n9400, n13295, n13309,
    n13418, n13173, n13416, n9399, n13294, n13122, n13160, n13145, n9574,
    n13437, n13120, n13119, n13062, n9355, n13081, n13080, n13117, n13061,
    n13010, n9346, n13344, n13009, n9345, n13296, n13142, n13342, n9569,
    n13341, n9553, n13140, n13269, n12983, n9167, n13462, n12862, n13041,
    n13139, n13074, n13214, n12958, n13248, n13452, n9166, n9756, n12957,
    n13040, n9155, n12942, n9310, n9258, n12953, n9755, n12940, n13171,
    n12881, n9206, n12939, n13357, n9087, n12849, n9327, n12847, n8485,
    n8996, n12873, n9204, n13322, n13349, n9304, n9325, n8428, n13089,
    n8994, n9182, n12767, n8427, n13088, n13157, n12785, n9323, n12753,
    n12766, n8940, n9180, n8992, n8991, n12803, n8800, n9178, n13156,
    n9322, n8890, n12789, n12781, n12751, n9081, n13085, n13230, n12780,
    n12996, n13153, n12920, n9177, n12750, n12919, n12796, n12662, n12995,
    n12871, n12720, n12739, n12897, n13082, n12820, n12679, n12992, n12793,
    n12916, n12526, n12815, n12896, n12475, n12674, n12870, n12715, n12714,
    n12673, n12832, n12483, n12517, n13520, n12471, n12489, n12867, n12445,
    n12893, n12506, n12535, n12829, n12497, n12443, n12049, n12615, n12442,
    n12101, n12496, n12825, n12044, n12700, n12655, n11597, n11844, n8486,
    n11768, n12469, n12611, n11757, n11945, n13213, n11766, n12822, n13194,
    n11841, n11588, n11622, n11943, n8476, n11978, n13407, n11765, n13212,
    n11423, n7662, n9736, n13193, n11563, n11899, n7660, n9735, n11556,
    n12026, n12689, n11421, n11973, n11283, n7661, n11246, n13211, n11348,
    n12508, n12687, n11420, n7659, n11885, n13209, n8433, n13107, n9731,
    n12683, n9768, n12413, n11346, n8431, n11916, n8417, n10992, n11548,
    n13072, n11037, n12633, n10996, n9767, n11412, n12213, n13020, n13207,
    n12976, n13205, n12628, n9739, n12396, n13070, n9727, n11035, n13068,
    n9597, n13033, n9596, n12199, n13345, n13280, n12461, n10831, n12434,
    n12653, n12432, n10672, n12627, n13188, n13031, n13066, n9385, n11698,
    n11682, n9764, n13202, n13327, n12574, n12548, n13129, n11666, n7646,
    n13102, n12559, n9595, n11690, n12648, n11711, n11674, n11024, n12109,
    n7645, n12230, n12250, n12222, n12138, n13539, n12266, n12238, n13039,
    n12125, n12956, n11438, n10571, n13271, n12258, n12647, n13325, n11817,
    n13324, n11834, n12924, n13533, n12278, n12117, n11826, n13128, n13130,
    n9583, n13510, n13125, n11861, n9575, n13494, n12879, n8997, n12886,
    n9183, n9328, n11414, n12861, n12943, n12737, n12955, n12563, n11839,
    n13545, n11930, n13444, n12933, n13215, n13036, n12736, n13551, n12609,
    n12211, n11701, n7636, n8076, n11758, n12740, n13148, n9374, n12329,
    n8055, n9382, n12248, n12210, n13078, n9573, n12979, n7588, n9330,
    n9579, n8053, n13243, n9414, n9749, n11613, n12136, n12744, n13449,
    n11882, n12467, n12595, n9568, n13346, n12435, n13443, n8088, n12729,
    n11339, n13409, n11463, n13311, n13489, n12276, n9148, n8077, n9387,
    n9586, n11626, n12986, n13268, n13011, n10665, n12240, n8479, n12058,
    n9168, n9570, n11738, n13425, n9563, n9744, n10908, n11986, n9748,
    n13218, n13513, n9404, n9384, n11624, n12568, n7586, n13388, n13369,
    n13147, n13076, n9411, n12206, n13303, n7973, n13399, n8074, n13428,
    n8087, n13442, n9147, n12888, n12931, n12591, n12855, n11658, n12149,
    n12728, n11503, n11484, n12038, n11915, n11946, n9181, n11977, n12606,
    n9326, n12412, n12768, n12203, n11995, n9577, n12037, n9403, n11747,
    n13413, n12504, n12592, n9144, n11914, n11447, n11985, n12590, n9771,
    n13441, n9314, n12816, n12850, n12158, n13396, n12848, n13384, n12395,
    n10632, n7585, n8085, n11735, n12778, n13144, n11583, n9333, n13288,
    n12310, n12055, n13497, n11937, n12326, n11502, n9146, n10330, n11976,
    n12144, n11461, n9562, n8056, n9130, n12981, n11171, n12067, n12909,
    n9347, n8165, n12414, n9564, n11971, n11936, n12499, n10889, n12155,
    n12064, n12431, n7007, n12323, n13557, n11495, n12604, n7582, n7971,
    n12775, n7640, n9354, n10800, n13300, n12834, n10630, n10510, n12839,
    n7635, n9184, n11253, n10602, n10906, n11264, n11300, n11459, n12300,
    n12397, n9781, n11744, n12713, n11311, n10560, n13110, n12408, n11382,
    n12493, n13500, n12672, n12200, n9129, n11994, n11363, n13249, n10508,
    n10495, n12141, n10547, n9365, n11732, n11446, n8037, n13479, n13359,
    n10558, n11479, n12833, n11981, n12773, n11959, n11894, n12306, n7638,
    n8173, n12052, n12492, n10904, n7969, n10786, n13000, n12197, n7634,
    n12783, n12201, n10600, n13423, n10798, n10557, n9779, n11290, n12304,
    n7633, n11430, n12514, n10506, n10654, n13524, n11383, n11275, n10887,
    n11614, n12722, n7626, n12523, n11731, n9557, n12140, n8026, n9128,
    n11980, n8027, n12051, n10796, n10538, n10312, n11427, n10692, n12837,
    n13415, n10536, n10614, n13378, n9364, n13531, n10583, n13001, n9369,
    n9560, n9121, n11606, n11918, n10525, n9124, n12612, n11475, n12043,
    n12128, n7629, n10652, n10396, n7639, n13563, n11476, n13555, n13549,
    n12593, n10395, n10496, n12999, n7628, n11443, n12028, n12600, n10651,
    n13049, n10304, n9127, n9589, n10535, n12944, n9368, n7984, n13299,
    n12721, n10794, n9205, n12635, n11546, n9120, n13251, n7556, n7595,
    n7538, n12577, n10597, n13138, n13507, n12285, n8144, n13504, n11442,
    n10533, n13340, n8132, n12617, n11712, n10649, n12949, n12936, n9319,
    n7537, n12298, n10331, n13559, n11655, n13185, n12154, n13229, n12968,
    n10694, n13169, n10581, n9551, n9161, n13355, n10673, n10613, n13099,
    n13016, n12057, n12063, n11743, n12472, n12764, n10555, n13183, n11737,
    n13333, n13475, n12907, n8965, n9754, n10504, n13293, n12946, n12148,
    n10797, n11155, n11494, n8954, n13334, n12053, n10928, n12801, n10492,
    n13176, n12636, n11733, n12543, n10449, n10444, n10403, n10458, n10419,
    n10436, n12147, n10427, n10415, n10411, n12142, n10431, n10440, n8964,
    n10453, n12338, n10407, n10423, n9163, n13571, n8128, n10781, n11810,
    n11636, n10169, n11456, n7423, n10677, n12322, n11992, n11714, n12805,
    n13472, n13199, n10456, n11591, n12308, n11627, n9541, n13391, n13467,
    n13565, n10451, n10080, n10079, n7410, n7536, n12490, n9539, n9705,
    n8972, n13348, n10674, n9598, n7935, n7590, n7650, n8951, n7988,
    n12307, n7664, n9497, n10242, n9100, n8496, n9456, n7995, n9536, n9302,
    n10865, n7560, n9075, n9496, n9298, n10211, n9251, n8123, n9249, n9073,
    n9416, n8933, n7485, n9297, n7540, n7378, n9208, n7488, n9070, n10857,
    n8974, n12476, n9103, n7421, n8930, n8749, n8707, n8789, n8944, n7561,
    n8968, n12527, n8668, n9498, n7370, n8892, n9299, n9248, n9455, n7399,
    n8629, n8666, n7484, n8582, n10468, n7480, n7419, n7570, n8751, n7368,
    n9067, n8627, n9139, n7367, n7381, n8711, n10077, n8084, n7474, n8081,
    n7389, n9096, n8821, n8541, n7362, n8143, n8670, n7405, n7964, n7366,
    n8116, n7371, n8345, n8071, n7468, n7513, n7417, n8122, n10983, n8141,
    n7341, n7369, n10824, n8430, n8156, n8663, n8059, n7360, n7374, n7402,
    n10821, n7445, n8044, n8342, n8172, n8229, n7623, n8306, n7314, n7448,
    n7433, n7507, n8041, n8384, n8472, n8046, n8421, n7321, n7968, n7472,
    n7384, n8493, n8537, n7954, n7993, n8154, n9500, n7346, n8803, n8624,
    n8070, n8130, n9391, n8830, n7991, n8881, n8827, n9197, n8813, n8032,
    n8884, n9194, n8139, n8848, n8110, n8083, n8872, n7461, n7388, n9131,
    n8164, n7435, n9457, n8851, n8869, n7385, n7966, n8842, n8170, n8875,
    n8309, n7442, n8949, n8854, n7432, n8274, n9711, n8833, n8845, n8878,
    n7930, n8266, n8857, n8839, n8191, n7933, n7313, n8264, n8863, n8836,
    n8182, n13186, n8866, n7471, n9394, n7616, n8341, n8860, n8492, n9418,
    n7431, n8747, n8705, n7396, n8068, n9093, n7428, n8787, n7436, n8928,
    n8825, n8019, n8189, n8501, n8272, n7992, n8193, n7926, n8580, n8308,
    n8263, n8109, n8422, n8162, n8180, n8152, n7430, n8092, n8344, n7333,
    n8491, n8819, n8002, n7318, n7335, n9110, n7395, n9707, n10240, n7356,
    n7337, n7464, n8065, n8812, n7508, n9132, n8228, n8058, n8488, n7315,
    n7929, n8418, n8376, n8004, n9723, n7702, n7950, n10245, n10748, n8260,
    n7732, n8226, n7332, n7792, n7731, n7762, n7701, n7823, n8267, n7703,
    n7117, n7822, n8259, n7885, n7330, n7917, n8258, n7886, n7793, n8413,
    n7853, n7852, n7763, n7918, n8414, n7722, n7723, n7884, n7310, n7309,
    n7836, n7790, n7883, n7777, n7902, n7851, n7916, n7850, n7791, n7901,
    n7776, n7733, n8227, n7806, n7761, n7683, n7807, n7821, n7760, n7697,
    n7746, n7696, n7213, n7212, n8261, n7227, n7226, n7820, n7747, n8256,
    n7837, n8257, n7870, n7245, n7915, n8242, n7244, n7869, n8243, n7259,
    n7258, n7196, n7237, n7829, n7054, n7243, n7720, n7236, n7818, n7137,
    n7862, n7819, n7721, n7812, n7729, n7504, n7913, n7700, n7156, n7813,
    n7728, n7694, n7758, n7804, n7695, n7759, n7805, n7799, n7688, n7689,
    n7798, n7093, n7709, n7848, n7077, n7849, n7708, n7842, n7893, n7062,
    n7843, n7881, n7900, n7834, n7835, n7307, n7899, n7882, n7875, n7876,
    n7113, n7867, n7715, n7284, n7828, n7908, n7868, n7907, n7894, n7256,
    n7257, n7714, n7251, n7177, n7914, n7861, n7774, n8184, n7775, n7744,
    n7745, n7738, n7782, n7679, n7788, n7739, n7768, n7753, n7682, n7789,
    n7769, n7752, n7327, n7064, n7811, n7103, n7202, n7272, n7271, n7282,
    n7281, n7889, n7296, n7295, n7306, n7247, n7305, n7892, n7891, n7503,
    n7239, n7896, n7895, n7234, n7898, n7897, n7052, n7904, n7903, n7053,
    n7041, n7906, n7905, n7783, n7042, n7910, n7678, n7699, n7698, n8176,
    n13417, n7276, n7275, n7280, n11877, n7233, n8378, n7304, n7269,
    n10585, n7290, n10489, n7300, n7293, n7265, n7680, n7270, n7264, n9672,
    n7289, n12690, n12691, n7493, n10893, n7478, n7502, n11700, n7641,
    n7456, n11269, n12271, n7051, n7046, n7047, n7040, n10615, n7035,
    n7036, n7890, n7909, n7810, n7165, n7192, n8270, n7140, n7121, n7166,
    n7189, n7133, n7172, n7120, n7149, n9647, n9673, n7139, n8167, n7171,
    n7129, n7125, n7162, n7184, n7163, n8959, n7143, n7182, n7174, n7153,
    n12243, n11284, n7124, n7181, n7130, n8187, n11247, n7455, n7173,
    n7050, n12562, n7132, n8943, n11258, n7325, n9535, n7477, n7499,
    n10074, n11357, n7279, n7152, n11445, n7492, n12131, n8159, n7303,
    n7039, n10485, n7323, n10374, n13515, n10486, n10034, n9789, n11809,
    n7043, n8146, n11480, n7665, n8958, n12821, n8269, n10638, n8586,
    n11488, n12502, n10490, n11628, n12324, n11497, n11813, n7393, n13257,
    n13112, n8134, n8891, n8963, n9056, n10637, n9058, n7497, n11478,
    n12681, n13498, n9757, n9782, n13505, n13496, n13447, n13495, n13476,
    n9769, n13466, n13488, n9554, n13347, n13362, n13458, n9760, n13246,
    n13438, n13454, n13381, n9580, n13307, n13170, n13149, n13245, n13261,
    n9388, n13220, n13404, n13305, n13216, n13159, n9409, n13287, n13395,
    n13058, n13281, n12921, n13115, n9386, n9338, n12872, n12898, n13393,
    n13007, n12987, n9738, n13100, n13478, n13108, n9737, n13184, n9337,
    n13021, n9552, n13017, n13195, n12969, n13238, n13073, n12977, n13450,
    n13094, n9546, n12925, n13093, n12887, n13172, n12908, n9306, n13034,
    n9331, n13092, n12880, n9254, n12950, n9543, n9153, n12962, n9083,
    n12937, n12860, n12945, n13356, n13320, n12901, n9202, n12845, n12899,
    n13319, n9143, n12854, n9252, n12763, n8936, n8425, n13083, n12787,
    n13228, n8809, n8795, n12800, n9250, n9320, n8987, n12747, n12777,
    n9175, n13151, n13525, n8998, n12738, n12660, n12701, n12813, n12989,
    n8976, n8973, n12791, n12914, n12665, n12988, n12891, n12480, n13532,
    n12470, n8975, n12533, n12703, n12864, n12487, n12516, n12656, n12863,
    n13526, n12823, n12097, n12046, n12494, n12039, n12439, n12610, n11755,
    n12528, n11595, n12478, n8424, n12694, n11929, n11585, n8474, n11840,
    n12602, n11619, n12438, n13401, n11762, n13445, n11891, n8423, n11838,
    n8500, n13191, n12748, n7649, n8432, n12686, n11417, n11243, n7654,
    n11280, n13343, n12742, n12411, n13308, n13106, n12685, n13189, n11241,
    n10990, n13141, n13328, n10994, n13019, n12474, n12693, n12440, n12975,
    n12692, n13131, n13075, n11240, n13366, n13204, n13538, n13365, n13206,
    n10828, n11763, n11661, n13065, n13067, n11669, n11862, n11685, n10984,
    n12541, n9576, n7663, n12552, n7643, n12923, n12954, n13028, n9398,
    n12972, n13127, n12745, n12819, n9582, n9313, n8482, n11859, n10825,
    n11028, n12858, n12959, n12878, n12885, n13023, n12941, n13509, n9150,
    n9207, n9203, n13493, n9142, n13289, n9187, n12932, n9591, n12890,
    n11178, n8040, n12608, n13219, n11608, n8093, n12911, n12856, n12732,
    n12704, n12818, n12978, n11295, n12268, n9381, n9378, n8052, n12982,
    n9413, n9329, n9186, n13402, n8094, n12678, n12436, n9179, n12731,
    n11873, n11706, n12910, n13385, n8889, n9373, n11831, n12127, n12743,
    n11248, n12466, n11358, n12677, n10350, n8051, n12605, n11259, n11944,
    n12852, n8072, n7972, n8183, n9745, n9743, n9566, n13403, n13241,
    n13302, n12984, n9407, n13286, n13146, n9185, n9324, n13278, n11623,
    n9747, n11306, n9741, n9200, n13240, n13217, n10460, n9122, n8049,
    n8038, n8029, n13054, n13487, n8888, n13398, n13434, n11377, n8887,
    n13121, n12712, n11270, n13265, n10903, n10351, n9171, n12786, n9401,
    n11285, n12810, n8039, n8993, n13256, n8158, n13060, n8017, n8036,
    n8064, n11477, n8166, n8048, n10598, n12427, n13114, n8035, n11547,
    n10493, n8047, n13118, n12667, n8157, n12705, n9344, n13523, n7584,
    n11966, n10545, n11317, n10305, n12481, n12664, n10676, n10783, n10901,
    n10681, n7600, n8145, n10548, n7627, n10621, n12030, n10320, n12663,
    n13008, n9778, n10590, n12047, n9165, n9588, n10541, n13371, n9775,
    n13250, n13298, n10523, n9361, n11846, n7577, n10335, n12782, n12765,
    n11847, n11707, n11931, n12498, n10319, n11316, n12842, n8986, n10526,
    n7956, n11244, n9734, n12926, n11718, n12040, n10989, n9191, n9174,
    n13071, n10642, n7983, n11594, n11586, n12716, n7593, n12675, n8129,
    n7555, n10779, n13528, n9321, n9176, n8990, n12417, n8102, n13069,
    n13029, n7006, n13210, n12938, n11326, n10321, n12554, n12369, n10544,
    n12358, n12569, n12538, n12346, n12312, n13460, n8484, n10233, n9545,
    n12334, n8808, n10234, n11646, n12317, n7948, n13335, n12330, n10442,
    n11620, n8989, n7949, n12749, n12994, n9544, n12792, n12794, n10586,
    n11422, n11347, n12098, n8426, n13175, n12752, n10447, n8935, n10425,
    n12444, n9253, n10405, n10434, n9305, n10438, n10413, n10417, n10421,
    n10203, n12828, n8117, n9082, n12895, n8794, n8011, n10455, n12799,
    n10409, n10429, n8014, n10450, n10401, n11767, n12869, n7947, n7990,
    n9108, n11481, n7422, n11632, n10402, n10215, n10426, n10414, n10410,
    n10435, n10430, n13091, n10439, n10418, n9693, n10422, n10406, n9105,
    n10616, n8126, n13164, n7955, n7543, n9106, n9537, n12960, n11830,
    n12588, n7591, n10488, n7987, n12900, n7941, n8127, n9098, n9704,
    n7542, n9079, n7539, n7936, n7486, n11553, n9071, n7557, n8999, n8931,
    n8495, n8709, n8932, n11402, n7505, n7489, n12699, n12654, n8790,
    n7377, n11319, n10038, n7495, n8750, n7392, n9101, n8708, n9114,
    n10035, n7475, n7463, n8824, n8073, n8581, n8664, n8630, n9247, n10938,
    n7379, n7452, n8947, n8626, n7458, n7416, n8583, n7970, n7407, n9097,
    n7386, n7446, n11023, n9135, n7940, n7986, n9134, n7473, n12025,
    n10032, n8538, n7361, n7946, n7406, n7934, n11239, n7339, n8499, n7994,
    n7451, n8822, n9095, n10391, n7412, n7376, n7347, n7444, n8818, n7466,
    n7958, n7462, n7352, n9156, n7483, n7418, n7359, n7408, n7937, n7354,
    n7364, n8140, n8121, n7945, n7967, n8069, n7439, n8471, n8153, n8536,
    n8802, n7963, n7351, n7336, n9094, n7230, n7425, n8380, n8539, n9117,
    n7344, n7938, n8419, n7350, n7957, n7953, n7944, n7343, n7357, n8114,
    n8852, n8843, n7952, n8879, n8861, n8828, n8882, n8837, n7962, n8864,
    n7199, n8147, n8870, n7319, n7482, n8383, n7931, n7443, n8873, n8834,
    n8846, n8867, n8855, n8811, n7460, n8831, n8138, n7311, n7518, n8169,
    n8849, n8858, n8840, n7438, n10241, n8876, n8080, n7467, n8416, n8151,
    n8489, n7615, n8435, n8060, n9074, n8490, n8535, n8703, n8746, n9259,
    n8667, n8179, n7481, n8188, n8066, n8108, n8579, n7312, n8379, n7923,
    n8161, n7320, n7856, n8786, n7429, n7413, n8470, n8120, n8628, n7317,
    n7427, n7961, n7925, n8271, n8841, n8829, n9210, n8816, n8853, n8856,
    n7459, n8950, n8859, n8835, n8850, n8817, n7613, n8192, n8101, n8810,
    n8575, n7924, n8868, n8381, n11637, n8792, n8838, n8832, n9686, n8826,
    n7922, n8031, n8847, n8273, n7345, n8862, n8801, n8865, n7996, n7887,
    n8844, n8815, n8343, n8042, n7921, n11156, n8265, n10499, n7231, n8003,
    n8225, n7261, n7057, n10574, n8190, n8304, n7260, n7331, n8338, n8303,
    n7114, n7198, n7115, n7031, n7071, n8181, n7101, n7070, n7085, n7030,
    n7197, n7084, n7100, n7178, n7205, n7210, n12347, n8171, n7204, n7055,
    n7211, n12345, n7112, n12359, n7157, n7136, n12313, n7092, n7225,
    n12301, n7098, n7224, n7107, n12333, n12335, n7218, n7023, n7099,
    n7022, n7082, n7029, n7083, n7106, n12549, n7028, n7219, n7195, n12555,
    n7076, n12560, n7242, n7063, n12368, n7250, n7308, n7283, n12544,
    n12570, n12357, n12536, n12370, n7069, n7068, n7194, n7186, n7168,
    n7111, n7187, n12754, n7109, n7104, n7674, n7175, n7110, n7072, n7176,
    n7074, n7108, n8163, n7167, n7089, n7065, n7154, n7155, n7091, n7145,
    n7060, n7146, n7080, n7067, n7061, n7134, n7090, n7135, n7058, n7066,
    n7059, n8953, n7126, n7081, n7127, n7102, n7078, n7193, n7079, n7795,
    n7911, n7912, n7794, n7846, n7847, n7844, n7845, n7840, n7841, n7838,
    n7839, n7832, n7830, n7826, n7827, n7201, n7200, n7203, n7824, n7726,
    n7206, n7727, n7825, n7724, n7725, n7816, n7817, n7814, n7815, n7808,
    n7809, n7802, n7803, n7800, n7796, n7797, n7209, n7736, n7873, n7878,
    n7874, n7735, n7249, n7773, n7770, n7877, n7737, n7771, n7740, n7248,
    n7743, n7880, n7871, n7742, n7027, n7879, n7872, n7024, n7025, n7749,
    n7766, n7748, n7246, n7020, n7767, n7021, n7866, n7253, n7019, n7255,
    n7222, n7863, n7751, n7864, n7750, n7686, n7223, n7254, n7859, n7755,
    n7860, n7858, n7754, n7684, n7220, n7757, n7772, n7756, n7764, n7238,
    n7685, n7232, n7716, n7221, n7208, n7765, n7681, n7235, n7705, n7785,
    n7704, n7217, n7241, n7673, n7787, n7215, n7707, n7780, n7706, n7781,
    n7240, n7214, n7786, n7784, n7778, n7190, n12511, n7150, n7779, n7741,
    n7734, n7144, n7185, n12991, n7002, n7207, n7710, n7216, n7865, n13451,
    n7857, n7801, n7252, n7676, n7677, n7294, n7301, n8178, n7833, n7831,
    n7073, n7075, n8160, n7088, n8155, n7095, n13057, n13306, n13382,
    n9766, n12866, n12840, n12779, n13456, n13363, n12762, n12826, n13508,
    n13006, n13262, n13162, n8585, n7286, n7288, n8195, n9057, n7324,
    n8196, n7454, n11849, n7299, n8262, n7470, n7491, n8168, n8307, n8142,
    n7476, n9855, n7338, n7498, n8551, n7032, n7526, n12835, n12680,
    n11893, n10341, n7003, n10223, n8061, n7391, n12718, n10934, n9140,
    n9138, n11896, n7358, n8194, n7170, n7038, n7034, n7268, n7263, n7602,
    n7123, n7119, n7888, n7928, n7594, n7580, n7579, n9172, n8984, n12576,
    n8823, n8107, n9303, n12696, n12734, n8095, n8086, n8078, n7589,
    n11444, n10690, n12145, n8814, n9318, n12033, n12726, n13196, n9316,
    n9339, n9340, n11589, n11087, n8807, n7322, n13079, n12912, n9332,
    n11940, n13405, n13521, n12524, n12624, n12459, n12646, n11653, n11656,
    n11648, n12295, n11957, n12859, n12853, n12913, n11088, n10867, n13536,
    n10667, n10668, n13542, n10470, n9308, n9256, n9085, n8938, n8798,
    n12658, n12297, n10322, n13152, n12473, n12391, n11649, n9758, n9363,
    n13376, n13375, n13380, n13259, n13258, n13004, n12758, n12760, n9160,
    n12510, n12515, n11892, n11890, n11561, n11560, n11559, n9116, n11576,
    n11395, n12114, n12106, n12122, n12134, n12320, n12341, n12353, n12364,
    n12375, n11454, n11470, n12255, n12263, n12274, n11380, n11868, n11880,
    n12219, n12246, n12227, n12235, n7355, n9641, n7690, n7691, n7693,
    n7692, n7687, n7675, n7713, n7712, n7718, n7719, n7717, n7711, n7348,
    n8020, n9050, n8548, n7960, n8592, n9417, n9209, n8403, n8300, n7976,
    n7450, n7469, n9052, n7179, n7180, n8199, n7188, n7160, n7164, n7161,
    n7044, n7049, n7285, n7291, n7287, n7298, n7302, n7297, n7273, n7278,
    n7277, n7274, n7342, n7372, n8659, n8660, n9490, n8584, n7141, n7142,
    n7138, n7151, n7147, n8590, n7131, n7128, n9296, n8745, n8578, n8465,
    n8375, n8374, n8235, n8241, n8254, n8255, n8248, n13279, n7611, n8043,
    n8034, n7932, n7939, n7951, n7501, n7496, n7500, n7409, n11441, n10898,
    n7169, n7037, n7033, n7266, n7262, n7403, n7404, n7400, n9317, n8434,
    n11717, n9762, n12874, n9389, n8622, n8224, n8207, n8206, n8175, n8137,
    n8174, n10467, n9634, n9540, n7122, n7118, n9548, n9295, n9454, n8969,
    n12707, n8339, n8240, n8249, n8013, n8136, n8113, n13429, n13190,
    n13101, n9198, n9195, n9315, n9192, n12695, n8877, n12733, n8874,
    n9162, n8477, n12771, n11086, n9088, n7612, n10864, n11886, n8057,
    n8075, n11552, n12202, n12207, n11401, n11318, n7541, n10484, n12302,
    n7919, n7583, n8980, n8945, n10043, n9732, n8988, n13338, n13136,
    n13064, n12970, n9717, n12973, n9713, n9397, n12882, n9392, n12947,
    n12948, n12934, n12935, n9173, n8985, n12717, n8871, n8960, n12670,
    n12669, n12607, n11969, n12448, n12644, n12587, n12585, n11948, n9300,
    n8885, n8883, n8966, n8880, n11584, n11590, n10986, n10856, n8820,
    n10932, n9494, n11752, n11647, n8487, n8131, n10297, n13471, n9692,
    n13453, n13332, n13234, n9408, n9405, n13161, n12951, n13352, n13315,
    n9077, n13224, n9383, n13227, n13150, n8710, n12601, n7671, n8382,
    n12463, n7670, n12390, n11645, n10927, n13468, n13400, n9765, n9773,
    n9366, n9201, n13419, n13059, n9375, n12844, n12755, n12761, n11237,
    n12776, n12509, n12770, n12512, n12468, n12491, n12437, n8089, n7316,
    n7624, n11921, n11919, n11558, n13374, n11397, n11432, n11325, n11330,
    n9126, n10582, n10372, n11638, n11458, n11607, n10679, n11376, n10902,
    n10629, n10628, n10617, n10057, n7648, n7449, n10039, n13037, n13022,
    n13506, n12928, n9190, n8962, n12811, n12735, n12725, n13527, n12711,
    n12035, n12613, n12598, n11942, n11934, n12410, n12406, n11909, n11912,
    n12379, n12394, n12389, n12387, n12425, n13440, n13264, n9343, n9342,
    n12045, n12841, n13548, n10352, n13554, n13562, n13181, n13097, n13014,
    n12966, n12905, n12798, n10206, n10283, n10446, n10293, n10273, n13473,
    n13457, n13455, n13168, n13353, n9578, n13225, n13154, n13086, n12917,
    n13056, n12993, n12985, n12990, n12894, n13005, n12868, n9334, n12827,
    n9151, n11939, n12741, n12465, n12441, n12433, n12495, n11764, n12616,
    n11419, n12428, n11344, n12449, n12634, n12575, n10325, n13480, n9349,
    n12838, n12769, n12501, n11928, n11926, n11436, n12003, n12001, n12011,
    n12009, n11989, n11987, n12019, n12017, n11167, n12550, n12539, n12566,
    n12564, n11185, n11659, n11677, n11675, n11683, n11667, n11704, n11702,
    n11693, n11691, n11159, n12181, n12179, n12165, n12163, n12173, n12171,
    n12152, n12150, n12190, n11361, n11492, n11542, n11534, n11526, n11518,
    n11510, n10693, n11007, n10999, n11795, n11771, n11769, n11779, n11741,
    n11739, n11803, n11874, n11787, n12061, n12059, n12074, n12072, n12090,
    n12082, n12650, n12418, n9956, n12632, n12462, n12652, n11657, n11652,
    n12594, n12299, n12296, n11729, n11960, n12702, n13522, n11090, n10868,
    n13537, n13543, n10471, n10935, n13394, n9309, n9257, n9086, n8939,
    n8799, n12659, n12532, n12486, n11025, n10822, n10360, n10172, n10163,
    n10127, n10119, n10107, n10103, n10099, n10095, n10091, n10087, n10123,
    n10083, n10115, n10111, n10167, n10143, n10200, n10155, n10151, n10180,
    n10184, n10135, n10192, n10131, n10147, n10139, n10207, n10176, n10196,
    n10188, n10159, n13570, n13155, n13087, n8429, n7672, n11843, n11842,
    n10569, n10481, n13360, n13503, n13499, n13379, n13260, n13055, n13003,
    n12759, n12784, n12525, n12518, n12505, n11898, n11897, n11562, n12214,
    n11411, n11405, n11582, n11104, n11103, n11092, n11396, n11835, n11833,
    n11818, n11827, n11863, n12116, n12108, n12124, n12137, n12331, n12343,
    n12355, n12366, n12377, n11464, n11472, n12257, n12265, n12277, n11870,
    n11883, n12221, n12249, n12229, n12237, n7004, n7005, n11852, n8018,
    n7008, n10027, n13481, n7009, n12415, n7010, n7011, n7597, n9883,
    n9102, n8970, n8148, n8533, n8268, n8377, n8971, n7012, n9169, n12638,
    n8001, n8067, n8177, n8185, n7013, n7014, n7015, n7016, n9657, n13491,
    n13222, n7017, n7292, n7373, n7855, n7329, n7045, n7183, n8119, n8783,
    n8467, n7148, n8924, n8186, n7487, n7546, n7959, n9572, n10780, n7398,
    n9726, n13163, n9080, n12309, n11483, n10534, n7601, n8796, n12477,
    n10076, n12961, n9301, n8540, n7669, n11593, n10787, n7657, n12963,
    n12790, n10441, n10432, n10826, n11578, n9918, n12676, n9648, n9501,
    n7018, n9053, n9636, n9051, n7267, n9640, n9522, n8587, n7026, n9642,
    n8591, n7056, n9665, n9602, n9599, n9656, n7087, n9662, n9607, n9610,
    n7086, n7614, n7094, n7097, n7096, n7105, n7116, n13389, n7465, n8498,
    n7159, n7158, n7191, n9092, n7229, n7228, n7441, n7394, n7411, n8574,
    n8791, n7326, n7349, n7328, n7334, n7382, n7383, n7401, n8082, n7340,
    n7365, n7353, n7363, n7375, n7380, n7387, n7390, n7397, n8946, n10075,
    n8948, n7516, n9107, n8804, n7414, n7415, n9099, n7420, n7424, n7592,
    n7426, n7434, n7506, n7447, n9111, n7440, n7437, n7453, n7457, n9787,
    n7568, n7567, n7559, n7479, n7558, n7490, n7494, n11440, n11854, n7512,
    n7510, n7509, n7511, n7514, n7515, n7517, n7519, n7520, n7544, n7523,
    n7522, n7524, n7525, n7534, n7545, n7527, n7528, n10363, n7532, n7529,
    n7530, n7531, n7533, n7535, n10362, n7587, n7554, n7547, n7552, n7550,
    n7548, n7549, n7551, n7553, n10338, n7581, n7569, n7566, n10373, n7562,
    n7564, n7563, n7565, n10369, n7575, n11949, n7574, n7572, n7571, n7573,
    n10383, n7576, n7578, n7596, n7598, n7599, n7609, n7604, n7603, n7607,
    n7605, n10055, n7606, n7608, n7610, n7617, n7619, n7618, n7621, n7620,
    n7622, n10071, n7625, n7630, n7632, n8978, n7647, n7642, n10063, n7644,
    n10056, n7651, n7652, n7653, n7655, n7656, n12684, n7658, n12305,
    n10060, n7666, n7668, n7667, n10209, n7730, n7943, n7854, n7920, n8079,
    n7927, n8090, n7942, n7975, n7974, n7965, n8063, n11820, n7982, n7978,
    n7977, n7979, n7980, n7981, n8016, n7985, n10327, n7989, n10886, n8000,
    n7998, n7997, n7999, n10216, n10224, n8007, n8005, n8006, n8010, n8009,
    n10222, n8012, n8015, n10328, n10474, n11845, n8024, n8021, n8022,
    n8023, n8025, n11332, n8028, n10473, n10476, n10565, n8033, n10566,
    n11027, n8050, n12196, n8054, n11029, n11338, n11340, n11413, n11415,
    n11759, n11761, n8096, n8097, n8098, n8099, n12746, n8100, n8478,
    n9633, n9708, n8103, n12292, n8104, n8106, n8105, n8115, n8112, n10213,
    n8124, n8125, n10313, n8149, n8150, n10461, n10666, n8198, n8197,
    n8203, n8201, n8200, n8202, n8205, n8204, n8209, n8208, n8213, n8211,
    n8210, n8212, n8221, n8215, n8214, n8219, n8217, n8216, n8218, n8220,
    n8223, n8222, n8231, n8230, n8233, n8232, n8234, n8237, n8236, n8239,
    n8238, n8245, n8244, n8247, n8246, n8251, n8250, n8253, n8252, n8276,
    n8275, n8280, n8278, n8277, n8279, n8288, n8282, n8281, n8286, n8284,
    n8283, n8285, n8287, n8290, n8289, n8294, n8292, n8291, n8293, n8302,
    n8296, n8295, n8298, n8297, n8299, n8301, n8305, n8311, n8310, n8315,
    n8313, n8312, n8314, n8323, n8317, n8316, n8321, n8319, n8318, n8320,
    n8322, n8325, n8324, n8329, n8327, n8326, n8328, n8337, n8331, n8330,
    n8335, n8333, n8332, n8334, n8336, n8340, n8347, n8346, n8351, n8349,
    n8348, n8350, n8359, n8353, n8352, n8357, n8355, n8354, n8356, n8358,
    n8361, n8360, n8365, n8363, n8362, n8364, n8373, n8367, n8366, n8371,
    n8369, n8368, n8370, n8372, n8386, n8385, n8390, n8388, n8387, n8389,
    n8398, n8392, n8391, n8396, n8394, n8393, n8395, n8397, n8400, n8399,
    n8404, n8402, n8401, n8412, n8406, n8405, n8410, n8408, n8407, n8409,
    n8411, n8415, n8420, n8468, n8475, n8473, n8437, n8436, n8441, n8439,
    n8438, n8440, n8449, n8443, n8442, n8447, n8445, n8444, n8446, n8448,
    n8451, n8450, n8455, n8453, n8452, n8454, n8463, n8457, n8456, n8461,
    n8459, n8458, n8460, n8462, n8464, n8466, n8469, n8480, n8481, n8483,
    n8494, n8497, n8503, n8502, n8507, n8505, n8504, n8506, n8515, n8509,
    n8508, n8513, n8511, n8510, n8512, n8514, n8531, n8517, n8516, n8521,
    n8519, n8518, n8520, n8529, n8523, n8522, n8527, n8525, n8524, n8526,
    n8528, n8530, n8532, n8534, n8543, n8542, n8547, n8545, n8544, n8546,
    n8573, n8550, n8549, n8555, n8553, n8552, n8554, n8571, n8557, n8556,
    n8561, n8559, n8558, n8560, n8569, n8563, n8562, n8567, n8565, n8564,
    n8566, n8568, n8570, n8572, n9696, n8576, n8577, n8589, n8588, n8597,
    n8595, n8594, n8596, n8601, n8599, n8598, n8600, n8621, n8603, n8602,
    n8607, n8605, n8604, n8606, n8615, n8609, n8608, n8613, n8611, n8610,
    n8612, n8614, n8619, n8617, n8616, n8618, n8620, n8623, n8625, n8632,
    n8631, n8636, n8634, n8633, n8635, n8644, n8638, n8637, n8642, n8640,
    n8639, n8641, n8643, n8646, n8645, n8650, n8648, n8647, n8649, n8658,
    n8652, n8651, n8656, n8654, n8653, n8655, n8657, n8661, n8669, n8662,
    n8665, n8672, n8671, n8676, n8674, n8673, n8675, n8684, n8678, n8677,
    n8682, n8680, n8679, n8681, n8683, n8700, n8686, n8685, n8690, n8688,
    n8687, n8689, n8698, n8692, n8691, n8696, n8694, n8693, n8695, n8697,
    n8699, n8701, n8706, n8702, n8704, n8713, n8712, n8717, n8715, n8714,
    n8716, n8725, n8719, n8718, n8723, n8721, n8720, n8722, n8724, n8741,
    n8727, n8726, n8731, n8729, n8728, n8730, n8739, n8733, n8732, n8737,
    n8735, n8734, n8736, n8738, n8740, n8742, n8748, n8743, n8744, n8753,
    n8752, n8757, n8755, n8754, n8756, n8765, n8759, n8758, n8763, n8761,
    n8760, n8762, n8764, n8781, n8767, n8766, n8771, n8769, n8768, n8770,
    n8779, n8773, n8772, n8777, n8775, n8774, n8776, n8778, n8780, n8782,
    n8788, n8784, n8785, n8793, n13177, n8797, n8805, n12208, n11887,
    n10987, n11238, n8967, n8886, n8894, n8893, n8898, n8896, n8895, n8897,
    n8906, n8900, n8899, n8904, n8902, n8901, n8903, n8905, n8922, n8908,
    n8907, n8912, n8910, n8909, n8911, n8920, n8914, n8913, n8918, n8916,
    n8915, n8917, n8919, n8921, n8923, n8929, n8927, n8925, n8926, n8934,
    n8937, n8961, n9951, n12603, n12029, n12380, n12630, n11911, n11975,
    n8941, n12447, n9994, n11654, n8942, n8955, n9091, n10061, n8952,
    n11630, n12651, n12631, n9984, n8956, n8957, n8995, n13330, n8977,
    n8982, n8979, n8981, n8983, n13197, n9078, n9001, n9000, n9005, n9003,
    n9002, n9004, n9029, n9007, n9006, n9011, n9009, n9008, n9010, n9019,
    n9013, n9012, n9017, n9015, n9014, n9016, n9018, n9027, n9021, n9020,
    n9025, n9023, n9022, n9024, n9026, n9028, n9031, n9030, n9035, n9033,
    n9032, n9034, n9066, n9037, n9036, n9041, n9039, n9038, n9040, n9049,
    n9043, n9042, n9047, n9045, n9044, n9046, n9048, n9064, n9055, n9054,
    n9062, n9060, n9059, n9061, n9063, n9065, n9068, n9076, n9069, n9072,
    n9084, n11406, n9119, n11557, n11920, n12500, n12513, n12519, n12774,
    n9089, n9090, n9104, n9109, n9125, n13043, n9112, n9113, n9115, n11324,
    n11579, n9118, n11569, n11407, n12520, n12836, n9348, n9357, n9360,
    n9123, n13377, n9157, n9133, n9137, n9136, n9141, n9145, n9152, n9149,
    n12830, n9154, n9159, n9158, n9164, n9170, n9311, n9189, n9188, n9193,
    n9199, n9196, n12875, n9212, n9211, n9216, n9214, n9213, n9215, n9224,
    n9218, n9217, n9222, n9220, n9219, n9221, n9223, n9240, n9226, n9225,
    n9230, n9228, n9227, n9229, n9238, n9232, n9231, n9236, n9234, n9233,
    n9235, n9237, n9239, n9260, n9241, n9242, n9245, n9243, n9244, n9246,
    n9255, n9262, n9261, n9266, n9264, n9263, n9265, n9270, n9268, n9267,
    n9269, n9290, n9272, n9271, n9276, n9274, n9273, n9275, n9284, n9278,
    n9277, n9282, n9280, n9279, n9281, n9283, n9288, n9286, n9285, n9287,
    n9289, n9291, n9294, n9292, n9293, n9307, n9312, n9335, n12889, n9336,
    n9341, n9356, n9351, n9350, n9352, n9353, n13272, n13484, n12998,
    n9558, n13048, n13053, n9561, n13372, n13410, n9555, n9776, n9359,
    n9358, n9362, n9559, n13044, n13373, n9367, n13274, n9772, n13501,
    n9371, n9370, n9372, n13109, n13002, n9567, n9379, n13111, n9376,
    n9377, n13270, n9380, n13283, n13370, n9406, n9390, n12883, n9393,
    n9714, n9396, n9395, n13244, n9410, n13239, n9415, n9780, n9412, n9420,
    n9419, n9424, n9422, n9421, n9423, n9432, n9426, n9425, n9430, n9428,
    n9427, n9429, n9431, n9448, n9434, n9433, n9438, n9436, n9435, n9437,
    n9446, n9440, n9439, n9444, n9442, n9441, n9443, n9445, n9447, n9458,
    n9449, n9450, n9452, n9451, n9453, n9460, n9459, n9464, n9462, n9461,
    n9463, n9488, n9466, n9465, n9470, n9468, n9467, n9469, n9478, n9472,
    n9471, n9476, n9474, n9473, n9475, n9477, n9486, n9480, n9479, n9484,
    n9482, n9481, n9483, n9485, n9487, n9499, n9489, n9495, n9493, n9491,
    n9492, n9503, n9502, n9507, n9505, n9504, n9506, n9515, n9509, n9508,
    n9513, n9511, n9510, n9512, n9514, n9532, n9517, n9516, n9521, n9519,
    n9518, n9520, n9530, n9524, n9523, n9528, n9526, n9525, n9527, n9529,
    n9531, n9635, n9533, n9542, n9534, n9538, n13132, n9547, n9550, n13133,
    n9549, n9556, n9565, n9571, n13077, n13414, n9740, n13314, n9581,
    n13026, n13126, n9587, n9888, n13200, n9594, n9590, n9592, n9593,
    n9601, n9600, n9606, n9604, n9603, n9605, n9616, n9609, n9608, n9614,
    n9612, n9611, n9613, n9615, n9632, n9618, n9617, n9622, n9620, n9619,
    n9621, n9630, n9624, n9623, n9628, n9626, n9625, n9627, n9629, n9631,
    n9682, n9681, n9695, n9638, n9637, n9646, n9639, n9644, n9643, n9645,
    n9652, n9650, n9649, n9651, n9679, n9655, n9654, n9661, n9659, n9658,
    n9660, n9671, n9664, n9663, n9669, n9667, n9666, n9668, n9670, n9677,
    n9675, n9674, n9676, n9678, n9694, n9683, n9680, n9685, n9684, n9691,
    n9689, n9687, n9688, n9690, n9697, n9703, n9701, n9699, n9700, n9702,
    n9706, n13174, n9712, n9710, n9709, n13464, n12971, n9716, n9715,
    n9761, n9719, n9718, n9720, n13187, n9722, n9721, n13103, n9725, n9724,
    n9729, n9728, n9730, n9733, n9742, n9746, n9750, n9751, n9753, n9752,
    n13297, n13301, n13273, n9759, n9763, n9770, n9774, n9777, n9783,
    n10023, n9784, n9861, n9786, n9785, n9788, n9791, n9790, n13517, n9793,
    n9792, n9795, n9794, n9797, n9796, n9799, n9798, n9801, n9800, n9803,
    n9802, n9807, n9805, n9804, n9806, n9815, n9809, n9808, n9813, n9811,
    n9810, n9812, n9814, n9831, n9817, n9816, n9821, n9819, n9818, n9820,
    n9829, n9823, n9822, n9827, n9825, n9824, n9826, n9828, n9830, n9850,
    n9852, n9839, n9836, n9849, n9833, n9840, n9832, n9834, n9835, n9837,
    n9838, n9844, n9841, n9845, n9842, n9843, n9846, n9848, n9847, n9851,
    n9854, n9853, n10018, n10011, n9858, n9863, n10012, n9856, n9864,
    n9857, n9860, n9859, n9862, n9866, n9865, n9867, n9868, n13514, n9870,
    n9869, n12031, n10001, n9872, n9999, n9871, n9874, n9873, n9876, n9897,
    n9875, n9878, n9877, n9880, n13221, n9879, n9882, n9881, n9885, n9884,
    n9887, n9886, n9890, n9889, n9892, n9891, n9894, n9893, n9896, n9895,
    n9899, n9898, n9901, n9900, n13035, n9903, n9902, n9905, n9904, n9907,
    n9906, n9909, n9908, n9957, n9911, n13024, n9910, n9913, n9912, n9915,
    n13124, n9914, n9917, n9916, n9920, n12817, n9919, n9922, n9921, n9967,
    n9924, n9989, n9923, n9926, n9925, n10000, n9928, n9927, n9930, n9929,
    n9932, n11901, n9931, n9934, n9933, n9936, n9935, n9938, n9937, n9940,
    n9939, n9942, n9941, n9944, n9943, n9946, n9945, n9962, n9948, n9947,
    n9950, n9949, n9953, n9952, n9955, n9954, n9959, n9958, n9961, n9960,
    n12284, n9964, n9963, n9966, n9965, n9969, n9968, n9971, n9970, n9973,
    n9972, n9975, n9974, n9977, n9976, n9979, n9978, n9981, n9980, n9983,
    n9982, n9986, n9985, n9988, n9987, n9991, n9990, n9993, n9992, n9996,
    n9995, n9998, n9997, n10003, n10002, n10005, n10004, n10006, n10007,
    n10008, n10010, n10009, n10017, n10015, n10013, n10014, n10016, n10022,
    n10020, n10019, n10021, n10025, n10024, n10028, n10026, n10031, n10029,
    n10030, n11631, n10037, n10036, n10042, n10040, n10041, n10069, n10044,
    n10049, n10048, n10046, n10047, n10051, n10050, n10053, n10052, n10054,
    n10059, n10058, n10062, n10064, n10068, n10202, n10065, n10066, n10067,
    n10073, n10070, n10072, n10078, n10082, n10081, n10084, n10086, n10085,
    n10088, n10090, n10089, n10092, n10094, n10093, n10096, n10098, n10097,
    n10100, n10102, n10101, n10104, n10106, n10105, n10108, n10110, n10109,
    n10112, n10114, n10113, n10116, n10118, n10117, n10120, n10122, n10121,
    n10124, n10126, n10125, n10128, n10130, n10129, n10132, n10134, n10133,
    n10136, n10138, n10137, n10140, n10142, n10141, n10144, n10146, n10145,
    n10148, n10150, n10149, n10152, n10154, n10153, n10156, n10158, n10157,
    n10160, n10162, n10161, n10164, n10166, n10165, n10168, n10171, n10170,
    n10173, n10175, n10174, n10177, n10179, n10178, n10181, n10183, n10182,
    n10185, n10187, n10186, n10189, n10191, n10190, n10193, n10195, n10194,
    n10197, n10199, n10198, n10201, n10205, n10204, n10208, n10210, n10221,
    n10212, n10214, n10219, n11390, n11388, n10217, n10218, n10220, n10225,
    n10226, n10229, n10227, n10228, n11093, n10232, n11094, n10230, n10231,
    n10239, n10237, n10235, n10236, n10238, n10244, n10243, n10246, n13566,
    n10248, n10247, n10249, n10251, n10250, n10252, n10254, n10253, n10255,
    n10257, n10256, n10258, n10260, n10259, n10261, n10263, n10262, n10264,
    n10266, n10265, n10267, n10269, n10268, n10270, n10272, n10271, n10274,
    n10276, n10275, n10277, n10279, n10278, n10280, n10282, n10281, n10284,
    n10286, n10285, n10287, n10289, n10288, n10290, n10292, n10291, n10294,
    n10296, n10295, n10299, n12099, n10298, n10399, n10301, n10300, n10303,
    n10302, n10454, n10309, n10307, n10306, n10308, n10311, n10310, n10315,
    n10859, n10314, n10317, n10316, n11567, n10318, n10326, n10324, n10323,
    n11573, n10329, n12507, n10333, n10332, n10334, n10336, n10337, n10349,
    n10346, n10370, n10339, n10371, n10344, n10342, n10343, n10345, n10347,
    n10348, n10355, n10353, n10354, n10357, n10356, n10359, n10358, n10361,
    n10365, n10364, n10366, n10368, n10367, n10379, n10377, n10375, n10376,
    n10378, n10380, n10382, n10381, n10387, n10385, n10384, n10386, n10388,
    n10390, n10389, n10393, n10392, n10394, n10398, n10397, n10400, n10404,
    n10408, n10412, n10416, n11753, n10420, n10459, n10424, n10428, n10433,
    n10437, n10443, n10445, n10448, n10452, n10457, n10464, n10462, n10463,
    n10466, n10465, n12286, n10469, n10472, n10482, n10478, n10475, n11333,
    n10477, n10480, n10479, n10483, n11321, n11699, n10503, n10487, n10491,
    n10543, n12316, n11828, n10542, n10494, n10498, n12537, n10497, n10501,
    n10747, n10500, n10502, n10512, n10505, n10507, n10509, n10511, n10519,
    n10514, n10513, n10517, n10516, n10518, n10521, n10520, n11872, n10532,
    n10584, n11730, n12287, n10522, n10524, n10528, n12092, n10527, n10530,
    n10529, n10531, n10540, n10537, n10539, n12561, n10554, n11979, n10546,
    n10550, n10549, n10552, n10551, n10553, n10562, n10556, n10559, n10561,
    n10564, n10563, n11424, n11429, n10567, n10568, n10570, n10578, n10573,
    n10572, n10576, n10575, n10577, n10580, n10579, n12126, n10596, n12050,
    n10587, n10589, n10588, n10592, n12239, n10591, n10594, n10593, n10595,
    n10604, n10599, n10601, n10603, n10610, n10606, n10605, n10608, n10607,
    n10609, n10612, n10611, n10627, n10675, n10892, n10618, n10620, n10619,
    n10623, n11301, n10622, n10625, n10624, n10626, n10634, n10631, n10633,
    n10636, n12183, n10648, n10784, n11451, n11457, n10639, n10641, n10640,
    n10644, n10643, n10646, n10645, n10647, n10656, n10650, n10653, n10655,
    n10662, n10658, n10657, n10660, n10659, n10661, n10664, n10663, n10670,
    n10669, n10671, n10688, n11489, n10680, n10684, n10678, n10683, n10682,
    n10686, n10685, n10687, n10696, n10689, n10691, n10695, n10702, n10698,
    n10697, n10700, n10699, n10701, n10704, n10703, n10710, n10706, n10705,
    n10708, n10707, n10709, n10712, n10711, n10716, n10714, n10713, n10715,
    n10720, n10718, n10717, n10719, n10724, n10722, n10721, n10723, n10728,
    n10726, n10725, n10727, n10732, n10730, n10729, n10731, n10736, n10734,
    n10733, n10735, n10740, n10738, n10737, n10739, n10744, n10742, n10741,
    n10743, n10752, n10746, n10745, n10750, n12350, n10749, n10751, n10754,
    n10753, n10760, n10756, n10755, n10758, n10757, n10759, n10762, n10761,
    n10766, n10764, n10763, n10765, n10770, n10768, n10767, n10769, n10776,
    n10772, n10771, n10774, n10773, n10775, n10778, n10777, n10793, n10782,
    n12139, n10785, n10789, n12267, n10788, n10791, n10790, n10792, n10802,
    n10795, n10799, n10801, n10808, n10804, n10803, n10806, n10805, n10807,
    n10810, n10809, n10814, n10812, n10811, n10813, n10818, n10816, n10815,
    n10817, n10820, n10819, n10823, n10829, n10827, n10830, n10837, n10833,
    n10832, n10835, n10834, n10836, n10839, n10838, n10843, n10841, n10840,
    n10842, n10847, n10845, n10844, n10846, n10851, n10849, n10848, n10850,
    n10855, n10853, n10852, n10854, n10858, n11629, n10861, n10860, n10863,
    n10862, n12381, n10866, n10869, n10875, n10871, n10870, n10873, n10872,
    n10874, n10877, n10876, n10881, n10879, n10878, n10880, n10885, n10883,
    n10882, n10884, n10897, n12146, n12065, n10888, n10891, n10890, n10895,
    n10894, n10896, n10910, n10899, n12156, n10900, n12056, n11851, n10905,
    n10907, n10909, n10916, n10912, n10911, n10914, n10913, n10915, n10918,
    n10917, n10924, n10920, n10919, n10922, n10921, n10923, n10926, n10925,
    n10931, n10929, n10930, n10936, n10933, n11954, n11713, n10940, n10939,
    n10942, n10941, n10946, n10944, n10943, n10945, n10950, n10948, n10947,
    n10949, n10954, n10952, n10951, n10953, n10958, n10956, n10955, n10957,
    n10962, n10960, n10959, n10961, n10966, n10964, n10963, n10965, n10972,
    n10968, n10967, n10970, n10969, n10971, n10974, n10973, n10980, n10976,
    n10975, n10978, n10977, n10979, n10982, n10981, n10985, n10988, n10991,
    n10993, n10995, n11000, n10998, n10997, n11004, n11002, n11001, n11003,
    n11008, n11006, n11005, n11012, n11010, n11009, n11011, n11016, n11014,
    n11013, n11015, n11020, n11018, n11017, n11019, n11022, n11021, n11026,
    n11036, n11032, n11030, n11031, n11034, n11033, n11398, n11043, n11039,
    n11038, n11041, n11040, n11042, n11045, n11044, n11049, n11047, n11046,
    n11048, n11053, n11051, n11050, n11052, n11057, n11055, n11054, n11056,
    n11061, n11059, n11058, n11060, n11065, n11063, n11062, n11064, n11069,
    n11067, n11066, n11068, n11073, n11071, n11070, n11072, n11077, n11075,
    n11074, n11076, n11081, n11079, n11078, n11080, n11085, n11083, n11082,
    n11084, n11089, n11091, n11102, n11096, n11095, n11100, n11097, n11098,
    n11099, n11101, n11110, n11106, n11105, n11108, n11107, n11109, n11112,
    n11111, n11116, n11114, n11113, n11115, n11120, n11118, n11117, n11119,
    n11124, n11122, n11121, n11123, n11128, n11126, n11125, n11127, n11134,
    n11130, n11129, n11132, n11131, n11133, n11136, n11135, n11142, n11138,
    n11137, n11140, n11139, n11141, n11144, n11143, n11150, n11146, n11145,
    n11148, n11147, n11149, n11152, n11151, n11160, n11154, n11153, n11158,
    n11157, n11162, n11161, n11168, n11164, n11163, n11166, n11165, n11170,
    n11169, n11177, n11173, n11172, n11175, n11174, n11176, n11180, n11179,
    n11186, n11182, n11181, n11184, n11183, n11188, n11187, n11192, n11190,
    n11189, n11191, n11196, n11194, n11193, n11195, n11200, n11198, n11197,
    n11199, n11204, n11202, n11201, n11203, n11208, n11206, n11205, n11207,
    n11212, n11210, n11209, n11211, n11216, n11214, n11213, n11215, n11220,
    n11218, n11217, n11219, n11224, n11222, n11221, n11223, n11228, n11226,
    n11225, n11227, n11232, n11230, n11229, n11231, n11236, n11234, n11233,
    n11235, n11242, n11245, n11252, n11250, n11249, n11251, n11257, n11255,
    n11254, n11256, n11263, n11261, n11260, n11262, n11268, n11266, n11265,
    n11267, n11274, n11272, n11271, n11273, n11279, n11277, n11276, n11278,
    n11281, n11282, n11289, n11287, n11286, n11288, n11294, n11292, n11291,
    n11293, n11299, n11297, n11296, n11298, n11305, n11303, n11302, n11304,
    n11310, n11308, n11307, n11309, n11315, n11313, n11312, n11314, n11323,
    n13558, n11320, n11322, n11337, n11568, n11331, n11327, n11329, n11328,
    n11335, n11334, n11336, n11343, n11341, n11342, n11345, n12204, n11352,
    n11350, n11349, n11351, n11356, n11354, n11353, n11355, n11362, n11360,
    n11359, n11367, n11365, n11364, n11366, n11371, n11369, n11368, n11370,
    n11375, n11373, n11372, n11374, n11381, n11379, n11378, n11387, n11385,
    n11384, n11386, n11389, n11394, n11392, n11391, n11393, n11400, n11399,
    n11404, n13552, n11403, n11409, n11408, n11410, n11418, n11416, n11549,
    n11426, n11425, n11439, n11428, n11437, n11435, n11431, n11433, n11434,
    n11455, n11474, n11991, n11448, n11450, n11449, n11453, n11452, n11465,
    n11460, n11462, n11983, n11471, n11467, n11466, n11469, n11468, n11473,
    n11493, n11487, n11498, n11745, n11485, n11482, n11486, n11491, n11496,
    n11490, n11505, n11500, n11734, n11499, n11501, n11504, n11511, n11507,
    n11506, n11509, n11508, n11513, n11512, n11519, n11515, n11514, n11517,
    n11516, n11521, n11520, n11527, n11523, n11522, n11525, n11524, n11529,
    n11528, n11535, n11531, n11530, n11533, n11532, n11537, n11536, n11543,
    n11539, n11538, n11541, n11540, n11545, n11544, n11551, n11550, n11555,
    n13540, n11554, n11917, n11580, n11564, n11565, n11577, n11566, n11572,
    n11570, n11571, n11575, n11574, n11581, n11587, n11592, n11596, n11601,
    n11599, n11598, n11600, n11605, n11603, n11602, n11604, n11612, n11610,
    n11609, n11611, n11618, n11616, n11615, n11617, n11621, n11625, n11642,
    n11635, n11633, n11634, n11640, n11639, n11641, n11644, n11643, n11651,
    n11650, n11662, n11660, n11664, n11663, n11665, n11670, n11668, n11672,
    n11671, n11673, n11678, n11676, n11680, n11679, n11681, n11686, n11684,
    n11688, n11687, n11689, n11694, n11692, n11696, n11695, n11697, n11705,
    n11703, n11709, n11708, n11710, n11727, n11723, n11716, n11715, n11721,
    n11719, n11720, n11722, n11725, n11724, n11726, n11728, n11742, n11740,
    n11736, n11751, n11746, n11749, n11748, n11750, n11754, n11756, n11760,
    n11889, n11772, n11770, n11776, n11774, n11773, n11775, n11780, n11778,
    n11777, n11784, n11782, n11781, n11783, n11788, n11786, n11785, n11792,
    n11790, n11789, n11791, n11796, n11794, n11793, n11800, n11798, n11797,
    n11799, n11804, n11802, n11801, n11808, n11806, n11805, n11807, n11812,
    n11811, n11815, n11853, n11822, n11814, n11816, n11819, n11821, n11824,
    n11823, n11825, n11829, n11832, n11837, n11836, n11848, n11850, n11858,
    n11856, n11855, n11857, n11860, n11869, n11865, n11864, n11867, n11866,
    n11871, n11881, n11876, n11875, n11879, n11878, n11884, n13534, n11888,
    n11895, n11910, n11906, n11900, n11902, n11904, n11903, n11905, n11908,
    n11907, n11913, n11927, n11923, n11922, n11925, n11924, n11938, n11933,
    n11932, n11935, n11941, n11947, n11958, n11953, n11951, n11950, n11952,
    n11956, n11955, n11962, n11961, n11974, n11964, n11963, n11972, n11965,
    n11970, n11968, n11967, n12398, n11990, n11988, n11982, n11984, n12000,
    n11996, n11993, n11998, n11997, n11999, n12004, n12002, n12008, n12006,
    n12005, n12007, n12012, n12010, n12016, n12014, n12013, n12015, n12020,
    n12018, n12024, n12022, n12021, n12023, n12027, n12034, n12032, n12036,
    n12042, n12041, n12048, n12062, n12060, n12054, n12071, n12066, n12069,
    n12068, n12070, n12075, n12073, n12079, n12077, n12076, n12078, n12083,
    n12081, n12080, n12087, n12085, n12084, n12086, n12091, n12089, n12088,
    n12096, n12094, n12093, n12095, n12100, n12107, n12103, n12102, n12105,
    n12104, n12115, n12111, n12110, n12113, n12112, n12123, n12119, n12118,
    n12121, n12120, n12135, n12130, n12129, n12133, n12132, n12153, n12151,
    n12143, n12303, n12328, n12162, n12157, n12160, n12159, n12161, n12166,
    n12164, n12170, n12168, n12167, n12169, n12174, n12172, n12178, n12176,
    n12175, n12177, n12182, n12180, n12187, n12185, n12184, n12186, n12191,
    n12189, n12188, n12195, n12193, n12192, n12194, n12198, n12212, n12205,
    n13546, n12209, n12220, n12216, n12215, n12218, n12217, n12228, n12224,
    n12223, n12226, n12225, n12236, n12232, n12231, n12234, n12233, n12247,
    n12242, n12241, n12245, n12244, n12256, n12252, n12251, n12254, n12253,
    n12264, n12260, n12259, n12262, n12261, n12275, n12270, n12269, n12273,
    n12272, n12281, n12279, n12280, n12283, n12282, n12291, n12289, n12288,
    n12290, n12294, n12293, n12321, n12311, n12315, n12314, n12319, n12318,
    n12332, n12325, n12327, n12342, n12337, n12336, n12340, n12339, n12344,
    n12354, n12349, n12348, n12352, n12351, n12356, n12365, n12361, n12360,
    n12363, n12362, n12367, n12376, n12372, n12371, n12374, n12373, n12378,
    n12388, n12383, n12382, n12384, n12386, n12385, n12393, n12392, n12399,
    n12400, n12407, n12402, n12401, n12403, n12405, n12404, n12409, n12426,
    n12416, n12424, n12422, n12420, n12419, n12421, n12423, n12430, n12429,
    n12446, n12460, n12451, n12450, n12458, n12452, n12456, n12454, n12453,
    n12455, n12457, n12464, n12479, n12482, n12485, n12484, n12488, n12503,
    n12522, n12521, n12529, n12531, n12530, n12534, n12542, n12540, n12546,
    n12545, n12547, n12553, n12551, n12557, n12556, n12558, n12567, n12565,
    n12572, n12571, n12573, n12586, n12582, n12578, n12580, n12579, n12581,
    n12584, n12583, n12589, n12599, n12597, n12596, n12614, n12629, n12625,
    n12618, n12620, n12619, n12621, n12623, n12622, n12626, n12649, n12645,
    n12637, n12643, n12641, n12639, n12640, n12642, n12657, n12661, n12666,
    n12671, n12668, n12682, n12688, n12698, n12697, n12706, n12708, n12710,
    n12709, n12719, n12730, n12724, n12723, n12727, n12757, n12756, n12772,
    n12788, n12795, n12797, n12802, n12804, n12809, n12807, n12806, n12808,
    n12812, n12814, n12824, n12831, n12843, n12846, n12851, n12857, n12865,
    n12876, n12877, n12884, n12980, n12892, n12902, n12906, n12904, n12903,
    n12915, n12918, n12922, n12927, n12930, n12952, n13232, n12967, n12965,
    n12964, n12974, n12997, n13015, n13013, n13012, n13018, n13042, n13032,
    n13025, n13027, n13030, n13038, n13047, n13046, n13052, n13050, n13051,
    n13063, n13084, n13331, n13098, n13096, n13095, n13104, n13105, n13123,
    n13113, n13116, n13143, n13137, n13135, n13134, n13166, n13165, n13167,
    n13182, n13180, n13179, n13192, n13198, n13208, n13201, n13203, n13231,
    n13223, n13226, n13233, n13236, n13235, n13237, n13242, n13255, n13252,
    n13253, n13254, n13276, n13275, n13277, n13282, n13284, n13285, n13436,
    n13432, n13290, n13292, n13291, n13397, n13426, n13304, n13313, n13318,
    n13317, n13321, n13326, n13339, n13337, n13336, n13351, n13350, n13354,
    n13361, n13390, n13392, n13431, n13430, n13482, n13411, n13412, n13420,
    n13427, n13433, n13435, n13439, n13446, n13470, n13469, n13474, n13483,
    n13485, n13486, n13492, n13502, n13511, n13512, n13516, n13519, n13518,
    n13530, n13529, n13535, n13544, n13541, n13550, n13547, n13556, n13553,
    n13564, n13561, n13569, n13568;
  assign n13567 = ~n10242 | ~n10241;
  assign n13560 = ~n8805 | ~n12691;
  assign n13178 = ~n8497 | ~n12691;
  assign n13329 = n8965 | n10937;
  assign n10033 = ~n7391 & ~n7390;
  assign n9698 = ~STATEBS16_REG_SCAN_IN & ~STATE2_REG_2__SCAN_IN;
  assign n8091 = ~n8064 | ~n8063;
  assign n8045 = ~n8030;
  assign n10635 = ~n7955 | ~n7954;
  assign n10937 = ~n10574 | ~n10515;
  assign n8008 = ~n7613;
  assign n10515 = ~n7159 | ~n7158;
  assign n9653 = ~n8593;
  assign n7048 = ~n10340 & ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n7521 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n7637 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7631 = INSTQUEUERD_ADDR_REG_3__SCAN_IN & INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n8135 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n8111 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n10340 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n8593 = ~n10374 | ~n7521;
  assign n8062 = ~n8045 | ~n7965;
  assign n8118 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n8030 = ~n7956 | ~n10635;
  assign n8133 = ~n10319 | ~n10321;
  assign n12929 = ~n8955 | ~n8954;
  assign n10045 = ~n9723;
  assign n13316 = ~n13164 | ~n7669;
  assign n13490 = ~n9161 | ~n9160;
  assign n13045 = ~n9161 | ~n9117;
  assign n8806 = n13560 | n13389;
  assign n13463 = ~n13451;
  assign n13465 = ~n7664 | ~n12691;
  assign n13448 = ~n13447 & ~n13446;
  assign n13368 = ~n13367 & ~n13366;
  assign n13477 = ~n13476 & ~n13475;
  assign n13358 = ~n13488 | ~n13348;
  assign n13461 = ~n13460 | ~n13459;
  assign n13424 = ~n13423 & ~n13422;
  assign n9585 = ~n9584 | ~n9583;
  assign n13387 = ~n13386 & ~n13385;
  assign n13367 = ~n13364 | ~n13363;
  assign n9584 = ~n13312 | ~n9141;
  assign n13422 = ~n13421 | ~n13420;
  assign n13247 = ~n13362 | ~n13348;
  assign n13323 = ~n13312 | ~n13348;
  assign n13364 = ~n13362 | ~n9141;
  assign n13267 = ~n13266 & ~n13265;
  assign n13459 = ~n13458 & ~n13457;
  assign n13408 = ~n13407 & ~n13406;
  assign n13386 = ~n13383 | ~n13382;
  assign n13266 = ~n13263 | ~n13262;
  assign n13383 = ~n9141 | ~n13381;
  assign n13158 = ~n13381 | ~n13348;
  assign n13421 = ~n13418 & ~n13417;
  assign n13312 = n9580 ^ n9579;
  assign n13310 = ~n13309 & ~n13308;
  assign n9402 = ~n9401 | ~n9400;
  assign n13406 = ~n13454 & ~n13504;
  assign n13090 = ~n13261 | ~n13348;
  assign n13263 = ~n9141 | ~n13261;
  assign n9400 = ~n9399 & ~n9398;
  assign n13295 = ~n13294 | ~n13293;
  assign n13309 = ~n13307 | ~n13306;
  assign n13418 = ~n13416 & ~n13504;
  assign n13173 = ~n13170 & ~n13169;
  assign n13416 = n13220 ^ n13219;
  assign n9399 = ~n9388 | ~n13162;
  assign n13294 = ~n13305 | ~n13348;
  assign n13122 = ~n13121 & ~n13120;
  assign n13160 = ~n13159;
  assign n13145 = ~n13080 | ~n13079;
  assign n9574 = ~n13216;
  assign n13437 = n13436 & n13435;
  assign n13120 = ~n13119 | ~n13118;
  assign n13119 = ~n13117 & ~n13116;
  assign n13062 = ~n13061 & ~n13060;
  assign n9355 = ~n9347 | ~n9346;
  assign n13081 = ~n13077 | ~n13078;
  assign n13080 = ~n13077;
  assign n13117 = ~n13504 & ~n13115;
  assign n13061 = ~n13058 | ~n13057;
  assign n13010 = ~n13009 & ~n13008;
  assign n9346 = ~n9345 & ~n9344;
  assign n13344 = ~n13343 & ~n13342;
  assign n13009 = ~n13007 | ~n13006;
  assign n9345 = ~n9338 | ~n12866;
  assign n13296 = ~n13269 & ~n13451;
  assign n13142 = ~n13141 & ~n13140;
  assign n13342 = ~n13341 | ~n13340;
  assign n9569 = ~n12912;
  assign n13341 = ~n13331 | ~n13330;
  assign n9553 = ~n9552 | ~n9551;
  assign n13140 = ~n13139 | ~n13138;
  assign n13269 = ~n13331;
  assign n12983 = ~n12980 & ~n12979;
  assign n9167 = ~n9166 | ~n9165;
  assign n13462 = ~n13452 & ~n13451;
  assign n12862 = ~n9337 & ~n9336;
  assign n13041 = ~n13040 & ~n13039;
  assign n13139 = ~n13132 | ~n13330;
  assign n13074 = ~n13073 | ~n13072;
  assign n13214 = ~n13450 | ~n13330;
  assign n12958 = ~n12957 & ~n12956;
  assign n13248 = n13238 & n13237;
  assign n13452 = ~n13450;
  assign n9166 = ~n9155 & ~n9154;
  assign n9756 = ~n9755 | ~n9754;
  assign n12957 = ~n12953 | ~n12952;
  assign n13040 = ~n13034 | ~n13033;
  assign n9155 = ~n13504 & ~n12830;
  assign n12942 = ~n12941 & ~n12940;
  assign n9310 = ~n9306 | ~n9305;
  assign n9258 = ~n9254 | ~n9253;
  assign n12953 = ~n12950 & ~n12949;
  assign n9755 = ~n12881 | ~n13463;
  assign n12940 = ~n12939 | ~n12938;
  assign n13171 = n12902 & n12901;
  assign n12881 = ~n12945;
  assign n9206 = ~n9205 | ~n9204;
  assign n12939 = ~n12937 & ~n12936;
  assign n13357 = ~n13356 & ~n13355;
  assign n9087 = ~n9083 | ~n9082;
  assign n12849 = n12848 & n12847;
  assign n9327 = ~n9326 | ~n9325;
  assign n12847 = ~n12846 & ~n12845;
  assign n8485 = ~n8484 | ~n8483;
  assign n8996 = ~n8995 | ~n8994;
  assign n12873 = ~n13349;
  assign n9204 = ~n9203 & ~n9202;
  assign n13322 = ~n13321 & ~n13320;
  assign n13349 = ~n9301 | ~n9252;
  assign n9304 = ~n9301 | ~n9300;
  assign n9325 = ~n9324 & ~n9323;
  assign n8428 = ~n8427 | ~n8426;
  assign n13089 = ~n13088 & ~n13087;
  assign n8994 = ~n8993 & ~n8992;
  assign n9182 = ~n9181 | ~n9180;
  assign n12767 = ~n12766 & ~n12765;
  assign n8427 = n8425 & n8424;
  assign n13088 = ~n13085 | ~n13262;
  assign n13157 = ~n13156 & ~n13155;
  assign n12785 = ~n12782 & ~n12781;
  assign n9323 = ~n9322 | ~n9321;
  assign n12753 = ~n12752 & ~n12751;
  assign n12766 = ~n12763 | ~n12762;
  assign n8940 = ~n8936 | ~n8935;
  assign n9180 = ~n9179 & ~n9178;
  assign n8992 = ~n8991 | ~n8990;
  assign n8991 = ~n8987 & ~n8986;
  assign n12803 = ~n12801 & ~n12800;
  assign n8800 = ~n8795 | ~n8794;
  assign n9178 = ~n9177 | ~n9176;
  assign n13156 = ~n13153 | ~n13382;
  assign n9322 = ~n9320 & ~n9319;
  assign n8890 = ~n8809 | ~n8808;
  assign n12789 = ~n12787 & ~n12786;
  assign n12781 = ~n12780 | ~n12779;
  assign n12751 = ~n12750 | ~n12749;
  assign n9081 = ~n9078 | ~n9077;
  assign n13085 = ~n13084 & ~n13083;
  assign n13230 = ~n13229 & ~n13228;
  assign n12780 = ~n12778 & ~n12777;
  assign n12996 = ~n12995 & ~n12994;
  assign n13153 = ~n13152 & ~n13151;
  assign n12920 = ~n12919 & ~n12918;
  assign n9177 = ~n9175 & ~n9174;
  assign n12750 = ~n12748 & ~n12747;
  assign n12919 = ~n12916 | ~n13057;
  assign n12796 = ~n12794 & ~n12793;
  assign n12662 = ~n12660 & ~n12659;
  assign n12995 = ~n12992 | ~n12991;
  assign n12871 = ~n12870 & ~n12869;
  assign n12720 = ~n12716 & ~n12715;
  assign n12739 = ~n12738 & ~n12737;
  assign n12897 = ~n12896 & ~n12895;
  assign n13082 = ~n8977 | ~n8976;
  assign n12820 = ~n12816 & ~n12815;
  assign n12679 = ~n12675 & ~n12674;
  assign n12992 = n12990 & n12989;
  assign n12793 = ~n12792 | ~n12791;
  assign n12916 = n12915 & n12914;
  assign n12526 = ~n12518 & ~n12517;
  assign n12815 = ~n12814 | ~n12813;
  assign n12896 = ~n12893 | ~n13006;
  assign n12475 = ~n12472 & ~n12471;
  assign n12674 = ~n12673 | ~n12672;
  assign n12870 = ~n12867 | ~n12866;
  assign n12715 = ~n12714 | ~n12713;
  assign n12714 = ~n12704 & ~n12703;
  assign n12673 = ~n12665 & ~n12664;
  assign n12832 = ~n12829 & ~n12828;
  assign n12483 = ~n12481 & ~n12480;
  assign n12517 = ~n12516 | ~n12515;
  assign n13520 = ~n12988;
  assign n12471 = ~n12511 | ~n12470;
  assign n12489 = ~n12487 & ~n12486;
  assign n12867 = ~n12865 & ~n12864;
  assign n12445 = ~n12444 & ~n12443;
  assign n12893 = ~n12892 & ~n12891;
  assign n12506 = ~n12498 & ~n12497;
  assign n12535 = ~n12533 & ~n12532;
  assign n12829 = ~n12826 | ~n12825;
  assign n12497 = ~n12496 | ~n12495;
  assign n12443 = ~n12442 | ~n12441;
  assign n12049 = ~n12047 & ~n12046;
  assign n12615 = ~n12612 & ~n12611;
  assign n12442 = ~n12440 & ~n12439;
  assign n12101 = ~n12098 & ~n12097;
  assign n12496 = ~n12494 & ~n12493;
  assign n12825 = ~n12824 & ~n12823;
  assign n12044 = ~n12039 & ~n12038;
  assign n12700 = ~n12655 & ~n12654;
  assign n12655 = ~n12528 | ~n12527;
  assign n11597 = ~n11595 & ~n11594;
  assign n11844 = ~n11842 & ~n11841;
  assign n8486 = ~n12840 | ~n8476;
  assign n11768 = ~n11767 & ~n11766;
  assign n12469 = ~n8097 | ~n12435;
  assign n12611 = ~n12610 | ~n12609;
  assign n11757 = ~n11755 & ~n11754;
  assign n11945 = ~n11944 & ~n11943;
  assign n13213 = ~n13212 & ~n13211;
  assign n11766 = ~n11765 | ~n11764;
  assign n12822 = ~n12027 | ~n12477;
  assign n13194 = ~n13193 & ~n13192;
  assign n11841 = ~n11921 | ~n11840;
  assign n11588 = ~n11586 & ~n11585;
  assign n11622 = ~n11620 & ~n11619;
  assign n11943 = ~n11942 | ~n11941;
  assign n8476 = ~n8475 & ~n8474;
  assign n11978 = ~n11974 & ~n11973;
  assign n13407 = ~n13401 | ~n13456;
  assign n11765 = ~n11763 & ~n11762;
  assign n13212 = ~n13329 & ~n13196;
  assign n11423 = ~n11422 & ~n11421;
  assign n7662 = ~n7661 | ~n7660;
  assign n9736 = ~n9735 & ~n9734;
  assign n13193 = ~n13528 & ~n13196;
  assign n11563 = ~n11894 & ~n11556;
  assign n11899 = ~n11891 & ~n11890;
  assign n7660 = ~n7659 & ~n7658;
  assign n9735 = ~n13329 & ~n13440;
  assign n11556 = ~n11555 | ~n11554;
  assign n12026 = n8500 & n8499;
  assign n12689 = ~n12688 | ~n12687;
  assign n11421 = ~n11420 | ~n11419;
  assign n11973 = ~n11972 | ~n11971;
  assign n11283 = ~n11281 & ~n11280;
  assign n7661 = ~n7649 | ~STATE2_REG_0__SCAN_IN;
  assign n11246 = ~n11244 & ~n11243;
  assign n13211 = ~n13210 | ~n13209;
  assign n11348 = ~n11347 & ~n11346;
  assign n12508 = ~n12683 | ~STATE2_REG_3__SCAN_IN;
  assign n12687 = ~n12686 | ~STATE2_REG_1__SCAN_IN;
  assign n11420 = ~n11418 & ~n11417;
  assign n7659 = ~n7654 & ~n7653;
  assign n11885 = ~n11761 | ~n11760;
  assign n13209 = ~n13208 & ~n13207;
  assign n8433 = ~n8431 | ~n8430;
  assign n13107 = ~n13106 & ~n13105;
  assign n9731 = ~n9727 & ~n13189;
  assign n12683 = ~n12685 | ~STATE2_REG_0__SCAN_IN;
  assign n9768 = ~n9767 | ~n9766;
  assign n12413 = ~n12412 & ~n12411;
  assign n11346 = ~n11345 | ~n11344;
  assign n8431 = ~n11241 | ~n7016;
  assign n11916 = ~n11910 & ~n11909;
  assign n8417 = ~n11241;
  assign n10992 = ~n10990 & ~n10989;
  assign n11548 = ~n11416 | ~n11415;
  assign n13072 = ~n13071 & ~n13070;
  assign n11037 = ~n11036 & ~n11035;
  assign n12633 = ~n12629 & ~n12628;
  assign n10996 = ~n10994 & ~n10993;
  assign n9767 = ~n13507 | ~n9765;
  assign n11412 = ~n12200 & ~n11405;
  assign n12213 = ~n12212 & ~n12211;
  assign n13020 = ~n13019 & ~n13018;
  assign n13207 = ~n13206 | ~n13205;
  assign n12976 = ~n12975 & ~n12974;
  assign n13205 = n13204 & n13203;
  assign n12628 = ~n12627 | ~n12626;
  assign n9739 = ~n9597 & ~n9596;
  assign n12396 = ~n12395 & ~n12394;
  assign n13070 = ~n13069 | ~n13068;
  assign n9727 = ~n13103 & ~n13190;
  assign n11035 = ~n11034 | ~n11033;
  assign n13068 = ~n13067 & ~n13066;
  assign n9597 = ~n13202 & ~n9883;
  assign n13033 = ~n13032 & ~n13031;
  assign n9596 = ~n9595 & ~REIP_REG_31__SCAN_IN;
  assign n12199 = ~n11341 | ~n11340;
  assign n13345 = ~n13327 | ~n13326;
  assign n13280 = ~n13279 & ~n13278;
  assign n12461 = ~n12460 & ~n12459;
  assign n10831 = ~n10829 & ~n10828;
  assign n12434 = ~n10985 | ~n11024;
  assign n12653 = ~n12649 & ~n12648;
  assign n12432 = ~n12426 & ~n12425;
  assign n10672 = ~n10670 & ~n10669;
  assign n12627 = ~n12625 & ~n12624;
  assign n13188 = ~n13187 & ~n13186;
  assign n13031 = ~n13030 | ~n13029;
  assign n13066 = ~n13065 | ~n13064;
  assign n9385 = n13271 & n9384;
  assign n11698 = ~n11694 & ~n11693;
  assign n11682 = ~n11678 & ~n11677;
  assign n9764 = ~n12973 | ~n9763;
  assign n13202 = ~n13324 | ~n9590;
  assign n13327 = ~n13324 | ~REIP_REG_29__SCAN_IN;
  assign n12574 = ~n12567 & ~n12566;
  assign n12548 = ~n12542 & ~n12541;
  assign n13129 = ~n13128 & ~REIP_REG_28__SCAN_IN;
  assign n11666 = ~n11662 & ~n11661;
  assign n7646 = ~n7645 | ~n7644;
  assign n13102 = ~n13187;
  assign n12559 = ~n12553 & ~n12552;
  assign n9595 = n13325 & n9594;
  assign n11690 = ~n11686 & ~n11685;
  assign n12648 = ~n12647 | ~n12646;
  assign n11711 = ~n11705 & ~n11704;
  assign n11674 = ~n11670 & ~n11669;
  assign n11024 = ~n10984 | ~n10983;
  assign n12109 = ~n12107 & ~n12106;
  assign n7645 = ~n7643 | ~n7642;
  assign n12230 = ~n12228 & ~n12227;
  assign n12250 = ~n12247 & ~n12246;
  assign n12222 = ~n12220 & ~n12219;
  assign n12138 = ~n12135 & ~n12134;
  assign n13539 = ~n10668 | ~n10667;
  assign n12266 = ~n12264 & ~n12263;
  assign n12238 = ~n12236 & ~n12235;
  assign n13039 = ~n13038 | ~n13037;
  assign n12125 = ~n12123 & ~n12122;
  assign n12956 = ~n12955 & ~n12954;
  assign n11438 = ~n11437 & ~n11436;
  assign n10571 = ~n10569 & ~n10568;
  assign n13271 = ~n9575 & ~n9577;
  assign n12258 = ~n12256 & ~n12255;
  assign n12647 = ~n12645 & ~n12644;
  assign n13325 = ~n13127 & ~n9593;
  assign n11817 = ~n11861 | ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n13324 = ~n9589 & ~n13125;
  assign n11834 = ~n11861 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n12924 = ~n12923 & ~n12922;
  assign n13533 = ~n10827 | ~n10826;
  assign n12278 = ~n12275 & ~n12274;
  assign n12117 = ~n12115 & ~n12114;
  assign n11826 = ~n11861 | ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n13128 = ~n13127 & ~n13126;
  assign n13130 = ~n13125 & ~n13124;
  assign n9583 = ~n9582 & ~n9581;
  assign n13510 = ~n13509 | ~n13508;
  assign n13125 = ~n9588 | ~n13036;
  assign n11861 = ~n11859;
  assign n9575 = ~n13215 | ~n13218;
  assign n13494 = ~n13493 & ~n13492;
  assign n12879 = ~n12878 & ~n12877;
  assign n8997 = ~n9313 & ~REIP_REG_20__SCAN_IN;
  assign n12886 = n12885 & n12884;
  assign n9183 = ~n9313 & ~n9170;
  assign n9328 = ~n9313 & ~n9312;
  assign n11414 = ~n8077 & ~n8076;
  assign n12861 = ~n12858 & ~n12857;
  assign n12943 = ~n12933 | ~n12932;
  assign n12737 = ~n12736 | ~n12735;
  assign n12955 = n13036 & REIP_REG_25__SCAN_IN;
  assign n12563 = ~n12330 | ~n12329;
  assign n11839 = ~n8094 & ~n8093;
  assign n13545 = ~n10462 | ~n10666;
  assign n11930 = ~n11927 & ~n11926;
  assign n13444 = ~n13468 | ~n13443;
  assign n12933 = ~n12928 | ~n12927;
  assign n13215 = ~n9383 & ~n13146;
  assign n13036 = ~n12926 | ~n9591;
  assign n12736 = ~n12732 | ~REIP_REG_17__SCAN_IN;
  assign n13551 = ~n10353 | ~n10352;
  assign n12609 = ~n12608 | ~n12607;
  assign n12211 = ~n12210 | ~n12209;
  assign n11701 = ~n11463 | ~n11983;
  assign n7636 = ~INSTQUEUEWR_ADDR_REG_4__SCAN_IN & ~n7588;
  assign n8076 = ~n8075 & ~INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n11758 = ~n8087 & ~n8088;
  assign n12740 = ~n12730 & ~n12729;
  assign n13148 = ~n13147 & ~n13146;
  assign n9374 = ~n12910 & ~n9748;
  assign n12329 = ~n12328 & ~n12327;
  assign n8055 = ~n8054;
  assign n9382 = ~n13147 & ~n9381;
  assign n12248 = ~n12058 | ~n12057;
  assign n12210 = ~n12206 & ~n12205;
  assign n13078 = ~n13076 | ~n13144;
  assign n9573 = ~n13147 & ~n9572;
  assign n12979 = ~n12978;
  assign n7588 = ~n7587 | ~n7586;
  assign n9330 = ~n9329;
  assign n9579 = ~n9578 & ~n9577;
  assign n8053 = ~n8052 & ~INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n13243 = ~n13242 & ~n13241;
  assign n9414 = ~n9413 & ~n9412;
  assign n9749 = ~n9748 & ~n9747;
  assign n11613 = ~n11485 & ~n11484;
  assign n12136 = ~n12330 | ~n11986;
  assign n12744 = ~n9147 | ~INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n13449 = ~n13428 | ~n13427;
  assign n11882 = ~n11738 | ~n11737;
  assign n12467 = ~n9147 | ~INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n12595 = ~n12592 & ~n12591;
  assign n9568 = ~n12910;
  assign n13346 = ~n9744 & ~n9743;
  assign n12435 = ~n9147 | ~INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n13443 = ~INSTADDRPOINTER_REG_30__SCAN_IN | ~n13442;
  assign n8088 = ~n8086 & ~n11893;
  assign n12729 = ~n12728 | ~n12727;
  assign n11339 = ~n8056 & ~n7973;
  assign n13409 = ~n13428 | ~n13399;
  assign n11463 = ~n12147 & ~n11462;
  assign n13311 = ~n13304 | ~n13303;
  assign n13489 = ~n12876 | ~n12883;
  assign n12276 = ~n12149 | ~n12148;
  assign n9148 = ~n9147 & ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n8077 = ~n8074 & ~n9088;
  assign n9387 = ~n9404 & ~n9407;
  assign n9586 = ~n9564 & ~n9563;
  assign n11626 = ~n11625 | ~n11624;
  assign n12986 = ~n12985 | ~n12984;
  assign n13268 = ~n13260 | ~n13259;
  assign n13011 = ~n13004 | ~n13003;
  assign n10665 = ~n8183 & ~n8182;
  assign n12240 = ~n12067 & ~n12066;
  assign n8479 = ~n9146 | ~n12835;
  assign n12058 = ~n12055 & ~n12054;
  assign n9168 = ~n9130 & ~n9129;
  assign n9570 = ~n12909;
  assign n11738 = ~n11735 & ~n11734;
  assign n13425 = ~n13413 | ~n13412;
  assign n9563 = ~n9562 & ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n9744 = ~n9745;
  assign n10908 = ~n12056 & ~n10907;
  assign n11986 = ~n11985 & ~n11984;
  assign n9748 = ~n13288 & ~INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n13218 = ~n13288 | ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n13513 = ~n13503 | ~n13502;
  assign n9404 = ~n13288 & ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n9384 = ~n9743 & ~n9747;
  assign n11624 = ~n11623 | ~n7597;
  assign n12568 = ~n12311 & ~n12310;
  assign n7586 = ~n7585 | ~n7584;
  assign n13388 = ~n13380 | ~n13379;
  assign n13369 = ~n13361 | ~n13360;
  assign n13147 = ~n13288 & ~INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n13076 = ~n13288 | ~INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n9411 = ~n13241;
  assign n12206 = ~n12203 & ~n12202;
  assign n13303 = ~n13302 | ~n13432;
  assign n7973 = ~n7972 & ~INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n13399 = ~n13441 | ~n13431;
  assign n8074 = ~n8073 & ~n8072;
  assign n13428 = ~n13396 | ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n8087 = ~n8085 & ~INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n13442 = ~INSTADDRPOINTER_REG_31__SCAN_IN & ~n13441;
  assign n9147 = ~n9146;
  assign n12888 = ~n13288 | ~INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n12931 = ~n9956 & ~n9185;
  assign n12591 = ~n12590 | ~n12589;
  assign n12855 = ~n12852 & ~n12851;
  assign n11658 = ~n11653 & ~n11652;
  assign n12149 = ~n12144 & ~n12143;
  assign n12728 = ~n12726 & ~n12725;
  assign n11503 = ~n11502 & ~n11501;
  assign n11484 = ~n11483 & ~n11494;
  assign n12038 = ~n12037 | ~n12036;
  assign n11915 = ~n11914 & ~n11913;
  assign n11946 = ~n11938 & ~n11937;
  assign n9181 = ~n9314 | ~REIP_REG_21__SCAN_IN;
  assign n11977 = ~REIP_REG_11__SCAN_IN | ~n11976;
  assign n12606 = ~REIP_REG_14__SCAN_IN & ~n12605;
  assign n9326 = ~n9314 | ~REIP_REG_22__SCAN_IN;
  assign n12412 = ~n12408 & ~REIP_REG_11__SCAN_IN;
  assign n12768 = ~n12760 | ~n12759;
  assign n12203 = ~n12201 & ~n12200;
  assign n11995 = ~n11994 & ~n11993;
  assign n9577 = ~n13434 & ~n13480;
  assign n12037 = ~n12726 & ~n12035;
  assign n9403 = ~n13500 & ~n13274;
  assign n11747 = ~n11744 & ~n11743;
  assign n13413 = ~n13487;
  assign n12504 = ~n12500 & ~n12499;
  assign n12592 = ~n12635 & ~n13557;
  assign n9144 = ~n13434 | ~n8481;
  assign n11914 = ~n11912 & ~REIP_REG_10__SCAN_IN;
  assign n11447 = ~n11459 & ~n11457;
  assign n11985 = ~n11994 & ~n11992;
  assign n12590 = ~n12586 & ~n12585;
  assign n9771 = ~n13398 | ~n9759;
  assign n13441 = ~n13398 | ~n13397;
  assign n9314 = ~n9184 & ~n12721;
  assign n12816 = ~n12812 | ~n12811;
  assign n12850 = ~n12834 | ~INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n12158 = ~n12155 & ~n12154;
  assign n13396 = ~n13300 | ~n13426;
  assign n12848 = ~n12839 | ~INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n13384 = ~n8888 | ~n8887;
  assign n12395 = ~n12389 & ~REIP_REG_9__SCAN_IN;
  assign n10632 = ~n10630 & ~n10797;
  assign n7585 = ~n7583 & ~n7582;
  assign n8085 = ~n8084 | ~n13434;
  assign n11735 = ~n11744 & ~n11733;
  assign n12778 = ~n12775 & ~n12774;
  assign n13144 = ~n13434 | ~n13257;
  assign n11583 = ~n11577 & ~n11576;
  assign n9333 = ~n13434 | ~n9375;
  assign n13288 = ~n13434;
  assign n12310 = ~n12323 & ~n12309;
  assign n12055 = ~n12064 & ~n12053;
  assign n13497 = ~n13487 & ~n13486;
  assign n11937 = ~n11936 | ~n11935;
  assign n12326 = ~n12323 & ~n12322;
  assign n11502 = n11495 & n11494;
  assign n9146 = ~n7007 | ~n8092;
  assign n10330 = ~n10326 & ~n10325;
  assign n11976 = ~REIP_REG_12__SCAN_IN & ~n12408;
  assign n12144 = ~n12155 & ~n12142;
  assign n11461 = ~n11459 & ~n11458;
  assign n9562 = ~n13487 & ~n13410;
  assign n8056 = ~n7971 & ~n12202;
  assign n9130 = ~n9122 & ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n12981 = ~n13434 | ~n13002;
  assign n11171 = ~n10889 & ~n10888;
  assign n12067 = ~n12064 & ~n12063;
  assign n12909 = ~n13434 & ~n13053;
  assign n9347 = ~n13000 | ~INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n8165 = ~n8158 & ~n8174;
  assign n12414 = ~n12407 & ~n12406;
  assign n9564 = ~n13479 & ~n13480;
  assign n11971 = ~n11970 & ~n11969;
  assign n11936 = ~n12726 & ~n11934;
  assign n12499 = ~n11920 | ~n11919;
  assign n10889 = ~n10904 & ~n7012;
  assign n12155 = ~n12141 | ~n12305;
  assign n12064 = ~n12052 | ~n12305;
  assign n12431 = ~n12430 & ~n12429;
  assign n7007 = n8091 & n8067;
  assign n12323 = ~n12306 | ~n12305;
  assign n13557 = ~n10307 | ~n10306;
  assign n11495 = ~n11480 & ~n11479;
  assign n12604 = ~n8959 | ~n12631;
  assign n7582 = ~n7581 & ~n7580;
  assign n7971 = ~n7970 & ~n7969;
  assign n12775 = ~n12773 | ~n12772;
  assign n7640 = ~n7638 & ~n7637;
  assign n9354 = ~n12833 & ~n9353;
  assign n10800 = ~n10798 & ~n10797;
  assign n13300 = ~n13359 | ~n13397;
  assign n12834 = ~INSTADDRPOINTER_REG_14__SCAN_IN & ~n12833;
  assign n10630 = ~n10629 & ~n10628;
  assign n10510 = ~n10508 & ~n10797;
  assign n12839 = ~n12838 | ~n12837;
  assign n7635 = ~n7634 | ~n7638;
  assign n9184 = ~n9171 & ~n9311;
  assign n11253 = ~n10495 & ~n10494;
  assign n10602 = ~n10600 & ~n10797;
  assign n10906 = ~n10904 & ~n10903;
  assign n11264 = ~n10547 & ~n10546;
  assign n11300 = ~n10620 & ~n10619;
  assign n11459 = ~n11446 & ~n11445;
  assign n12300 = ~n12296 & ~n12295;
  assign n12397 = ~n12388 & ~n12387;
  assign n9781 = ~n13359 & ~n9780;
  assign n11744 = ~n11732 | ~n12305;
  assign n12713 = ~n12712 & ~n12711;
  assign n11311 = ~n10589 & ~n10588;
  assign n10560 = ~n10558 & ~n10797;
  assign n13110 = ~n13001 & ~n13000;
  assign n12408 = ~n12398 | ~n12631;
  assign n11382 = n10680 & n10679;
  assign n12493 = ~n12501 & ~n12492;
  assign n13500 = ~n9365 & ~n9364;
  assign n12672 = ~n12671 & ~n12670;
  assign n12200 = n12196 & n12197;
  assign n9129 = ~n13000 & ~n9349;
  assign n11994 = ~n11981 | ~n12305;
  assign n11363 = ~n10786 & ~n10785;
  assign n13249 = ~n13052 | ~n13051;
  assign n10508 = ~n10506 & ~n10505;
  assign n10495 = ~n10504 & ~n10506;
  assign n12141 = ~n12140 | ~STATEBS16_REG_SCAN_IN;
  assign n10547 = ~n10555 & ~n10557;
  assign n9365 = ~n9362 | ~n9557;
  assign n11732 = ~n11731 | ~STATEBS16_REG_SCAN_IN;
  assign n11446 = ~n11444 & ~n11443;
  assign n8037 = ~n8036 & ~INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n13479 = ~n9557 | ~n9556;
  assign n13359 = n9779 & n9778;
  assign n10558 = ~n10557 & ~n10556;
  assign n11479 = ~n11478 & ~n11477;
  assign n12833 = ~n12836;
  assign n11981 = ~n11980 | ~STATEBS16_REG_SCAN_IN;
  assign n12773 = ~n12514 & ~n12513;
  assign n11959 = ~n11958 & ~n11957;
  assign n11894 = ~INSTADDRPOINTER_REG_7__SCAN_IN & ~n12514;
  assign n12306 = ~n12304 | ~STATEBS16_REG_SCAN_IN;
  assign n7638 = n7633 & n7632;
  assign n8173 = ~n8166 | ~n9633;
  assign n12052 = ~n12051 | ~STATEBS16_REG_SCAN_IN;
  assign n12492 = ~n11918 & ~n11917;
  assign n10904 = ~n10887 & ~n11830;
  assign n7969 = n8166 & n8092;
  assign n10786 = ~n10794 & ~n10796;
  assign n13000 = ~n9128 | ~n12524;
  assign n12197 = ~n11430 & ~n11432;
  assign n7634 = n7626 & n7625;
  assign n12783 = ~n12524 | ~n12523;
  assign n12201 = ~n12524 | ~n11410;
  assign n10600 = ~n10599 & ~n10598;
  assign n13423 = ~n13415 & ~n13414;
  assign n10798 = ~n10796 & ~n10795;
  assign n10557 = ~n10545 & ~n11445;
  assign n9779 = ~n13377 & ~n9775;
  assign n11290 = ~n10525 & ~n10524;
  assign n12304 = ~n12561 | ~n12537;
  assign n7633 = ~n7629 | ~n7628;
  assign n11430 = ~n11317 & ~n11316;
  assign n12514 = ~n11547 & ~n11546;
  assign n10506 = ~n10493 & ~n11445;
  assign n10654 = ~n10652 & ~n10797;
  assign n13524 = ~n13523 | ~n13522;
  assign n11383 = ~n10901;
  assign n11275 = ~n10641 & ~n10640;
  assign n10887 = ~n10614 & ~n11480;
  assign n11614 = ~n11475;
  assign n12722 = ~n12705 & ~n8961;
  assign n7626 = ~n7639 & ~n7610;
  assign n12523 = ~n12522 & ~n12521;
  assign n11731 = ~n11874 | ~n11872;
  assign n9557 = ~n9361 & ~n13377;
  assign n12140 = ~n12267 | ~n12183;
  assign n8026 = ~n8025;
  assign n9128 = ~n9124 & ~n9123;
  assign n11980 = ~n12126 | ~n12128;
  assign n8027 = ~n8025 & ~INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n12051 = ~n12239 | ~n12092;
  assign n10796 = ~n10783 & ~n11445;
  assign n10538 = ~n10536 & ~n10797;
  assign n10312 = ~n8157 | ~n8156;
  assign n11427 = ~n11331 & ~n11330;
  assign n10692 = ~n10676 & ~n11480;
  assign n12837 = ~n12758 & ~n13377;
  assign n13415 = ~n13378 & ~n13377;
  assign n10536 = ~n10535 & ~n10534;
  assign n10614 = ~n10621 & ~n11478;
  assign n13378 = ~n13376 | ~n13375;
  assign n9364 = ~n9363 & ~n13484;
  assign n13531 = ~n13530 | ~n13529;
  assign n10583 = ~n10590 | ~STATEBS16_REG_SCAN_IN;
  assign n13001 = ~n12999 & ~n12998;
  assign n9369 = ~n9366 & ~n11579;
  assign n9560 = ~n11579 & ~n9558;
  assign n9121 = ~n12754 & ~n11579;
  assign n11606 = ~n11476;
  assign n11918 = ~n11920 & ~n12999;
  assign n10525 = ~n10533 & ~n10535;
  assign n9124 = ~n13049 & ~n9357;
  assign n12612 = ~n12600 | ~n12805;
  assign n11475 = ~n10681 & ~n10674;
  assign n12043 = ~n12042 & ~n12041;
  assign n12128 = ~n10548 | ~n10886;
  assign n7629 = n7627 & n11813;
  assign n10652 = ~n10651 & ~n10650;
  assign n10396 = ~n10395;
  assign n7639 = ~n7600 | ~n7599;
  assign n13563 = ~n13562 | ~n13561;
  assign n11476 = ~n11847 & ~n10886;
  assign n13555 = ~n13554 | ~n13553;
  assign n13549 = ~n13548 | ~n13547;
  assign n12593 = ~n12285 | ~n11656;
  assign n10395 = ~n10335 | ~n10334;
  assign n10496 = ~n10541 & ~n11810;
  assign n12999 = ~n13374 & ~n13371;
  assign n7628 = ~n7556 & ~n7555;
  assign n11443 = ~n11442 & ~n11830;
  assign n12028 = ~n11931 & ~n8960;
  assign n12600 = ~n12599 & ~n12598;
  assign n10651 = ~n11445 & ~n11442;
  assign n13049 = ~n13371;
  assign n10304 = ~n8144 & ~n8143;
  assign n9127 = ~n9126 | ~n8001;
  assign n9589 = ~REIP_REG_28__SCAN_IN & ~n12721;
  assign n10535 = ~n10523 & ~n11445;
  assign n12944 = ~n13329;
  assign n9368 = ~n13045 & ~n9772;
  assign n7984 = ~n7983 & ~INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n13299 = ~n11324 | ~n13045;
  assign n12721 = ~n12926;
  assign n10794 = ~n10782 & ~n11357;
  assign n9205 = ~n9191 & ~n9190;
  assign n12635 = ~n12298;
  assign n11546 = ~n13045 & ~n11558;
  assign n9120 = ~n13045 & ~n12755;
  assign n13251 = ~n13045 & ~n9559;
  assign n7556 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~n10331;
  assign n7595 = ~n7594 | ~n7593;
  assign n7538 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~n10331;
  assign n12577 = ~n11655 | ~REIP_REG_1__SCAN_IN;
  assign n10597 = ~n10585 & ~n10587;
  assign n13138 = ~n13137 & ~n13136;
  assign n13507 = ~n13490;
  assign n12285 = ~n11714 & ~n11718;
  assign n8144 = ~n11852 & ~n8174;
  assign n13504 = ~n9141;
  assign n11442 = ~n10642 & ~n11480;
  assign n10533 = ~n11284 & ~n10522;
  assign n13340 = ~n13339 & ~n13338;
  assign n8132 = ~n8129;
  assign n12617 = ~n12418 & ~n12417;
  assign n11712 = ~n10235 | ~n10321;
  assign n10649 = ~n11269 & ~n10639;
  assign n12949 = ~n12948 | ~n12947;
  assign n12936 = ~n12935 | ~n12934;
  assign n9319 = ~n9318 | ~n9317;
  assign n7537 = ~n7592 & ~n10362;
  assign n12298 = ~n12946 | ~n11648;
  assign n10331 = ~n7592;
  assign n13559 = ~n13528;
  assign n11655 = ~n12929;
  assign n13185 = ~n8806;
  assign n12154 = ~n12142;
  assign n13229 = ~n13226 | ~n13225;
  assign n12968 = ~n12967 & ~n12966;
  assign n10694 = ~n10689 & ~n10797;
  assign n13169 = ~n13168 | ~n13167;
  assign n10581 = ~n11820 | ~n10635;
  assign n9551 = ~n9550 & ~n9549;
  assign n9161 = ~n9125;
  assign n13355 = ~n13354 | ~n13353;
  assign n10673 = ~n11820 & ~n7990;
  assign n10613 = ~n11820 & ~n11810;
  assign n13099 = ~n13098 & ~n13097;
  assign n13016 = ~n13015 & ~n13014;
  assign n12057 = ~n12056 & ~n12147;
  assign n12063 = ~n12053;
  assign n11743 = ~n11733;
  assign n12472 = ~n12465 | ~n12464;
  assign n12764 = ~n11593 | ~n11592;
  assign n10555 = ~n10544 & ~n11258;
  assign n13183 = ~n13182 & ~n13181;
  assign n11737 = ~n12147 & ~n11736;
  assign n13333 = ~n13197;
  assign n13475 = ~n13474 | ~n13473;
  assign n12907 = ~n12906 & ~n12905;
  assign n8965 = ~EBX_REG_31__SCAN_IN | ~n8964;
  assign n9754 = ~n9753 & ~n9752;
  assign n10504 = ~n11247 & ~n10492;
  assign n13293 = ~n13292 & ~n13291;
  assign n12946 = ~n13330;
  assign n12148 = ~n12328 & ~n12147;
  assign n10797 = ~n11456 | ~n10507;
  assign n11155 = ~n10747;
  assign n11494 = ~n11482 | ~n12307;
  assign n8954 = ~n8980 & ~n11636;
  assign n13334 = ~n13199;
  assign n12053 = ~n10586 & ~n12307;
  assign n10928 = ~n13560;
  assign n12801 = ~n12798 | ~n12797;
  assign n10492 = ~n10542 & ~n12307;
  assign n13176 = ~n12799;
  assign n12636 = ~n11714 & ~n8957;
  assign n11733 = ~n10586 & ~n7936;
  assign n12543 = ~n11456 | ~DATAI_5_;
  assign n10449 = ~n10456 & ~n10447;
  assign n10444 = ~n10451 & ~n10442;
  assign n10403 = ~n10401 & ~n10400;
  assign n10458 = ~n10456 & ~n10455;
  assign n10419 = ~n10417 & ~n10416;
  assign n10436 = ~n10434 & ~n10433;
  assign n12147 = ~n11456 | ~n12302;
  assign n10427 = ~n10425 & ~n10424;
  assign n10415 = ~n10413 & ~n10412;
  assign n10411 = ~n10409 & ~n10408;
  assign n12142 = ~n10781 & ~n12307;
  assign n10431 = ~n10429 & ~n10428;
  assign n10440 = ~n10438 & ~n10437;
  assign n8964 = ~n8963 & ~n11636;
  assign n10453 = ~n10451 & ~n10450;
  assign n12338 = n10515 & n10747;
  assign n10407 = ~n10405 & ~n10404;
  assign n10423 = ~n10421 & ~n10420;
  assign n9163 = ~n11589 | ~n11584;
  assign n13571 = ~n13565 & ~n8533;
  assign n8128 = ~n10215;
  assign n10781 = ~n11854 | ~n12287;
  assign n11810 = ~n7990;
  assign n11636 = ~STATE2_REG_2__SCAN_IN | ~n11632;
  assign n10169 = ~n10080;
  assign n11456 = ~n11627;
  assign n7423 = ~n7410 & ~READY_N;
  assign n10677 = ~n11481 & ~n11828;
  assign n12322 = ~n12308 & ~n12307;
  assign n11992 = ~n12308 & ~n7936;
  assign n11714 = ~n11632;
  assign n12805 = ~n11632 | ~n11631;
  assign n13472 = ~n13316;
  assign n13199 = ~n11632 | ~STATE2_REG_3__SCAN_IN;
  assign n10456 = ~n10446 & ~n10445;
  assign n11591 = ~n11238 | ~n11237;
  assign n12308 = ~n11854 | ~n10616;
  assign n11627 = ~n10491 | ~n10490;
  assign n9541 = ~n9540 | ~n9539;
  assign n13391 = ~n13178;
  assign n13467 = ~n13164;
  assign n13565 = ~n7005;
  assign n10451 = n13566 & DATAI_14_;
  assign n10080 = ~n10078 | ~n10076;
  assign n10079 = ~n10078 | ~n10077;
  assign n7410 = ~n7409 & ~n8944;
  assign n7536 = ~n11854 & ~n7561;
  assign n12490 = ~n10988 | ~n11087;
  assign n9539 = ~n9538 & ~n9537;
  assign n9705 = ~n13332 & ~n9789;
  assign n8972 = ~n9598 | ~PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n13348 = ~n13465;
  assign n10674 = ~n10886;
  assign n9598 = ~n9704 & ~n8971;
  assign n7935 = ~n7988;
  assign n7590 = ~n7539 | ~n7540;
  assign n7650 = ~n10033;
  assign n8951 = ~n10033 | ~n8945;
  assign n7988 = ~n7995 | ~n8090;
  assign n12307 = ~n7936;
  assign n7664 = ~n10033 & ~n9134;
  assign n9497 = ~n13234 & ~n9789;
  assign n10242 = ~n10033 & ~n10032;
  assign n9100 = ~n10033 & ~n7641;
  assign n8496 = ~n7392 & ~n10033;
  assign n9456 = ~n13161 & ~n9789;
  assign n7995 = ~n7927 | ~n7991;
  assign n9536 = ~n9496 & ~n9490;
  assign n9302 = ~n9299 & ~n9298;
  assign n10865 = ~n11887 | ~n11886;
  assign n7560 = ~n7558 | ~n7557;
  assign n9075 = ~n9074 & ~n9073;
  assign n9496 = ~n9416 | ~PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n9298 = ~n12951 & ~n9789;
  assign n10211 = ~n8123 | ~n8122;
  assign n9251 = ~n9249 & ~n9248;
  assign n8123 = ~n11949 | ~n9633;
  assign n9249 = ~n13352 & ~n9789;
  assign n9073 = ~n9072 | ~n9071;
  assign n9416 = ~n9297 & ~n8970;
  assign n8933 = ~n8932;
  assign n7485 = ~n7489;
  assign n9297 = ~n9208 | ~PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n7540 = ~n7494 | ~n7493;
  assign n7378 = ~n7377 | ~n7376;
  assign n9208 = ~n9070 & ~n8969;
  assign n7488 = ~n7487;
  assign n9070 = ~n8968 | ~PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n10857 = ~n11319 & ~n11318;
  assign n8974 = ~n8750 | ~n8749;
  assign n12476 = ~n8583 | ~n8582;
  assign n9103 = ~n9102 & ~n9101;
  assign n7421 = ~n9099 & ~n7420;
  assign n8930 = ~n8929 | ~n8928;
  assign n8749 = ~n8748 | ~n8747;
  assign n8707 = ~n8706 | ~n8705;
  assign n8789 = ~n8788 | ~n8787;
  assign n8944 = ~n7602 & ~n7516;
  assign n7561 = ~n9114 & ~n7517;
  assign n8968 = ~n8892 & ~n8891;
  assign n12527 = ~n8630 | ~n8629;
  assign n8668 = ~n8667 & ~n8666;
  assign n9498 = ~n9495 & ~n9494;
  assign n7370 = ~n7369 & ~n7368;
  assign n8892 = ~n8751 | ~PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n9299 = ~n9296 & ~n9295;
  assign n9248 = ~n9247 | ~n9246;
  assign n9455 = ~n9454 | ~n9453;
  assign n7399 = ~n7570 | ~n8949;
  assign n8629 = ~n8628 & ~n8627;
  assign n8666 = ~n8665 | ~n8664;
  assign n7484 = ~n7480;
  assign n8582 = ~n8581 | ~n8580;
  assign n10468 = ~n8824 & ~n8823;
  assign n7480 = ~n7452 | ~STATE2_REG_0__SCAN_IN;
  assign n7419 = ~n7417 & ~n7416;
  assign n7570 = ~n10077;
  assign n8751 = ~n8711 & ~n8710;
  assign n7368 = ~n7367 | ~n7366;
  assign n9067 = ~n9696;
  assign n8627 = ~n8626 | ~n8625;
  assign n9139 = ~n7316 | ~n7996;
  assign n7367 = ~n7363 | ~n7362;
  assign n7381 = n7341 & n7340;
  assign n8711 = ~n8670 | ~PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n10077 = ~n8946 & ~n10245;
  assign n8084 = ~n8081 | ~n8080;
  assign n7474 = ~n7473 & ~n7472;
  assign n8081 = ~n8060 & ~n8059;
  assign n7389 = ~n7406;
  assign n9096 = ~n9095 | ~n9094;
  assign n8821 = ~n8820 | ~n10934;
  assign n8541 = ~n12868;
  assign n7362 = n7361 & n7360;
  assign n8143 = ~n8142 | ~n8141;
  assign n8670 = ~n8663 & ~n12707;
  assign n7405 = ~n7403 | ~n7402;
  assign n7964 = ~n8044;
  assign n7366 = ~n7365 | ~n7364;
  assign n8116 = ~n8115 & ~n8114;
  assign n7371 = ~n7346 & ~n7356;
  assign n8345 = ~n8309 | ~n8342;
  assign n8071 = ~n8070 | ~n8069;
  assign n7468 = ~n7467 & ~n7466;
  assign n7513 = ~n7418 & ~n7314;
  assign n7417 = ~n7507 & ~n7415;
  assign n8122 = ~n8121 & ~n8120;
  assign n10983 = ~n8274 | ~n8306;
  assign n8141 = ~n8140 & ~n8139;
  assign n7341 = ~n7401 | ~n7336;
  assign n7369 = ~n7348 & ~n7347;
  assign n10824 = ~n8191 | ~n8229;
  assign n8430 = ~n8422 | ~n8421;
  assign n8156 = ~n8155 & ~n8154;
  assign n8663 = ~n8624 | ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n8059 = ~n8041 | ~n7887;
  assign n7360 = ~n7359 | ~n7358;
  assign n7374 = ~n7404 | ~n7373;
  assign n7402 = ~n7401 & ~n7400;
  assign n10821 = ~n8266 & ~n7009;
  assign n7445 = ~n7444 & ~n7466;
  assign n8044 = ~n7958 | ~n7957;
  assign n8342 = ~n8341 | ~n8340;
  assign n8172 = ~n8171 & ~n8170;
  assign n8229 = ~n8341 | ~n8228;
  assign n7623 = ~n7616 | ~n7615;
  assign n8306 = ~n8341 | ~n8305;
  assign n7314 = ~n7313 | ~n7312;
  assign n7448 = ~n8949 & ~n10937;
  assign n7433 = ~n7432 | ~n7431;
  assign n7507 = ~n7414 | ~n7443;
  assign n8041 = ~n7856 & ~n8032;
  assign n8384 = ~n8380 & ~n7015;
  assign n8472 = ~n8471 & ~n7014;
  assign n8046 = ~n7963 & ~n7962;
  assign n8421 = ~n8420 & ~n8419;
  assign n7321 = ~n8949 & ~n7320;
  assign n7968 = ~n8058 | ~n7966;
  assign n7472 = ~n7471 | ~n7470;
  assign n7384 = ~n7383 | ~n11628;
  assign n8493 = ~n8802 | ~n11647;
  assign n8537 = ~n8536 & ~n7013;
  assign n7954 = ~n7953 & ~n7952;
  assign n7993 = ~n7991;
  assign n8154 = ~n8153 | ~n8152;
  assign n9500 = ~n9458 & ~n9457;
  assign n7346 = ~n7344 & ~n7343;
  assign n8803 = ~n8802 | ~n8801;
  assign n8624 = ~n8539 & ~n12821;
  assign n8070 = ~n8067 & ~n8066;
  assign n8130 = ~n8110 | ~n8109;
  assign n9391 = ~n9390 | ~n9389;
  assign n8830 = ~n8829 | ~n8828;
  assign n7991 = ~n7926 | ~n7925;
  assign n8881 = ~n8880 | ~n8879;
  assign n8827 = ~n8826 | ~n8825;
  assign n9197 = ~n9196 | ~n9195;
  assign n8813 = ~n8812 | ~n8811;
  assign n8032 = ~n8020 | ~n8019;
  assign n8884 = ~n8883 | ~n8882;
  assign n9194 = ~n9193 | ~n9192;
  assign n8139 = ~n8138 | ~n8137;
  assign n8848 = ~n8847 | ~n8846;
  assign n8110 = ~n8147 | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n8083 = ~n8090 & ~n8082;
  assign n8872 = ~n8871 | ~n8870;
  assign n7461 = ~n7460 | ~n7459;
  assign n7388 = ~n8068 | ~n8092;
  assign n9131 = ~n7482 | ~n7481;
  assign n8164 = ~n8163 | ~n8162;
  assign n7435 = ~n7436 & ~n7601;
  assign n9457 = ~n9418 | ~n9417;
  assign n8851 = ~n8850 | ~n8849;
  assign n8869 = ~n8868 | ~n8867;
  assign n7385 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n7382;
  assign n7966 = ~n7959;
  assign n8842 = ~n8841 | ~n8840;
  assign n8170 = ~n8169 | ~n8168;
  assign n8875 = ~n8874 | ~n8873;
  assign n8309 = n8308 & n8307;
  assign n7442 = ~n7441;
  assign n8949 = ~n7319 | ~n8008;
  assign n8854 = ~n8853 | ~n8852;
  assign n7432 = ~n7428 | ~n9102;
  assign n8274 = n8273 & n8272;
  assign n9711 = ~n9710 | ~n9709;
  assign n8833 = ~n8832 | ~n8831;
  assign n8845 = ~n8844 | ~n8843;
  assign n8878 = ~n8877 | ~n8876;
  assign n7930 = ~n7932 & ~n7929;
  assign n8266 = ~n8193 & ~n8260;
  assign n8857 = ~n8856 | ~n8855;
  assign n8839 = ~n8838 | ~n8837;
  assign n8191 = n8190 & n8189;
  assign n7933 = ~n7932 & ~n8003;
  assign n7313 = ~n7311 | ~n11637;
  assign n8264 = ~n8263 | ~n8262;
  assign n8863 = ~n8862 | ~n8861;
  assign n8836 = ~n8835 | ~n8834;
  assign n8182 = ~n8181 | ~n8180;
  assign n13186 = ~n9722 | ~n9721;
  assign n8866 = ~n8865 | ~n8864;
  assign n7471 = ~n7199 | ~n10076;
  assign n9394 = ~n9393 | ~n9392;
  assign n7616 = n7612 & n7611;
  assign n8341 = ~n8193;
  assign n8860 = ~n8859 | ~n8858;
  assign n8492 = ~n8490 | ~n8489;
  assign n9418 = ~n9260 & ~n9259;
  assign n7431 = ~n7430 | ~n7429;
  assign n8747 = ~n8746 & ~n8745;
  assign n8705 = ~n8704 & ~n8703;
  assign n7396 = ~n7394;
  assign n8068 = ~n7961;
  assign n9093 = ~n8796;
  assign n7428 = ~n8491 | ~n7427;
  assign n8787 = ~n8786 & ~n8785;
  assign n7436 = ~n7465;
  assign n8928 = ~n8927 & ~n8926;
  assign n8825 = ~n10932 | ~EBX_REG_2__SCAN_IN;
  assign n8019 = ~n7976 | ~n8002;
  assign n8189 = ~n8188 & ~n8187;
  assign n8501 = ~n8435 & ~n8434;
  assign n8272 = ~n8271 & ~n8270;
  assign n7992 = ~n7919 | ~n7928;
  assign n8193 = ~n9633 | ~n8192;
  assign n7926 = ~n7923 | ~n7922;
  assign n8580 = ~n8579 & ~n8578;
  assign n8308 = ~n9707 | ~EAX_REG_11__SCAN_IN;
  assign n8263 = ~n9707 | ~EAX_REG_9__SCAN_IN;
  assign n8109 = ~n8108 & ~n8107;
  assign n8422 = ~n9707 | ~EAX_REG_13__SCAN_IN;
  assign n8162 = ~n8161 & ~n8160;
  assign n8180 = ~n8179 & ~n8178;
  assign n8152 = ~n8151 & ~n8150;
  assign n7430 = ~n9132 & ~n9102;
  assign n8092 = ~n8082;
  assign n8344 = ~n12463 & ~n9789;
  assign n7333 = n7372 & INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n8491 = ~n7614;
  assign n8819 = ~n8817 & ~n8816;
  assign n8002 = ~n7855 | ~n7854;
  assign n7318 = ~n8791 | ~n7231;
  assign n7335 = ~n8065;
  assign n9110 = ~n8488 & ~n8101;
  assign n7395 = ~n7508 | ~n10748;
  assign n9707 = ~n9686;
  assign n10240 = ~n10076;
  assign n7356 = ~n7345 | ~n7601;
  assign n7337 = ~n9092 & ~n10490;
  assign n7464 = ~n9092 & ~n10748;
  assign n8065 = ~n9092 | ~STATE2_REG_0__SCAN_IN;
  assign n8812 = ~n10937 | ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n7508 = ~n9102;
  assign n9132 = ~n7231;
  assign n8228 = ~n8227 | ~n8226;
  assign n8058 = ~n7703 | ~n7702;
  assign n8488 = ~n9102 | ~n10748;
  assign n7315 = ~n13389 & ~n7231;
  assign n7929 = ~n8079;
  assign n8418 = ~n8414 & ~n8413;
  assign n8376 = ~n8375 & ~n8374;
  assign n8004 = ~n7823 & ~n7822;
  assign n9723 = ~n10515 | ~n8814;
  assign n7702 = ~n7701 & ~n7700;
  assign n7950 = ~n7763 & ~n7762;
  assign n10245 = ~n10515;
  assign n10748 = ~n8814;
  assign n8260 = ~n8259 & ~n8258;
  assign n7732 = ~n7731 & ~n7730;
  assign n8226 = ~n8225 & ~n8224;
  assign n7332 = ~n7331 | ~n7330;
  assign n7792 = ~n7791 | ~n7790;
  assign n7731 = ~n7723 | ~n7722;
  assign n7762 = ~n7761 | ~n7760;
  assign n7701 = ~n7697 | ~n7696;
  assign n7823 = ~n7807 | ~n7806;
  assign n8267 = ~n8261 & ~n7670;
  assign n7703 = ~n7683 & ~n7682;
  assign n7117 = ~n7101 | ~n7100;
  assign n7822 = ~n7821 | ~n7820;
  assign n8259 = ~n8243 | ~n8242;
  assign n7885 = ~n7884 | ~n7883;
  assign n7330 = ~n7329 | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n7917 = ~n7916 | ~n7915;
  assign n8258 = ~n8257 | ~n8256;
  assign n7886 = ~n7870 | ~n7869;
  assign n7793 = ~n7777 | ~n7776;
  assign n8413 = ~n8412 | ~n8411;
  assign n7853 = ~n7837 | ~n7836;
  assign n7852 = ~n7851 | ~n7850;
  assign n7763 = ~n7747 | ~n7746;
  assign n7918 = ~n7902 | ~n7901;
  assign n8414 = ~n8398 | ~n8397;
  assign n7722 = ~n7721 & ~n7720;
  assign n7723 = ~n7715 & ~n7714;
  assign n7884 = ~n7876 & ~n7875;
  assign n7310 = ~n7284 & ~n7283;
  assign n7309 = ~n7308 & ~n7307;
  assign n7836 = ~n7835 & ~n7834;
  assign n7790 = ~n7789 & ~n7788;
  assign n7883 = ~n7882 & ~n7881;
  assign n7777 = ~n7769 & ~n7768;
  assign n7902 = ~n7894 & ~n7893;
  assign n7851 = ~n7843 & ~n7842;
  assign n7916 = ~n7908 & ~n7907;
  assign n7850 = ~n7849 & ~n7848;
  assign n7791 = ~n7783 & ~n7782;
  assign n7901 = ~n7900 & ~n7899;
  assign n7776 = ~n7775 & ~n7774;
  assign n7733 = ~n7709 & ~n7708;
  assign n8227 = ~n8207 & ~n8206;
  assign n7806 = ~n7805 & ~n7804;
  assign n7761 = ~n7753 & ~n7752;
  assign n7683 = ~n7679 | ~n7678;
  assign n7807 = ~n7799 & ~n7798;
  assign n7821 = ~n7813 & ~n7812;
  assign n7760 = ~n7759 & ~n7758;
  assign n7697 = ~n7689 & ~n7688;
  assign n7746 = ~n7745 & ~n7744;
  assign n7696 = ~n7695 & ~n7694;
  assign n7213 = ~n7205 & ~n7204;
  assign n7212 = ~n7211 & ~n7210;
  assign n8261 = ~n8184 | ~PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n7227 = ~n7219 & ~n7218;
  assign n7226 = ~n7225 & ~n7224;
  assign n7820 = ~n7819 & ~n7818;
  assign n7747 = ~n7739 & ~n7738;
  assign n8256 = ~n8255 & ~n8254;
  assign n7837 = ~n7829 & ~n7828;
  assign n8257 = ~n8249 & ~n8248;
  assign n7870 = ~n7862 & ~n7861;
  assign n7245 = ~n7237 & ~n7236;
  assign n7915 = ~n7914 & ~n7913;
  assign n8242 = ~n8241 & ~n8240;
  assign n7244 = ~n7243 & ~n7242;
  assign n7869 = ~n7868 & ~n7867;
  assign n8243 = ~n8235 & ~n8234;
  assign n7259 = ~n7251 & ~n7250;
  assign n7258 = ~n7257 & ~n7256;
  assign n7196 = ~n7187 | ~n7186;
  assign n7237 = ~n7233 | ~n7232;
  assign n7829 = ~n7825 | ~n7824;
  assign n7054 = ~n7053 | ~n7052;
  assign n7243 = ~n7239 | ~n7238;
  assign n7720 = ~n7719 | ~n7718;
  assign n7236 = ~n7235 | ~n7234;
  assign n7818 = ~n7817 | ~n7816;
  assign n7137 = ~n7127 | ~n7126;
  assign n7862 = ~n7858 | ~n7857;
  assign n7819 = ~n7815 | ~n7814;
  assign n7721 = ~n7717 | ~n7716;
  assign n7812 = ~n7811 | ~n7810;
  assign n7729 = ~n7725 | ~n7724;
  assign n7504 = ~n7503 | ~n7502;
  assign n7913 = ~n7912 | ~n7911;
  assign n7700 = ~n7699 | ~n7698;
  assign n7156 = ~n7155 | ~n7154;
  assign n7813 = ~n7809 | ~n7808;
  assign n7728 = ~n7727 | ~n7726;
  assign n7694 = ~n7693 | ~n7692;
  assign n7758 = ~n7757 | ~n7756;
  assign n7804 = ~n7803 | ~n7802;
  assign n7695 = ~n7691 | ~n7690;
  assign n7759 = ~n7755 | ~n7754;
  assign n7805 = ~n7801 | ~n7800;
  assign n7799 = ~n7795 | ~n7794;
  assign n7688 = ~n7687 | ~n7686;
  assign n7689 = ~n7685 | ~n7684;
  assign n7798 = ~n7797 | ~n7796;
  assign n7093 = ~n7089 | ~n7088;
  assign n7709 = ~n7705 | ~n7704;
  assign n7848 = ~n7847 | ~n7846;
  assign n7077 = ~n7073 | ~n7072;
  assign n7849 = ~n7845 | ~n7844;
  assign n7708 = ~n7707 | ~n7706;
  assign n7842 = ~n7841 | ~n7840;
  assign n7893 = ~n7892 | ~n7891;
  assign n7062 = ~n7061 | ~n7060;
  assign n7843 = ~n7839 | ~n7838;
  assign n7881 = ~n7880 | ~n7879;
  assign n7900 = ~n7896 | ~n7895;
  assign n7834 = ~n7833 | ~n7832;
  assign n7835 = ~n7831 | ~n7830;
  assign n7307 = ~n7306 | ~n7305;
  assign n7899 = ~n7898 | ~n7897;
  assign n7882 = ~n7878 | ~n7877;
  assign n7875 = ~n7874 | ~n7873;
  assign n7876 = ~n7872 | ~n7871;
  assign n7113 = ~n7109 | ~n7108;
  assign n7867 = ~n7866 | ~n7865;
  assign n7715 = ~n7711 | ~n7710;
  assign n7284 = ~n7272 | ~n7271;
  assign n7828 = ~n7827 | ~n7826;
  assign n7908 = ~n7904 | ~n7903;
  assign n7868 = ~n7864 | ~n7863;
  assign n7907 = ~n7906 | ~n7905;
  assign n7894 = ~n7890 | ~n7889;
  assign n7256 = ~n7255 | ~n7254;
  assign n7257 = ~n7253 | ~n7252;
  assign n7714 = ~n7713 | ~n7712;
  assign n7251 = ~n7247 | ~n7246;
  assign n7177 = ~n7176 | ~n7175;
  assign n7914 = ~n7910 | ~n7909;
  assign n7861 = ~n7860 | ~n7859;
  assign n7774 = ~n7773 | ~n7772;
  assign n8184 = ~n8176 & ~n12415;
  assign n7775 = ~n7771 | ~n7770;
  assign n7744 = ~n7743 | ~n7742;
  assign n7745 = ~n7741 | ~n7740;
  assign n7738 = ~n7737 | ~n7736;
  assign n7782 = ~n7781 | ~n7780;
  assign n7679 = n7674 & n7673;
  assign n7788 = ~n7787 | ~n7786;
  assign n7739 = ~n7735 | ~n7734;
  assign n7768 = ~n7767 | ~n7766;
  assign n7753 = ~n7749 | ~n7748;
  assign n7682 = ~n7681 | ~n7680;
  assign n7789 = ~n7785 | ~n7784;
  assign n7769 = ~n7765 | ~n7764;
  assign n7752 = ~n7751 | ~n7750;
  assign n7327 = ~n7349 & ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n7064 = ~n9653 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n7811 = ~n9653 | ~INSTQUEUE_REG_4__0__SCAN_IN;
  assign n7103 = ~n9501 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n7202 = ~n7002 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n7272 = ~n7265 & ~n7264;
  assign n7271 = ~n7270 & ~n7269;
  assign n7282 = ~n7276 & ~n7275;
  assign n7281 = ~n7280 & ~n7279;
  assign n7889 = ~n9501 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n7296 = ~n7290 & ~n7289;
  assign n7295 = ~n7294 & ~n7293;
  assign n7306 = ~n7301 & ~n7300;
  assign n7247 = ~n9636 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n7305 = ~n7304 & ~n7303;
  assign n7892 = ~n9599 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n7891 = ~n9673 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n7503 = ~n11440 | ~n7500;
  assign n7239 = ~n9648 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n7896 = ~n9672 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n7895 = ~n9647 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n7234 = ~n9653 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n7898 = ~n9602 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n7897 = ~n9522 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n7052 = ~n7051 & ~n7050;
  assign n7904 = ~n9648 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n7903 = ~n9636 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n7053 = ~n7047 & ~n7046;
  assign n7041 = ~n7040 & ~n7039;
  assign n7906 = ~n9665 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n7905 = ~n9653 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n7783 = ~n7779 | ~n7778;
  assign n7042 = ~n7036 & ~n7035;
  assign n7910 = ~n9656 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n7678 = ~n7677 & ~n7676;
  assign n7699 = ~n9522 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n7698 = ~n9636 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n8176 = ~n8167 | ~PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n13417 = ~n13222 & ~n13221;
  assign n7276 = ~n8195 & ~n7273;
  assign n7275 = ~n8196 & ~n7274;
  assign n7280 = ~n8585 & ~n7277;
  assign n11877 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n11730;
  assign n7233 = ~n9662 | ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n8378 = ~n9535 & ~n8382;
  assign n7304 = ~n8593 & ~n7302;
  assign n7269 = ~n8591 & ~n7268;
  assign n10585 = ~n11488 & ~n12050;
  assign n7290 = ~n7286 & ~n7285;
  assign n10489 = ~n10487 | ~n10486;
  assign n7300 = ~n7299 & ~n7298;
  assign n7293 = ~n9053 & ~n7292;
  assign n7265 = ~n9640 & ~n7262;
  assign n7680 = ~n9607 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n7270 = ~n7267 & ~n7266;
  assign n7264 = ~n8587 & ~n7263;
  assign n9672 = ~n7267;
  assign n7289 = ~n7288 & ~n7287;
  assign n12690 = ~n10057 & ~n9789;
  assign n12691 = ~n10074;
  assign n7493 = ~n7492 & ~n7491;
  assign n10893 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n10892;
  assign n7478 = ~n7477 & ~n7476;
  assign n7502 = ~n7501 | ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n11700 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n11451;
  assign n7641 = ~n9855;
  assign n7456 = ~n7455 | ~n7454;
  assign n11269 = ~n11488 & ~n11451;
  assign n12271 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n12139;
  assign n7051 = ~n8591 & ~n7049;
  assign n7046 = ~n8593 & ~n7045;
  assign n7047 = ~n7286 & ~n7044;
  assign n7040 = ~n7288 & ~n7037;
  assign n10615 = ~n11488 & ~n10892;
  assign n7035 = ~n8196 & ~n7034;
  assign n7036 = ~n8585 & ~n7033;
  assign n7890 = ~n9662 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n7909 = ~n9607 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n7810 = ~n9607 | ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n7165 = ~n8591 & ~n7164;
  assign n7192 = ~n8593 & ~n9056;
  assign n8270 = ~n9535 & ~n8269;
  assign n7140 = ~n7286 & ~n8584;
  assign n7121 = ~n9640 & ~n7118;
  assign n7166 = ~n7267 & ~n8548;
  assign n7189 = ~n7299 & ~n8199;
  assign n7133 = ~n8585 & ~n8592;
  assign n7172 = ~n8195 & ~n7169;
  assign n7120 = ~n8587 & ~n7119;
  assign n7149 = ~n7299 & ~n7148;
  assign n9647 = ~n8587;
  assign n9673 = ~n8591;
  assign n7139 = ~n7288 & ~n7138;
  assign n8167 = ~n8159 & ~n12638;
  assign n7171 = ~n8196 & ~n7170;
  assign n7129 = ~n8196 & ~n7128;
  assign n7125 = ~n7267 & ~n7122;
  assign n7162 = ~n8587 & ~n7161;
  assign n7184 = ~n9053 & ~n7183;
  assign n7163 = ~n9640 & ~n7160;
  assign n8959 = ~n11975 & ~n8941;
  assign n7143 = ~n9053 & ~n7142;
  assign n7182 = ~n7286 & ~n7179;
  assign n7174 = ~n8585 & ~n9052;
  assign n7153 = ~n8593 & ~n7151;
  assign n12243 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n12050;
  assign n11284 = ~n11488 & ~n11730;
  assign n7124 = ~n8591 & ~n7123;
  assign n7181 = ~n7288 & ~n7180;
  assign n7130 = ~n8195 & ~n8590;
  assign n8187 = ~n9535 & ~n8186;
  assign n11247 = ~n11488 & ~n12316;
  assign n7455 = ~n7665 | ~n11488;
  assign n7173 = ~n9642 & ~n8194;
  assign n7050 = ~n8551 & ~n7960;
  assign n12562 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n12316;
  assign n7132 = ~n9642 & ~n7131;
  assign n8943 = ~n10486 & ~n7655;
  assign n11258 = ~n11488 & ~n11979;
  assign n7325 = ~n7326 & ~n8111;
  assign n9535 = ~n9708;
  assign n7477 = ~n11441 & ~n7665;
  assign n7499 = ~n7498 & ~n12145;
  assign n10074 = ~n9787 | ~STATE2_REG_0__SCAN_IN;
  assign n11357 = n12145 & n7498;
  assign n7279 = ~n9642 & ~n7278;
  assign n7152 = ~n8551 & ~n8586;
  assign n11445 = ~STATEBS16_REG_SCAN_IN & ~n11480;
  assign n7492 = ~n7665 & ~n10898;
  assign n12131 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n11979;
  assign n8159 = ~n8146 | ~PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n7303 = ~n8551 & ~n7951;
  assign n7039 = ~n9642 & ~n7038;
  assign n10485 = ~n11497 & ~n11813;
  assign n7323 = ~n11488 | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n10374 = ~n10341;
  assign n13515 = STATE_REG_1__SCAN_IN & n9861;
  assign n10486 = ~n11497 | ~n11813;
  assign n10034 = ~n11813 | ~n12305;
  assign n9789 = ~n9698;
  assign n11809 = ~STATEBS16_REG_SCAN_IN | ~n12305;
  assign n7043 = ~n8118 & ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n8146 = ~n8134 & ~n12576;
  assign n11480 = ~n12305;
  assign n7665 = ~n12681 | ~n10490;
  assign n8958 = ~n12447 & ~n12650;
  assign n12821 = ~PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n8269 = ~PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n10638 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n8586 = ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n11488 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n12502 = ~INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n10490 = ~STATE2_REG_0__SCAN_IN;
  assign n11628 = ~INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n12324 = ~STATE2_REG_3__SCAN_IN;
  assign n11497 = ~STATE2_REG_2__SCAN_IN;
  assign n11813 = ~STATE2_REG_1__SCAN_IN;
  assign n7393 = ~STATE_REG_2__SCAN_IN;
  assign n13257 = ~INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n13112 = ~INSTADDRPOINTER_REG_17__SCAN_IN | ~INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n8134 = ~PHYADDRPOINTER_REG_1__SCAN_IN | ~PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n8891 = ~PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n8963 = ~STATEBS16_REG_SCAN_IN & ~READY_N;
  assign n9056 = ~INSTQUEUE_REG_3__0__SCAN_IN;
  assign n10637 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n9058 = ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n7497 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n11478 = ~STATEBS16_REG_SCAN_IN;
  assign n12681 = ~STATE2_REG_3__SCAN_IN & ~STATE2_REG_1__SCAN_IN;
  assign n13498 = ~n13497 & ~n13496;
  assign n9757 = ~n13505 & ~n13465;
  assign n9782 = ~n9771 | ~n9770;
  assign n13505 = n9750 ^ n9749;
  assign n13496 = ~n13495 | ~n13494;
  assign n13447 = ~n13466 & ~n13504;
  assign n13495 = ~n13488 | ~n9141;
  assign n13476 = ~n13466 & ~n13465;
  assign n9769 = ~n9760 & ~n13504;
  assign n13466 = n13439 ^ INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n13488 = ~n13347 ^ n13346;
  assign n9554 = ~n9760 & ~n13465;
  assign n13347 = ~n9742 | ~n9741;
  assign n13362 = ~n13246 & ~n13245;
  assign n13458 = ~n13454 & ~n13465;
  assign n9760 = ~n9415 ^ n9414;
  assign n13246 = ~n13239 & ~n13241;
  assign n13438 = ~n13430 & ~n13429;
  assign n13454 = n13430 ^ n13405;
  assign n13381 = ~n13149 ^ n13148;
  assign n9580 = ~n9740 | ~n9576;
  assign n13307 = ~n9141 | ~n13305;
  assign n13170 = ~n13160 & ~n13465;
  assign n13149 = ~n13145 | ~n13144;
  assign n13245 = ~n13244 & ~n13243;
  assign n13261 = ~n13081 | ~n13145;
  assign n9388 = ~n9141 | ~n13159;
  assign n13220 = ~n13216 | ~n13215;
  assign n13404 = ~n13436 | ~n13402;
  assign n13305 = n13436 ^ n13289;
  assign n13216 = ~n13077 | ~n9573;
  assign n13159 = n9406 ^ n9387;
  assign n9409 = ~n9406 | ~n9405;
  assign n13287 = ~n13281 | ~n13280;
  assign n13395 = ~n13393 | ~n13392;
  assign n13058 = ~n9141 | ~n13056;
  assign n13281 = ~n13270;
  assign n12921 = ~n13056 | ~n13348;
  assign n13115 = n12987 ^ n12986;
  assign n9386 = ~n13270 | ~n9382;
  assign n9338 = ~n9141 | ~n12862;
  assign n12872 = ~n12862 | ~n13348;
  assign n12898 = ~n13005 | ~n13348;
  assign n13393 = ~n13390 | ~n13391;
  assign n13007 = ~n9141 | ~n13005;
  assign n12987 = ~n12983 & ~n12982;
  assign n9738 = ~n9737 | ~n9736;
  assign n13100 = ~n13331 | ~n13176;
  assign n13478 = ~n13464 | ~n13463;
  assign n13108 = ~n13331 | ~n13185;
  assign n9737 = ~n13464 | ~n13330;
  assign n13184 = ~n13450 | ~n13176;
  assign n9337 = ~n12889 & ~n9332;
  assign n13021 = ~n13132 | ~n13185;
  assign n9552 = ~n13132 | ~n13463;
  assign n13017 = ~n13132 | ~n13176;
  assign n13195 = ~n13450 | ~n13185;
  assign n12969 = ~n13232 | ~n13176;
  assign n13238 = ~n13232 | ~n13463;
  assign n13073 = ~n13232 | ~n13330;
  assign n12977 = ~n13232 | ~n13185;
  assign n13450 = n13175 ^ n13174;
  assign n13094 = ~n13174;
  assign n9546 = ~n12963 & ~n9545;
  assign n12925 = ~n13171 | ~n13185;
  assign n13093 = ~n13092 & ~n13091;
  assign n12887 = ~n12881 | ~n13185;
  assign n13172 = ~n13171 | ~n13463;
  assign n12908 = ~n13171 | ~n13176;
  assign n9306 = ~n13176 | ~n12881;
  assign n13034 = ~n13171 | ~n13330;
  assign n9331 = ~n9149 | ~n9150;
  assign n13092 = ~n9543 & ~n9544;
  assign n12880 = ~n12873 | ~n13185;
  assign n9254 = ~n13176 | ~n12873;
  assign n12950 = ~n12946 & ~n12945;
  assign n9543 = ~n12961 | ~n12960;
  assign n9153 = ~n9152 | ~n9151;
  assign n12962 = ~n12961 & ~n12960;
  assign n9083 = ~n13176 | ~n12859;
  assign n12937 = ~n12946 & ~n13349;
  assign n12860 = ~n13185 | ~n12859;
  assign n12945 = ~n9304 | ~n12899;
  assign n13356 = ~n13349 & ~n13451;
  assign n13320 = ~n13319 & ~n13451;
  assign n12901 = ~n12900 | ~n12899;
  assign n9202 = ~n12946 & ~n13319;
  assign n12845 = ~n13504 & ~n12844;
  assign n12899 = ~n9303 | ~n9302;
  assign n13319 = ~n9081 | ~n9250;
  assign n9143 = ~n8480 | ~n8479;
  assign n12854 = ~n13185 | ~n12853;
  assign n9252 = ~n9251 | ~n9250;
  assign n12763 = ~n9141 | ~n12761;
  assign n8936 = ~n13176 | ~n12853;
  assign n8425 = ~n13348 | ~n12761;
  assign n13083 = ~n13082 & ~n13451;
  assign n12787 = ~n8806 & ~n13082;
  assign n13228 = ~n13227 & ~n13451;
  assign n8809 = ~n13185 | ~n8807;
  assign n8795 = ~n13176 | ~n8807;
  assign n12800 = ~n12799 & ~n13082;
  assign n9250 = ~n9080 | ~n9079;
  assign n9320 = ~n12946 & ~n13227;
  assign n8987 = ~n12946 & ~n13082;
  assign n12747 = ~n13465 & ~n12776;
  assign n12777 = ~n13504 & ~n12776;
  assign n9175 = ~n12946 & ~n13150;
  assign n13151 = ~n13150 & ~n13451;
  assign n13525 = ~n8806 & ~n13520;
  assign n8998 = ~n8973 | ~n8933;
  assign n12738 = ~n12946 & ~n13520;
  assign n12660 = ~n12799 & ~n13520;
  assign n12701 = ~n13185 | ~n12913;
  assign n12813 = ~n13330 | ~n12913;
  assign n12989 = ~n12988 | ~n13463;
  assign n8976 = ~n8975 | ~n8974;
  assign n8973 = ~n8975 & ~n8974;
  assign n12791 = ~n13176 | ~n12913;
  assign n12914 = ~n12913 | ~n13463;
  assign n12665 = ~n12946 & ~n12863;
  assign n12988 = ~n12656 & ~n12700;
  assign n12891 = ~n13526 & ~n13451;
  assign n12480 = ~n8806 & ~n12863;
  assign n13532 = ~n8806 & ~n13526;
  assign n12470 = ~n13348 | ~n12512;
  assign n8975 = ~n12700 | ~n8709;
  assign n12533 = ~n12799 & ~n13526;
  assign n12703 = ~n12946 & ~n13526;
  assign n12864 = ~n12863 & ~n13451;
  assign n12487 = ~n12799 & ~n12863;
  assign n12516 = ~n9141 | ~n12512;
  assign n12656 = n12655 & n12654;
  assign n12863 = ~n12479 | ~n12478;
  assign n13526 = ~n12529 | ~n12655;
  assign n12823 = ~n12822 & ~n13451;
  assign n12097 = ~n12799 & ~n12822;
  assign n12046 = ~n8806 & ~n12822;
  assign n12494 = ~n13504 & ~n12491;
  assign n12039 = ~n12946 & ~n12822;
  assign n12439 = ~n13465 & ~n12491;
  assign n12610 = ~n13330 | ~n12602;
  assign n11755 = ~n12799 & ~n11752;
  assign n12528 = ~n12477 & ~n12476;
  assign n11595 = ~n8806 & ~n11752;
  assign n12478 = ~n12477 | ~n12476;
  assign n8424 = ~n11940 | ~n13463;
  assign n12694 = ~n12690 & ~n12689;
  assign n11929 = ~n9141 | ~n11928;
  assign n11585 = ~n8806 & ~n12601;
  assign n8474 = ~n12601 & ~n13451;
  assign n11840 = ~n13348 | ~n11928;
  assign n12602 = ~n12601;
  assign n11619 = ~n12799 & ~n12601;
  assign n12438 = ~n8096 | ~n8095;
  assign n13401 = ~n13507 | ~n13400;
  assign n11762 = ~n13465 & ~n11885;
  assign n13445 = ~n13490 & ~n13440;
  assign n11891 = ~n13504 & ~n11885;
  assign n8423 = ~n8432 | ~n8431;
  assign n11838 = ~n11761 | ~n8089;
  assign n8500 = ~n8433 | ~n8432;
  assign n13191 = ~n13189 & ~n13188;
  assign n12748 = ~n12742 & ~n13451;
  assign n7649 = ~n11831 | ~n12685;
  assign n8432 = ~n8417 | ~n8416;
  assign n12686 = ~n12685 | ~n12684;
  assign n11417 = ~n13465 & ~n11548;
  assign n11243 = ~n8806 & ~n12742;
  assign n7654 = ~n12685;
  assign n11280 = ~n12799 & ~n12742;
  assign n13343 = ~n13329 & ~n13328;
  assign n12742 = ~n11242 | ~n11241;
  assign n12411 = ~n12410 | ~n12409;
  assign n13308 = ~n13490 & ~n13328;
  assign n13106 = ~n13528 & ~n13328;
  assign n12685 = ~n7648 | ~STATE2_REG_2__SCAN_IN;
  assign n13189 = ~n9726 & ~n10045;
  assign n11241 = ~n11240 | ~n11239;
  assign n10990 = ~n8806 & ~n12434;
  assign n13141 = ~n13329 & ~n13131;
  assign n13328 = ~n13104 | ~n13103;
  assign n10994 = ~n12799 & ~n12434;
  assign n13019 = ~n13528 & ~n13131;
  assign n12474 = ~n12473 | ~n13463;
  assign n12693 = ~n12692 | ~n12691;
  assign n12440 = ~n12434 & ~n13451;
  assign n12975 = ~n13528 & ~n13365;
  assign n12692 = ~n7647 | ~n7646;
  assign n13131 = ~n13187 | ~n9764;
  assign n13075 = ~n13329 & ~n13365;
  assign n11240 = ~n11024 & ~n11023;
  assign n13366 = ~n13490 & ~n13365;
  assign n13204 = ~REIP_REG_30__SCAN_IN | ~n13202;
  assign n13538 = ~n8806 & ~n13533;
  assign n13365 = ~n12973 | ~n12972;
  assign n13206 = ~n13325 | ~n13201;
  assign n10828 = ~n12799 & ~n13533;
  assign n11763 = ~n13533 & ~n13451;
  assign n11661 = ~n11660 | ~n11659;
  assign n13065 = ~REIP_REG_27__SCAN_IN | ~n13125;
  assign n13067 = ~n13127 & ~REIP_REG_27__SCAN_IN;
  assign n11669 = ~n11668 | ~n11667;
  assign n11862 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n11861;
  assign n11685 = ~n11684 | ~n11683;
  assign n10984 = ~n10826 & ~n10821;
  assign n12541 = ~n12540 | ~n12539;
  assign n9576 = ~n9575;
  assign n7663 = ~n7643 & ~n10074;
  assign n12552 = ~n12551 | ~n12550;
  assign n7643 = ~n7636 & ~n7635;
  assign n12923 = ~n13528 & ~n13022;
  assign n12954 = ~n13023 & ~REIP_REG_25__SCAN_IN;
  assign n13028 = ~n13023;
  assign n9398 = ~n13490 & ~n13022;
  assign n12972 = ~n12971 | ~n12970;
  assign n13127 = ~n13023 | ~n9592;
  assign n12745 = ~n12744 | ~n12743;
  assign n12819 = ~n12818 | ~n12817;
  assign n9582 = ~n13490 & ~n12856;
  assign n9313 = ~REIP_REG_19__SCAN_IN | ~n12818;
  assign n8482 = ~n9142 | ~n9144;
  assign n11859 = ~n11627 | ~n11626;
  assign n10825 = ~n10666 & ~n10665;
  assign n11028 = ~n8054 & ~n8053;
  assign n12858 = ~n13528 & ~n12856;
  assign n12959 = ~n12944 | ~n13506;
  assign n12878 = ~n13528 & ~n13489;
  assign n12885 = ~n13559 | ~n13506;
  assign n13023 = ~n12929 & ~n9591;
  assign n12941 = ~n13329 & ~n13489;
  assign n13509 = ~n13507 | ~n13506;
  assign n9150 = ~n9329 & ~n9148;
  assign n9207 = ~n12931 & ~n9187;
  assign n9203 = ~n13329 & ~n12856;
  assign n13493 = ~n13490 & ~n13489;
  assign n9142 = ~n9147 | ~INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n13289 = ~n13402 | ~n13403;
  assign n9187 = ~n9186 | ~n12926;
  assign n12932 = ~n12931 | ~n12930;
  assign n9591 = ~REIP_REG_24__SCAN_IN | ~n12931;
  assign n12890 = ~n12978 | ~n12981;
  assign n11178 = ~n12330 | ~n10908;
  assign n8040 = ~n10565 | ~n10566;
  assign n12608 = ~n12721 & ~n12606;
  assign n13219 = ~n13218 | ~n13217;
  assign n11608 = ~n12330 | ~n11503;
  assign n8093 = ~n9147 & ~INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n12911 = ~n12910 & ~n12909;
  assign n12856 = ~n9201 | ~n9200;
  assign n12732 = ~REIP_REG_18__SCAN_IN & ~n12731;
  assign n12704 = ~n12731 & ~REIP_REG_17__SCAN_IN;
  assign n12818 = ~n8961 & ~n12731;
  assign n12978 = ~n13288 | ~INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n11295 = ~n10632 | ~n10631;
  assign n12268 = ~n12158 & ~n12157;
  assign n9381 = ~n13288 & ~n13283;
  assign n9378 = ~n13288 | ~n9377;
  assign n8052 = ~n8051;
  assign n12982 = ~n12981;
  assign n9413 = ~n13288 & ~INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n9329 = ~n9146 & ~n9349;
  assign n9186 = ~n9956 | ~n9185;
  assign n13402 = ~n13288 | ~INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n8094 = ~n9146 & ~n12502;
  assign n12678 = ~n12677 | ~n12676;
  assign n12436 = ~n9146 | ~n12501;
  assign n9179 = ~n13329 & ~n13384;
  assign n12731 = ~REIP_REG_16__SCAN_IN | ~n12677;
  assign n11873 = ~n11747 & ~n11746;
  assign n11706 = ~n11448 & ~n11447;
  assign n12910 = ~n13288 & ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n13385 = ~n13490 & ~n13384;
  assign n8889 = ~n13528 & ~n13384;
  assign n9373 = ~n12984 | ~n12981;
  assign n11831 = ~n11623 | ~n10485;
  assign n12127 = ~n11996 & ~n11995;
  assign n12743 = ~n13434 | ~n12771;
  assign n11248 = ~n10510 | ~n10509;
  assign n12466 = ~n13434 | ~n12770;
  assign n11358 = ~n10800 | ~n10799;
  assign n12677 = ~n8960 & ~n12604;
  assign n10350 = ~n8165 & ~n8164;
  assign n8051 = ~n8050 & ~n8049;
  assign n12605 = ~n12604 & ~n12603;
  assign n11259 = ~n10560 | ~n10559;
  assign n11944 = ~n12604 & ~REIP_REG_13__SCAN_IN;
  assign n12852 = ~n13528 & ~n13419;
  assign n8072 = ~n8175 & ~n8082;
  assign n7972 = ~n7971;
  assign n8183 = ~n8175 & ~n8174;
  assign n9745 = ~n13434 | ~n13481;
  assign n9743 = ~n13434 & ~n13481;
  assign n9566 = ~n13434 & ~n9565;
  assign n13403 = ~n13434 | ~n13432;
  assign n13241 = ~n13434 & ~n9410;
  assign n13302 = ~n13398 | ~n13301;
  assign n12984 = ~n13434 | ~n13109;
  assign n9407 = ~n13434 & ~n13274;
  assign n13286 = ~n13434 | ~n13285;
  assign n13146 = ~n13434 & ~n13370;
  assign n9185 = ~REIP_REG_22__SCAN_IN | ~n9184;
  assign n9324 = ~n13329 & ~n13419;
  assign n13278 = ~n13434 & ~n13277;
  assign n11623 = ~n7640 & ~n7639;
  assign n9747 = ~n13434 & ~n13272;
  assign n11306 = ~n10602 | ~n10601;
  assign n9741 = ~n13434 | ~n13480;
  assign n9200 = ~n9199 | ~n9198;
  assign n13240 = ~n13434 | ~n9410;
  assign n13217 = ~n13434 | ~n13414;
  assign n10460 = ~n8173 | ~n8172;
  assign n9122 = ~n12833 & ~n9348;
  assign n8049 = ~n8158 & ~n8082;
  assign n8038 = ~n8039;
  assign n8029 = ~n8028;
  assign n13054 = ~n13256 & ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n13487 = ~n13256 | ~n9561;
  assign n8888 = ~n9316;
  assign n13398 = ~n9758 & ~n9773;
  assign n13434 = ~n8091 | ~n8083;
  assign n11377 = ~n10694 | ~n10693;
  assign n8887 = ~n8886 | ~n8885;
  assign n13121 = ~n13114 & ~n13113;
  assign n12712 = ~n12706 & ~n12721;
  assign n11270 = ~n10654 | ~n10653;
  assign n13265 = ~n13490 & ~n13264;
  assign n10903 = ~n10902 | ~n7012;
  assign n10351 = ~n10313 | ~n10312;
  assign n9171 = ~REIP_REG_19__SCAN_IN | ~n12722;
  assign n12786 = ~n13528 & ~n13264;
  assign n9401 = ~n13501 | ~n9372;
  assign n11285 = ~n10538 | ~n10537;
  assign n12810 = ~n12722 & ~n12721;
  assign n8039 = ~n8036 | ~INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n8993 = ~n13329 & ~n13264;
  assign n13256 = ~n13114 & ~n13112;
  assign n8158 = ~n8048 | ~n8062;
  assign n13060 = ~n13490 & ~n13059;
  assign n8017 = ~n10327 | ~n10328;
  assign n8036 = ~n8035 | ~n8034;
  assign n8064 = ~n8062;
  assign n11477 = ~n11476 & ~n11475;
  assign n8166 = ~n8062 ^ n8063;
  assign n8048 = ~n8047 | ~n8046;
  assign n10598 = ~n12305 | ~n10583;
  assign n12427 = ~n8958 | ~n12651;
  assign n13114 = ~n9560 & ~n13251;
  assign n8035 = ~n8145 | ~n8092;
  assign n11547 = ~n11557 & ~n11579;
  assign n10493 = ~n10496 & ~n11480;
  assign n8047 = ~n8045 | ~n8044;
  assign n13118 = ~n13507 | ~n13521;
  assign n12667 = ~n12028 & ~n12721;
  assign n8157 = ~n8145 | ~n9633;
  assign n12705 = ~REIP_REG_16__SCAN_IN | ~n12028;
  assign n9344 = ~n13490 & ~n12663;
  assign n13523 = ~n13559 | ~n13521;
  assign n7584 = ~n7627 | ~n12145;
  assign n11966 = ~n12030 & ~n12721;
  assign n10545 = ~n10548 & ~n11480;
  assign n11317 = ~n11325 & ~n11579;
  assign n10305 = ~n8133 | ~n10320;
  assign n12481 = ~n13528 & ~n12663;
  assign n12664 = ~n13329 & ~n12663;
  assign n10676 = ~n10681 & ~n11478;
  assign n10783 = ~n10787 & ~n11480;
  assign n10901 = ~n10681 & ~n10886;
  assign n10681 = ~n11845 | ~n10673;
  assign n7600 = ~n7595 | ~n11813;
  assign n8145 = ~n8030 ^ n8044;
  assign n10548 = ~n10541 & ~n7990;
  assign n7627 = ~n7538 & ~n7537;
  assign n10621 = ~n11845 | ~n10613;
  assign n12030 = ~n11931;
  assign n10320 = ~n8132 | ~n8131;
  assign n12663 = ~n9343 | ~n12718;
  assign n13008 = ~n13490 & ~n13527;
  assign n9778 = ~n9777 | ~n13371;
  assign n10590 = ~n11846;
  assign n12047 = ~n13528 & ~n12045;
  assign n9165 = ~n13507 | ~n12040;
  assign n9588 = ~n9587 | ~n12926;
  assign n10541 = ~n11852 | ~n10484;
  assign n13371 = ~n11324 | ~n13043;
  assign n9775 = ~n13045 & ~n9774;
  assign n13250 = ~n8001 & ~n11324;
  assign n13298 = ~n11326 | ~n13043;
  assign n10523 = ~n10526 & ~n11480;
  assign n9361 = ~n13045 & ~n9367;
  assign n11846 = ~n10582 | ~n7990;
  assign n7577 = ~n10331 | ~n10369;
  assign n10335 = ~n10331 | ~n12691;
  assign n12782 = ~n13490 & ~n12769;
  assign n12765 = ~n13490 & ~n12764;
  assign n11847 = ~n10780 | ~n7990;
  assign n11707 = ~n10642 | ~n10886;
  assign n11931 = ~n12617 | ~n8959;
  assign n12498 = ~n12490 & ~n13490;
  assign n10319 = ~n8129 | ~n8130;
  assign n11316 = ~n13045 & ~n11569;
  assign n12842 = ~n13490 & ~n12841;
  assign n8986 = ~n8985 | ~n8984;
  assign n10526 = ~n10581 & ~n7990;
  assign n7956 = ~n8018;
  assign n11244 = ~n13528 & ~n12769;
  assign n9734 = ~n9733 | ~n9732;
  assign n12926 = ~n11632 | ~n12929;
  assign n11718 = ~n12929 & ~REIP_REG_1__SCAN_IN;
  assign n12040 = ~n9164 & ~n9339;
  assign n10989 = ~n13528 & ~n12490;
  assign n9191 = ~n13315 & ~n13333;
  assign n9174 = ~n9173 | ~n9172;
  assign n13071 = ~n13333 & ~n13234;
  assign n10642 = ~n10779 & ~n7990;
  assign n7983 = ~n7982 | ~n7981;
  assign n11594 = ~n13528 & ~n12764;
  assign n11586 = ~n13528 & ~n12841;
  assign n12716 = ~n13333 & ~n12894;
  assign n7593 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n7592;
  assign n12675 = ~n13333 & ~n12868;
  assign n8129 = ~n8102 | ~n9535;
  assign n7555 = ~n7592 & ~n10338;
  assign n10779 = ~n11820 | ~n10636;
  assign n13528 = ~n10928 | ~n13389;
  assign n9321 = ~n13197 | ~n13224;
  assign n9176 = ~n13197 | ~n13154;
  assign n8990 = ~n13197 | ~n13086;
  assign n12417 = ~n12636 | ~n8958;
  assign n8102 = ~n11820 | ~n9633;
  assign n13069 = ~n13334 | ~PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n13029 = ~n13335 | ~EBX_REG_26__SCAN_IN;
  assign n7006 = ~n7231 & ~n11155;
  assign n13210 = ~n13453 | ~n13197;
  assign n12938 = ~n13197 | ~n13352;
  assign n11326 = ~n9125 | ~n13222;
  assign n10321 = ~n10234 | ~n10233;
  assign n12554 = ~n11456 | ~DATAI_2_;
  assign n12369 = ~n11456 | ~DATAI_7_;
  assign n10544 = ~n10542 & ~n7936;
  assign n12358 = ~n11456 | ~DATAI_4_;
  assign n12569 = ~n11456 | ~DATAI_6_;
  assign n12538 = n10499 & n10747;
  assign n12346 = ~n11456 | ~DATAI_3_;
  assign n12312 = ~n11456 | ~DATAI_0_;
  assign n13460 = ~n13453 | ~n13472;
  assign n8484 = ~n13472 | ~n12613;
  assign n10233 = ~n8128 & ~n8127;
  assign n9545 = ~n9544;
  assign n12334 = ~n11456 | ~DATAI_1_;
  assign n8808 = ~n13560 | ~EBX_REG_21__SCAN_IN;
  assign n10234 = ~n8117 | ~n8116;
  assign n11646 = ~n11636;
  assign n12317 = n10574 & n10747;
  assign n7948 = ~n7974;
  assign n13335 = ~n8983 & ~n11636;
  assign n12330 = ~n11627 & ~n10900;
  assign n10442 = ~n13565 & ~n10441;
  assign n11620 = ~n8467 & ~n13391;
  assign n8989 = ~n11632 | ~STATE2_REG_1__SCAN_IN;
  assign n7949 = ~n7975;
  assign n12749 = ~n13467 | ~PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n12994 = ~n13316 & ~n12993;
  assign n9544 = ~n9542 & ~n9541;
  assign n12792 = ~n7008 | ~DATAI_19_;
  assign n12794 = ~n13391 & ~n12790;
  assign n10586 = ~n12588 | ~n12287;
  assign n11422 = ~n12428 & ~n13316;
  assign n11347 = ~n12449 & ~n13316;
  assign n12098 = ~n8533 & ~n13391;
  assign n8426 = ~n13467 | ~PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n13175 = ~n9693 | ~n9692;
  assign n12752 = ~n12741 & ~n13316;
  assign n10447 = ~n13565 & ~n12790;
  assign n8935 = ~n13177 | ~DATAI_6_;
  assign n10425 = ~n13565 & ~n10459;
  assign n12444 = ~n12433 & ~n13316;
  assign n9253 = ~n13177 | ~DATAI_8_;
  assign n10405 = ~n13565 & ~n8377;
  assign n10434 = ~n13565 & ~n10432;
  assign n9305 = ~n13177 | ~DATAI_9_;
  assign n10438 = ~n13565 & ~n8268;
  assign n10413 = ~n13565 & ~n8177;
  assign n10417 = ~n13565 & ~n8148;
  assign n10421 = ~n13565 & ~n11753;
  assign n10203 = ~n10080 | ~n10079;
  assign n12828 = ~n13316 & ~n12827;
  assign n8117 = ~n7990 | ~n9633;
  assign n9082 = ~n13177 | ~DATAI_7_;
  assign n12895 = ~n13316 & ~n12894;
  assign n8794 = ~n13177 | ~DATAI_5_;
  assign n8011 = ~n10224 | ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n10455 = ~n13565 & ~n10454;
  assign n12799 = ~n13391 | ~n10297;
  assign n10409 = ~n13565 & ~n8185;
  assign n10429 = ~n13565 & ~n8119;
  assign n8014 = ~n10224 & ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n10450 = ~n13565 & ~n8467;
  assign n10401 = ~n13565 & ~n10399;
  assign n11767 = ~n12616 & ~n13316;
  assign n12869 = ~n13316 & ~n12868;
  assign n7947 = ~n10616 & ~STATE2_REG_0__SCAN_IN;
  assign n7990 = ~n7989 ^ n7988;
  assign n9108 = ~n9106 | ~n9105;
  assign n11481 = ~n12588 | ~n10616;
  assign n7422 = ~n8804 | ~n7421;
  assign n11632 = ~n8953 | ~n8952;
  assign n10402 = ~n13566 | ~DATAI_1_;
  assign n10215 = ~n8126 | ~n7017;
  assign n10426 = ~n13566 | ~DATAI_6_;
  assign n10414 = ~n13566 | ~DATAI_7_;
  assign n10410 = ~n13566 | ~DATAI_8_;
  assign n10435 = ~n13566 | ~DATAI_5_;
  assign n10430 = ~n13566 | ~DATAI_0_;
  assign n13091 = ~n9706 & ~n9705;
  assign n10439 = ~n13566 | ~DATAI_10_;
  assign n10418 = ~n13566 | ~DATAI_4_;
  assign n9693 = ~n13453 | ~n9698;
  assign n10422 = ~n13566 | ~DATAI_13_;
  assign n10406 = ~n13566 | ~DATAI_12_;
  assign n9105 = ~n9104 | ~n9103;
  assign n10616 = ~n7590 | ~n7543;
  assign n8126 = ~n10213 | ~STATE2_REG_2__SCAN_IN;
  assign n13164 = ~n13465 | ~n7666;
  assign n7955 = ~n12588 | ~n10490;
  assign n7543 = ~n7542 | ~n7541;
  assign n9106 = ~n9099 & ~n9098;
  assign n9537 = ~n9548 & ~n9789;
  assign n12960 = ~n9498 & ~n9497;
  assign n11830 = ~n10886 & ~n11480;
  assign n12588 = n7590 ^ n7589;
  assign n7591 = ~n7590 & ~n7589;
  assign n10488 = ~STATE2_REG_3__SCAN_IN | ~n7650;
  assign n7987 = ~n7941 | ~n7940;
  assign n12900 = ~n9456 & ~n9455;
  assign n7941 = ~n7936 | ~n10490;
  assign n8127 = ~n7017 & ~n9698;
  assign n9098 = ~n10033 & ~n9097;
  assign n9704 = ~n9536 | ~PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n7542 = ~n7539;
  assign n9079 = ~n9076 | ~n9075;
  assign n7539 = ~n7490 | ~n7557;
  assign n7936 = n7560 ^ n7559;
  assign n7486 = ~n7559;
  assign n11553 = ~n12208 | ~n12207;
  assign n9071 = ~n9698 | ~n13315;
  assign n7557 = ~n7489 | ~n7488;
  assign n8999 = ~n8931 | ~n8930;
  assign n8931 = ~n13224 | ~n9698;
  assign n8495 = ~n8494 | ~n8493;
  assign n8709 = ~n12699;
  assign n8932 = ~n8790 | ~n8789;
  assign n11402 = ~n10857 | ~n10856;
  assign n7505 = ~n7496 & ~n8135;
  assign n7489 = ~n7479 | ~n7478;
  assign n12699 = ~n8708 | ~n8707;
  assign n12654 = n8669 & n8668;
  assign n8790 = ~n13154 | ~n9698;
  assign n7377 = ~n7375 | ~n7374;
  assign n11319 = ~n10468 | ~n10467;
  assign n10038 = ~n10035 | ~n10032;
  assign n7495 = ~n7453 | ~n7480;
  assign n8750 = ~n13086 | ~n9698;
  assign n7392 = ~n7322 & ~n7321;
  assign n9101 = ~n8948 | ~n12680;
  assign n8708 = ~n12917 | ~n9698;
  assign n9114 = ~n7514 | ~n7513;
  assign n10035 = ~n8948 | ~n8947;
  assign n7475 = ~n7463 | ~n7462;
  assign n7463 = ~n7458 | ~n9092;
  assign n8824 = ~n10938 & ~n10937;
  assign n8073 = ~n8061 & ~n10240;
  assign n8581 = ~n8575 | ~n9696;
  assign n8664 = ~n9698 | ~n12993;
  assign n8630 = ~n8622 | ~n9696;
  assign n9247 = ~n9241 | ~n9696;
  assign n10938 = ~n8822 | ~n8821;
  assign n7379 = ~n7341 & ~n7340;
  assign n7452 = ~n9135 | ~n7451;
  assign n8947 = ~n8946 & ~n10074;
  assign n8626 = ~n12894 | ~n9698;
  assign n7458 = ~n7506 & ~n9110;
  assign n7416 = ~n8946;
  assign n8583 = ~n8541 | ~n9698;
  assign n7970 = ~n7888 & ~n10240;
  assign n7407 = ~n7405 & ~n7404;
  assign n9097 = ~n9096 | ~n9102;
  assign n7386 = ~n7406 | ~n7966;
  assign n7446 = ~n7445 & ~n10490;
  assign n11023 = ~n8345 & ~n8344;
  assign n9135 = ~n10391 & ~n7448;
  assign n7940 = ~n7939 & ~n7938;
  assign n7986 = ~n7934 | ~n7933;
  assign n9134 = ~n7624 | ~n10499;
  assign n7473 = ~n7468 & ~n10245;
  assign n12025 = ~n8538 | ~n8537;
  assign n10032 = ~n9091 | ~n8950;
  assign n8538 = ~n12827 | ~n9698;
  assign n7361 = ~n7354 | ~n7388;
  assign n7946 = ~n7945 | ~n7944;
  assign n7406 = ~n7385 | ~n7384;
  assign n7934 = ~n7937 | ~n8065;
  assign n11239 = ~n8384 | ~n8383;
  assign n7339 = ~n7401 | ~n8068;
  assign n8499 = ~n8473 | ~n8472;
  assign n7994 = ~n7993 | ~n7992;
  assign n7451 = ~n9156 | ~n7450;
  assign n8822 = ~n8818 | ~n8819;
  assign n9095 = ~n9091 | ~n9090;
  assign n10391 = ~n7408 & ~n7601;
  assign n7412 = ~n7411 | ~n10515;
  assign n7376 = ~n7404 | ~n7966;
  assign n7347 = ~n7966 | ~n7356;
  assign n7444 = ~n7440 | ~n7439;
  assign n8818 = ~n8813 ^ n10045;
  assign n7466 = ~n7443 | ~n7442;
  assign n7958 = ~n8031 | ~n7966;
  assign n7462 = ~n7461 | ~n10574;
  assign n7352 = ~n7350 | ~n10499;
  assign n9156 = ~n8949 & ~n10240;
  assign n7483 = ~n9131 & ~n10490;
  assign n7418 = ~n7471 | ~n7230;
  assign n7359 = ~n7357 & ~n7356;
  assign n7408 = ~n7397 | ~n9093;
  assign n7937 = ~n7931 & ~n7930;
  assign n7354 = ~n7966 | ~n7358;
  assign n7364 = ~n7388 | ~n7353;
  assign n8140 = ~n8136 & ~n8135;
  assign n8121 = ~n8136 & ~n8118;
  assign n7945 = ~n7943 | ~n7966;
  assign n7967 = ~n8068 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n8069 = ~n8068 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n7439 = ~n7438 & ~n7437;
  assign n8471 = ~n8193 & ~n8466;
  assign n8153 = ~n8147 | ~INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n8536 = ~n8193 & ~n8532;
  assign n8802 = ~n8492 & ~n8491;
  assign n7963 = ~n8042 & ~n7959;
  assign n7351 = ~n7959 & ~n10245;
  assign n7336 = ~n7959 | ~n8092;
  assign n9094 = ~n9093 & ~n9092;
  assign n7230 = ~n7441 | ~n10574;
  assign n7425 = ~n7518;
  assign n8380 = ~n8193 & ~n8376;
  assign n8539 = ~n8501 | ~PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n9117 = ~n7519 & ~n7518;
  assign n7344 = ~n7403 & ~n8068;
  assign n7938 = ~n7959 & ~n8003;
  assign n8419 = ~n11939 & ~n9789;
  assign n7350 = ~n8068 | ~n7400;
  assign n7957 = ~n8068 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n7953 = ~n7950 & ~n7959;
  assign n7944 = ~n8068 | ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n7343 = n7403 & n7959;
  assign n7357 = ~n7932 & ~n7355;
  assign n8114 = ~n8113 | ~n8112;
  assign n8852 = ~n10932 | ~EBX_REG_11__SCAN_IN;
  assign n8843 = ~n10932 | ~EBX_REG_8__SCAN_IN;
  assign n7952 = ~n7961 & ~n7951;
  assign n8879 = ~n10932 | ~EBX_REG_20__SCAN_IN;
  assign n8861 = ~n10932 | ~EBX_REG_14__SCAN_IN;
  assign n8828 = ~n10932 | ~EBX_REG_3__SCAN_IN;
  assign n8882 = ~n10932 | ~EBX_REG_21__SCAN_IN;
  assign n8837 = ~n10932 | ~EBX_REG_6__SCAN_IN;
  assign n7962 = ~n7961 & ~n7960;
  assign n8864 = ~n10932 | ~EBX_REG_15__SCAN_IN;
  assign n7199 = ~n7465 | ~n8498;
  assign n8147 = ~n8796 & ~n11497;
  assign n8870 = ~n10932 | ~EBX_REG_17__SCAN_IN;
  assign n7319 = ~n7318 & ~n7317;
  assign n7482 = ~n8796 & ~n7601;
  assign n8383 = ~n12741 | ~n9698;
  assign n7931 = ~n7961 & ~n8586;
  assign n7443 = ~n7413 | ~n7231;
  assign n8873 = ~n10932 | ~EBX_REG_18__SCAN_IN;
  assign n8834 = ~n10932 | ~EBX_REG_5__SCAN_IN;
  assign n8846 = ~n10932 | ~EBX_REG_9__SCAN_IN;
  assign n8867 = ~n10932 | ~EBX_REG_16__SCAN_IN;
  assign n8855 = ~n10932 | ~EBX_REG_12__SCAN_IN;
  assign n8811 = ~n10932 | ~EBX_REG_1__SCAN_IN;
  assign n7460 = ~n8008 | ~n7231;
  assign n8831 = ~n10932 | ~EBX_REG_4__SCAN_IN;
  assign n8138 = ~n9707 | ~EAX_REG_3__SCAN_IN;
  assign n7311 = ~n7394 | ~n8488;
  assign n7518 = ~n7315 | ~n7413;
  assign n8169 = ~n9707 | ~EAX_REG_6__SCAN_IN;
  assign n8849 = ~n10932 | ~EBX_REG_10__SCAN_IN;
  assign n8858 = ~n10932 | ~EBX_REG_13__SCAN_IN;
  assign n8840 = ~n10932 | ~EBX_REG_7__SCAN_IN;
  assign n7438 = ~n8008 | ~n10574;
  assign n10241 = ~n10240 | ~READY_N;
  assign n8876 = ~n10932 | ~EBX_REG_19__SCAN_IN;
  assign n8080 = ~n10240 & ~n8079;
  assign n7467 = ~n7465 | ~n7464;
  assign n8416 = n8415 & n9633;
  assign n8151 = ~n9686 & ~n8148;
  assign n8489 = ~n8488;
  assign n7615 = ~n7614 & ~n7613;
  assign n8435 = ~n8381 | ~PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n8060 = ~n8058;
  assign n9074 = ~n9686 & ~n9069;
  assign n8490 = ~n8791 & ~n9132;
  assign n8535 = ~n9686 & ~n8533;
  assign n8703 = ~n9686 & ~n12790;
  assign n8746 = ~n9686 & ~n8743;
  assign n9259 = ~n9210 | ~n9209;
  assign n8667 = ~n9686 & ~n8662;
  assign n8179 = ~n9686 & ~n8177;
  assign n7481 = ~n8488 & ~n10499;
  assign n8188 = ~n9686 & ~n8185;
  assign n8066 = ~n8065 & ~n8079;
  assign n8108 = ~n9686 & ~n8103;
  assign n8579 = ~n9686 & ~n8576;
  assign n7312 = ~n7613 | ~n10574;
  assign n8379 = ~n9686 & ~n8377;
  assign n7923 = ~n7921 | ~n9132;
  assign n8161 = ~n9686 & ~n10432;
  assign n7320 = ~n8801 | ~n12680;
  assign n7856 = ~n8031;
  assign n8786 = ~n9686 & ~n8783;
  assign n7429 = ~n8792 & ~n11156;
  assign n7413 = ~n8498;
  assign n8470 = ~n9686 & ~n8467;
  assign n8120 = ~n9686 & ~n8119;
  assign n8628 = ~n9686 & ~n8623;
  assign n7317 = ~n8792 | ~n11156;
  assign n7427 = ~n9132 | ~n11156;
  assign n7961 = ~n7337 | ~n9132;
  assign n7925 = ~n7924 & ~n10490;
  assign n8271 = ~n9686 & ~n8268;
  assign n8841 = ~n10937 | ~INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n8829 = ~n10937 | ~INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n9210 = ~n9029 | ~n9028;
  assign n8816 = ~n8815 & ~n8814;
  assign n8853 = ~n10937 | ~INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n8856 = ~n10937 | ~INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n7459 = ~n10515 | ~n9102;
  assign n8950 = ~n9092 & ~n10074;
  assign n8859 = ~n10937 | ~INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n8835 = ~n10937 | ~INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n8850 = ~n10937 | ~INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n8817 = ~n9723 & ~EBX_REG_0__SCAN_IN;
  assign n7613 = ~n8814 | ~n9102;
  assign n8192 = ~n10574 | ~n7231;
  assign n8101 = ~n11156;
  assign n8810 = ~n10574 | ~n10748;
  assign n8575 = ~n8573 | ~n8572;
  assign n7924 = ~n10574 & ~n8004;
  assign n8868 = ~n10937 | ~INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n8381 = ~n8343 & ~n7671;
  assign n11637 = ~n10574 & ~n10245;
  assign n8792 = ~n10499;
  assign n8838 = ~n10937 | ~INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n8832 = ~n10937 | ~INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n9686 = ~n13389 | ~STATE2_REG_2__SCAN_IN;
  assign n8826 = ~n10937 | ~INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n7922 = ~n7231 | ~n8079;
  assign n8031 = ~n7733 | ~n7732;
  assign n8847 = ~n10937 | ~INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n8273 = ~n12433 | ~n9698;
  assign n7345 = ~n10245 | ~n10499;
  assign n8862 = ~n10937 | ~INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n8801 = ~n10937;
  assign n8865 = ~n10937 | ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n7996 = ~n10748 & ~n10574;
  assign n7887 = ~n8042;
  assign n8844 = ~n10937 | ~INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n8815 = ~n10574 | ~EBX_REG_0__SCAN_IN;
  assign n8343 = ~n8267 | ~PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n8042 = ~n7886 & ~n7885;
  assign n7921 = ~n10574 | ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n11156 = ~n7087 & ~n7086;
  assign n8265 = ~n12390 & ~n9789;
  assign n10499 = ~n7057 | ~n7056;
  assign n7231 = ~n7229 & ~n7228;
  assign n8003 = ~n7853 & ~n7852;
  assign n8225 = ~n8221 | ~n8220;
  assign n7261 = ~n7245 | ~n7244;
  assign n7057 = n7031 & n7030;
  assign n10574 = ~n7198 | ~n7197;
  assign n8190 = ~n12616 | ~n9698;
  assign n8304 = ~n8288 | ~n8287;
  assign n7260 = ~n7259 | ~n7258;
  assign n7331 = ~n7342 | ~n10637;
  assign n8338 = ~n8337 | ~n8336;
  assign n8303 = ~n8302 | ~n8301;
  assign n7114 = ~n7113 & ~n7112;
  assign n7198 = ~n7178 & ~n7177;
  assign n7115 = ~n7107 & ~n7106;
  assign n7031 = ~n7023 & ~n7022;
  assign n7071 = ~n7063 & ~n7062;
  assign n8181 = ~n12428 | ~n9698;
  assign n7101 = ~n7093 & ~n7092;
  assign n7070 = ~n7069 & ~n7068;
  assign n7085 = ~n7077 & ~n7076;
  assign n7030 = ~n7029 & ~n7028;
  assign n7197 = ~n7196 & ~n7195;
  assign n7084 = ~n7083 & ~n7082;
  assign n7100 = ~n7099 & ~n7098;
  assign n7178 = ~n7168 | ~n7167;
  assign n7205 = ~n7201 | ~n7200;
  assign n7210 = ~n7209 | ~n7208;
  assign n12347 = ~n13463 | ~DATAI_27_;
  assign n8171 = n12449 & n9698;
  assign n7204 = ~n7203 | ~n7202;
  assign n7055 = ~n7042 | ~n7041;
  assign n7211 = ~n7207 | ~n7206;
  assign n12345 = ~n13463 | ~DATAI_19_;
  assign n7112 = ~n7111 | ~n7110;
  assign n12359 = ~n13463 | ~DATAI_28_;
  assign n7157 = ~n7146 | ~n7145;
  assign n7136 = ~n7135 | ~n7134;
  assign n12313 = ~n13463 | ~DATAI_16_;
  assign n7092 = ~n7091 | ~n7090;
  assign n7225 = ~n7221 | ~n7220;
  assign n12301 = ~n13463 | ~DATAI_24_;
  assign n7098 = ~n7097 | ~n7096;
  assign n7224 = ~n7223 | ~n7222;
  assign n7107 = ~n7103 | ~n7102;
  assign n12333 = ~n13463 | ~DATAI_25_;
  assign n12335 = ~n13463 | ~DATAI_17_;
  assign n7218 = ~n7217 | ~n7216;
  assign n7023 = ~n7019 | ~n7018;
  assign n7099 = ~n7095 | ~n7094;
  assign n7022 = ~n7021 | ~n7020;
  assign n7082 = ~n7081 | ~n7080;
  assign n7029 = ~n7025 | ~n7024;
  assign n7083 = ~n7079 | ~n7078;
  assign n7106 = ~n7105 | ~n7104;
  assign n12549 = ~n13463 | ~DATAI_18_;
  assign n7028 = ~n7027 | ~n7026;
  assign n7219 = ~n7215 | ~n7214;
  assign n7195 = ~n7194 | ~n7193;
  assign n12555 = ~n13463 | ~DATAI_26_;
  assign n7076 = ~n7075 | ~n7074;
  assign n12560 = ~n13463 | ~DATAI_30_;
  assign n7242 = ~n7241 | ~n7240;
  assign n7063 = ~n7059 | ~n7058;
  assign n12368 = ~n13463 | ~DATAI_31_;
  assign n7250 = ~n7249 | ~n7248;
  assign n7308 = ~n7296 | ~n7295;
  assign n7283 = ~n7282 | ~n7281;
  assign n12544 = ~n13463 | ~DATAI_29_;
  assign n12570 = ~n13463 | ~DATAI_22_;
  assign n12357 = ~n13463 | ~DATAI_20_;
  assign n12536 = ~n13463 | ~DATAI_21_;
  assign n12370 = ~n13463 | ~DATAI_23_;
  assign n7069 = ~n7065 | ~n7064;
  assign n7068 = ~n7067 | ~n7066;
  assign n7194 = ~n7190 & ~n7189;
  assign n7186 = ~n7185 & ~n7184;
  assign n7168 = ~n7163 & ~n7162;
  assign n7111 = ~n9522 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n7187 = ~n7182 & ~n7181;
  assign n12754 = ~n12519 | ~n12774;
  assign n7109 = ~n9648 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n7104 = ~n9673 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n7674 = ~n9647 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n7175 = ~n7174 & ~n7173;
  assign n7110 = ~n9647 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n7072 = ~n9648 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n7176 = ~n7172 & ~n7171;
  assign n7074 = ~n9610 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n7108 = ~n9636 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n8163 = ~n12634 | ~n9698;
  assign n7167 = ~n7166 & ~n7165;
  assign n7089 = ~n9672 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n7065 = ~n9599 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n7154 = ~n7153 & ~n7152;
  assign n7155 = ~n7150 & ~n7149;
  assign n7091 = ~n9656 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n7145 = ~n7144 & ~n7143;
  assign n7060 = ~n9672 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n7146 = ~n7140 & ~n7139;
  assign n7080 = ~n9657 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n7067 = ~n9656 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n7061 = ~n9636 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n7134 = ~n7133 & ~n7132;
  assign n7090 = ~n7003 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n7135 = ~n7130 & ~n7129;
  assign n7058 = ~n9602 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n7066 = ~n9647 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n7059 = ~n9665 | ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n8953 = ~n12690 & ~n8943;
  assign n7126 = ~n7125 & ~n7124;
  assign n7081 = ~n9522 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n7127 = ~n7121 & ~n7120;
  assign n7102 = ~n9653 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n7078 = ~n9673 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n7193 = ~n7192 & ~n7191;
  assign n7079 = ~n9501 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n7795 = ~n9648 | ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n7911 = ~n9657 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n7912 = ~n9610 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n7794 = ~n9636 | ~INSTQUEUE_REG_3__0__SCAN_IN;
  assign n7846 = ~n9657 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n7847 = ~n9522 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n7844 = ~n9647 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n7845 = ~n9656 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n7840 = ~n9610 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n7841 = ~n9602 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n7838 = ~n9599 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n7839 = ~n9648 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n7832 = ~n9673 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n7830 = ~n9653 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n7826 = ~n9672 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n7827 = ~n9665 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n7201 = ~n9665 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n7200 = ~n9599 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n7203 = ~n9636 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n7824 = ~n9501 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n7726 = ~n9602 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n7206 = ~n9653 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n7727 = ~n9656 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n7825 = ~n9636 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n7724 = ~n9653 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n7725 = ~n9657 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n7816 = ~n7003 | ~INSTQUEUE_REG_0__0__SCAN_IN;
  assign n7817 = ~n9673 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n7814 = ~n9610 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n7815 = ~n9656 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n7808 = ~n9602 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n7809 = ~n9501 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n7802 = ~n9647 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n7803 = ~n9522 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n7800 = ~n9665 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n7796 = ~n9672 | ~INSTQUEUE_REG_6__0__SCAN_IN;
  assign n7797 = ~n9599 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n7209 = ~n9648 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n7736 = ~n9636 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n7873 = ~n9602 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n7878 = ~n9648 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n7874 = ~n9522 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n7735 = ~n9501 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n7249 = ~n9602 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n7773 = ~n9599 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n7770 = ~n9665 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n7877 = ~n9653 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n7737 = ~n9522 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n7771 = ~n9501 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n7740 = ~n9653 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n7248 = ~n9610 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n7743 = ~n9610 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n7880 = ~n9599 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n7871 = ~n9647 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n7742 = ~n9648 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n7027 = ~n9647 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n7879 = ~n9673 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n7872 = ~n9656 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n7024 = ~n9522 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n7025 = ~n9672 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n7749 = ~n9656 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n7766 = ~n9522 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n7748 = ~n9673 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n7246 = ~n9599 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n7020 = ~n9610 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n7767 = ~n9656 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n7021 = ~n9636 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n7866 = ~n9610 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n7253 = ~n9656 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n7019 = ~n9648 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n7255 = ~n9522 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n7222 = ~n9647 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n7863 = ~n9672 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n7751 = ~n9602 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n7864 = ~n9501 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n7750 = ~n9647 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n7686 = ~n9665 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n7223 = ~n9522 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n7254 = ~n9647 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n7859 = ~n9636 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n7755 = ~n9665 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n7860 = ~n9665 | ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n7858 = ~n7003 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n7754 = ~n9672 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n7684 = ~n9653 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n7220 = ~n9673 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n7757 = ~n9599 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n7772 = ~n9636 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n7756 = ~n9657 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n7764 = ~n9673 | ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n7238 = ~n9672 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n7685 = ~n9599 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n7232 = ~n9501 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n7716 = ~n9636 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n7221 = ~n9672 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n7208 = ~n9610 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n7765 = ~n9672 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n7681 = ~n9610 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n7235 = ~n9665 | ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n7705 = ~n9647 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n7785 = ~n9648 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n7704 = ~n9648 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n7217 = ~n9656 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n7241 = ~n9673 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n7673 = ~n9602 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n7787 = ~n9653 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n7215 = ~n9501 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n7707 = ~n9501 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n7780 = ~n9647 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n7706 = ~n9610 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n7781 = ~n9602 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n7240 = ~n9657 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n7214 = ~n9602 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n7786 = ~n7003 | ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n7784 = ~n9610 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n7778 = ~n9607 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n7190 = ~n9051 & ~n7188;
  assign n12511 = ~n13491 | ~REIP_REG_11__SCAN_IN;
  assign n7150 = ~n9051 & ~n7147;
  assign n7779 = ~n9662 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n7741 = ~n9607 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n7734 = ~n9662 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n7144 = ~n9057 & ~n7141;
  assign n7185 = ~n9057 & ~n9050;
  assign n12991 = ~n13491 | ~REIP_REG_18__SCAN_IN;
  assign n7002 = ~n9057;
  assign n7207 = ~n9662 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n7710 = ~n9607 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n7216 = ~n9607 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n7865 = ~n9662 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n13451 = ~n10063 | ~n11849;
  assign n7857 = ~n9607 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n7801 = ~n9662 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n7252 = ~n9607 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n7676 = ~n8591 & ~n7675;
  assign n7677 = ~n9057 & ~n9641;
  assign n7294 = ~n9057 & ~n7291;
  assign n7301 = ~n9051 & ~n7297;
  assign n8178 = ~n9535 & ~n12415;
  assign n7833 = ~n9607 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n7831 = ~n9662 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n7073 = ~n9662 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n7075 = ~n9607 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n8160 = ~n9535 & ~n12638;
  assign n7088 = ~n9607 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n8155 = ~n11645 & ~n9789;
  assign n7095 = ~n9662 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n13057 = ~n13491 | ~REIP_REG_19__SCAN_IN;
  assign n13306 = ~n13491 | ~REIP_REG_29__SCAN_IN;
  assign n13382 = ~n13491 | ~REIP_REG_21__SCAN_IN;
  assign n9766 = ~n13491 | ~REIP_REG_28__SCAN_IN;
  assign n12866 = ~n13491 | ~REIP_REG_16__SCAN_IN;
  assign n12840 = ~n13491 | ~REIP_REG_14__SCAN_IN;
  assign n12779 = ~n13491 | ~REIP_REG_12__SCAN_IN;
  assign n13456 = ~n13491 | ~REIP_REG_30__SCAN_IN;
  assign n13363 = ~n13491 | ~REIP_REG_27__SCAN_IN;
  assign n12762 = ~n13491 | ~REIP_REG_13__SCAN_IN;
  assign n12826 = ~n13491 | ~REIP_REG_15__SCAN_IN;
  assign n13508 = ~n13491 | ~REIP_REG_25__SCAN_IN;
  assign n13006 = ~n13491 | ~REIP_REG_17__SCAN_IN;
  assign n13262 = ~n13491 | ~REIP_REG_20__SCAN_IN;
  assign n13162 = ~n13491 | ~REIP_REG_26__SCAN_IN;
  assign n8585 = ~n7032 | ~n7048;
  assign n7286 = ~n7526 | ~n7043;
  assign n7288 = ~n7526 | ~n7637;
  assign n8195 = ~n7526 | ~n7032;
  assign n9057 = ~n7631 | ~n10374;
  assign n7324 = ~n10374 & ~n7323;
  assign n8196 = ~n7043 | ~n7521;
  assign n7454 = ~n9787 | ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n11849 = ~n11809;
  assign n7299 = ~n7048 | ~n7637;
  assign n8262 = ~n9708 | ~PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n7470 = ~n7469 & ~n10490;
  assign n7491 = ~n9787 & ~n10637;
  assign n8168 = ~n9708 | ~PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n8307 = ~n9708 | ~PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n8142 = ~n12575 | ~n9698;
  assign n7476 = ~n9787 & ~n10638;
  assign n9855 = ~n7449 & ~STATE_REG_0__SCAN_IN;
  assign n7338 = ~n10490 | ~INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n7498 = ~n10637 & ~n7497;
  assign n8551 = ~n7521 | ~n7637;
  assign n7032 = ~n8111 & ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n7526 = ~n8135 & ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n12835 = ~INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n12680 = ~READY_N;
  assign n11893 = ~INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n10341 = ~INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n7003 = ~n9057;
  assign n10223 = ~n7990 | ~n8092;
  assign n8061 = n8079 ^ n8081;
  assign n7391 = n7387 & n7386;
  assign n12718 = ~n9339 | ~n9340;
  assign n10934 = ~n8819;
  assign n9140 = ~n9139 | ~n9138;
  assign n9138 = ~n9137 & ~n9136;
  assign n11896 = ~INSTADDRPOINTER_REG_8__SCAN_IN | ~n11895;
  assign n7358 = ~INSTQUEUERD_ADDR_REG_0__SCAN_IN ^ INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n8194 = ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n7170 = ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n7038 = ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n7034 = ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n7268 = ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n7263 = ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n7602 = ~n8948;
  assign n7123 = ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n7119 = ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n7888 = n8058 ^ n8059;
  assign n7928 = ~n9132 & ~n10490;
  assign n7594 = ~n11638 | ~n10391;
  assign n7580 = ~n7579 | ~n7578;
  assign n7579 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n7576;
  assign n9172 = ~n13335 | ~EBX_REG_21__SCAN_IN;
  assign n8984 = ~n13335 | ~EBX_REG_20__SCAN_IN;
  assign n12576 = ~PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n8823 = ~n8822;
  assign n8107 = ~n8106 | ~n8105;
  assign n9303 = ~n9251 & ~n9250;
  assign n12696 = ~n12734 | ~n12733;
  assign n12734 = ~n12718 & ~n12717;
  assign n8095 = ~n8094;
  assign n8086 = ~n8085;
  assign n8078 = ~n8077;
  assign n7589 = ~n7505 & ~n7504;
  assign n11444 = ~n11699;
  assign n10690 = ~n10684 | ~n10678;
  assign n12145 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n8814 = ~n7310 | ~n7309;
  assign n9318 = ~n13334 | ~PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n12033 = ~n12667 | ~n12032;
  assign n12726 = ~n12805;
  assign n13196 = ~n13400;
  assign n9316 = ~n8886 & ~n8885;
  assign n9339 = ~n9163 & ~n9162;
  assign n9340 = n8869 ^ n10045;
  assign n11589 = ~n11591 & ~n11590;
  assign n11087 = ~n10987 | ~n10986;
  assign n8807 = ~n13150;
  assign n7322 = ~n9139;
  assign n13079 = ~n13078;
  assign n12912 = ~n9567 & ~n9566;
  assign n9332 = ~n12888;
  assign n11940 = ~n8423 ^ n8430;
  assign n13405 = ~n13434 ^ INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n13521 = n12734 ^ n12733;
  assign n12524 = ~n13377;
  assign n12624 = ~n12623 | ~n12622;
  assign n12459 = ~n12458 | ~n12457;
  assign n12646 = ~n13335 | ~EBX_REG_5__SCAN_IN;
  assign n11653 = ~n11644 | ~n11643;
  assign n11656 = ~n11655 | ~n11654;
  assign n11648 = ~n11647 | ~n11646;
  assign n12295 = ~n12294 | ~n12293;
  assign n11957 = ~n11956 | ~n11955;
  assign n12859 = ~n13319;
  assign n12853 = ~n13227;
  assign n12913 = ~n12700 ^ n12699;
  assign n11088 = ~n13559 | ~n12509;
  assign n10867 = ~n13559 | ~n12381;
  assign n13536 = ~n13559 | ~n13534;
  assign n10667 = ~n10666 | ~n10665;
  assign n10668 = ~n10825;
  assign n13542 = ~n13559 | ~n13540;
  assign n10470 = ~n13559 | ~n12286;
  assign n9308 = ~n7008 | ~DATAI_25_;
  assign n9256 = ~n7008 | ~DATAI_24_;
  assign n9085 = ~n7008 | ~DATAI_23_;
  assign n8938 = ~n7008 | ~DATAI_22_;
  assign n8798 = ~n7008 | ~DATAI_21_;
  assign n12658 = ~n7008 | ~DATAI_18_;
  assign n12297 = n10322 ^ n10321;
  assign n10322 = ~n10320 | ~n10319;
  assign n13152 = n13467 & PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n12473 = n11024 ^ n11023;
  assign n12391 = n10826 ^ n10821;
  assign n11649 = n10313 ^ n10312;
  assign n9758 = ~n13501;
  assign n9363 = ~n13299;
  assign n13376 = ~n13372 | ~n13371;
  assign n13375 = ~n13374 | ~n13373;
  assign n13380 = ~n13487 | ~n13370;
  assign n13259 = ~n13258 | ~n13257;
  assign n13258 = ~n13256 | ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n13004 = ~n13110 | ~INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n12758 = ~n12757 | ~n12756;
  assign n12760 = ~n12833 | ~n12835;
  assign n9160 = ~n9159 | ~n9158;
  assign n12510 = ~n12509 | ~n13507;
  assign n12515 = ~n12773 | ~n12770;
  assign n11892 = ~INSTADDRPOINTER_REG_7__SCAN_IN | ~n11919;
  assign n11890 = ~n11889 | ~n11888;
  assign n11561 = ~n11560 | ~n11559;
  assign n11560 = ~n11557 | ~n13371;
  assign n11559 = ~n13374 | ~n11558;
  assign n9116 = ~n13043;
  assign n11576 = ~n11575 | ~n11574;
  assign n11395 = ~n8001 | ~n13299;
  assign n12114 = ~n12113 | ~n12112;
  assign n12106 = ~n12105 | ~n12104;
  assign n12122 = ~n12121 | ~n12120;
  assign n12134 = ~n12133 | ~n12132;
  assign n12320 = ~n12319 | ~n12318;
  assign n12341 = ~n12340 | ~n12339;
  assign n12353 = ~n12352 | ~n12351;
  assign n12364 = ~n12363 | ~n12362;
  assign n12375 = ~n12374 | ~n12373;
  assign n11454 = ~n11453 | ~n11452;
  assign n11470 = ~n11469 | ~n11468;
  assign n12255 = ~n12254 | ~n12253;
  assign n12263 = ~n12262 | ~n12261;
  assign n12274 = ~n12273 | ~n12272;
  assign n11380 = ~n11379 | ~n11378;
  assign n11868 = ~n11867 | ~n11866;
  assign n11880 = ~n11879 | ~n11878;
  assign n12219 = ~n12218 | ~n12217;
  assign n12246 = ~n12245 | ~n12244;
  assign n12227 = ~n12226 | ~n12225;
  assign n12235 = ~n12234 | ~n12233;
  assign n7355 = ~n10499 | ~n10574;
  assign n9641 = ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n7690 = ~n9662 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n7691 = ~n9656 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n7693 = ~n9672 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n7692 = ~n9648 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n7687 = ~n9501 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n7675 = ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n7713 = ~n9672 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n7712 = ~n9673 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n7718 = ~n9662 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n7719 = ~n9665 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n7717 = ~n9599 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n7711 = ~n9522 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n7348 = ~n7403;
  assign n8020 = ~n7950;
  assign n9050 = ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n8548 = ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n7960 = ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n8592 = ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n9417 = ~n9290 | ~n9289;
  assign n9209 = ~n9066 | ~n9065;
  assign n8403 = ~n8402 | ~n8401;
  assign n8300 = ~n8296 | ~n8295;
  assign n7976 = ~n7943;
  assign n7450 = ~n7449;
  assign n7469 = ~n12681;
  assign n9052 = ~INSTQUEUE_REG_6__0__SCAN_IN;
  assign n7179 = ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n7180 = ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n8199 = ~INSTQUEUE_REG_4__0__SCAN_IN;
  assign n7188 = ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n7160 = ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n7164 = ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n7161 = ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n7044 = ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n7049 = ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n7285 = ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n7291 = ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n7287 = ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n7298 = ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n7302 = ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n7297 = ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n7273 = ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n7278 = ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n7277 = ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n7274 = ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n7342 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ n7328;
  assign n7372 = n7332 ^ INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n8659 = ~n8658 | ~n8657;
  assign n8660 = ~n8644 | ~n8643;
  assign n9490 = ~PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n8584 = ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n7141 = ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n7142 = ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n7138 = ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n7151 = ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n7147 = ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n8590 = ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n7131 = ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n7128 = ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n9296 = n9291 & n9696;
  assign n8745 = ~n9789 | ~n8744;
  assign n8578 = ~n9789 | ~n8577;
  assign n8465 = ~n8449 | ~n8448;
  assign n8375 = ~n8359 | ~n8358;
  assign n8374 = ~n8373 | ~n8372;
  assign n8235 = ~n8231 | ~n8230;
  assign n8241 = ~n8237 | ~n8236;
  assign n8254 = ~n8253 | ~n8252;
  assign n8255 = ~n8251 | ~n8250;
  assign n8248 = ~n8247 | ~n8246;
  assign n13279 = ~n13271;
  assign n7611 = ~n8192;
  assign n8043 = n8042 ^ n8041;
  assign n8034 = ~n8033 | ~n10076;
  assign n7932 = ~n7928;
  assign n7939 = ~n7937;
  assign n7951 = ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n7501 = ~n9787;
  assign n7496 = ~n7495;
  assign n7500 = ~n7665;
  assign n7409 = ~n10075;
  assign n11441 = n11488 ^ INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n10898 = INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ n7497;
  assign n7169 = ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n7037 = ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n7033 = ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n7266 = ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n7262 = ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n7403 = ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ n7342;
  assign n7404 = n7372 ^ INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n7400 = n7349 ^ n10638;
  assign n9317 = ~n13335 | ~EBX_REG_22__SCAN_IN;
  assign n8434 = ~PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n11717 = ~n11637 | ~n11646;
  assign n9762 = n9720 ^ n10045;
  assign n12874 = n9391 ^ n10045;
  assign n9389 = ~n10932 | ~EBX_REG_24__SCAN_IN;
  assign n8622 = ~n8621 | ~n8620;
  assign n8224 = ~n8223 | ~n8222;
  assign n8207 = ~n8203 | ~n8202;
  assign n8206 = ~n8205 | ~n8204;
  assign n8175 = n8091 ^ n8071;
  assign n8137 = ~n9708 | ~PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n8174 = ~n9633;
  assign n10467 = n8827 ^ n10045;
  assign n9634 = ~n9500 | ~n9499;
  assign n9540 = ~n9707 | ~EAX_REG_28__SCAN_IN;
  assign n7122 = ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n7118 = ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n9548 = PHYADDRPOINTER_REG_28__SCAN_IN ^ n9536;
  assign n9295 = ~n9294 | ~n9293;
  assign n9454 = ~n9449 | ~n9696;
  assign n8969 = ~PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n12707 = ~PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n8339 = ~n8323 | ~n8322;
  assign n8240 = ~n8239 | ~n8238;
  assign n8249 = ~n8245 | ~n8244;
  assign n8013 = ~n10223;
  assign n8136 = ~n8147;
  assign n8113 = ~n9707 | ~EAX_REG_1__SCAN_IN;
  assign n13429 = ~n13434 | ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n13190 = ~n9725 | ~n9724;
  assign n13101 = ~n13186 ^ n9723;
  assign n9198 = ~n9197 ^ n10045;
  assign n9195 = ~n10932 | ~EBX_REG_23__SCAN_IN;
  assign n9315 = n9194 ^ n10045;
  assign n9192 = ~n10932 | ~EBX_REG_22__SCAN_IN;
  assign n12695 = ~n8878 ^ n10045;
  assign n8877 = ~n10937 | ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n12733 = n8875 ^ n10045;
  assign n8874 = ~n10937 | ~INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n9162 = ~n8866 ^ n10045;
  assign n8477 = n9147 ^ INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n12771 = ~INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n11086 = ~n8854 ^ n10045;
  assign n9088 = ~INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n7612 = ~n8796 | ~n10499;
  assign n10864 = ~n8848 ^ n10045;
  assign n11886 = n8845 ^ n10045;
  assign n8057 = ~n8056;
  assign n8075 = ~n8074;
  assign n11552 = ~n8842 ^ n10045;
  assign n12202 = ~INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n12207 = n8839 ^ n10045;
  assign n11401 = ~n8836 ^ n10045;
  assign n11318 = ~n8830 ^ n10045;
  assign n7541 = ~n7540;
  assign n10484 = ~n11820;
  assign n12302 = ~n10898 | ~STATE2_REG_2__SCAN_IN;
  assign n7919 = n8079 ^ n8004;
  assign n7583 = n10637 & n7628;
  assign n8980 = ~n8963;
  assign n8945 = ~n8944;
  assign n10043 = ~n10039 | ~n7608;
  assign n9732 = ~n13335 | ~EBX_REG_31__SCAN_IN;
  assign n8988 = PHYADDRPOINTER_REG_31__SCAN_IN ^ n8972;
  assign n13338 = ~n13337 | ~n13336;
  assign n13136 = ~n13135 | ~n13134;
  assign n13064 = ~EBX_REG_27__SCAN_IN | ~n13335;
  assign n12970 = ~n9717 ^ n10045;
  assign n9717 = ~n9716 | ~n9715;
  assign n12973 = ~n9761;
  assign n9713 = n9397 ^ n10045;
  assign n9397 = ~n9396 | ~n9395;
  assign n12882 = ~n9394 ^ n10045;
  assign n9392 = ~n10932 | ~EBX_REG_25__SCAN_IN;
  assign n12947 = ~n13335 | ~EBX_REG_25__SCAN_IN;
  assign n12948 = ~n13334 | ~PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n12934 = ~n13335 | ~EBX_REG_24__SCAN_IN;
  assign n12935 = ~n13334 | ~PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n9173 = ~n13334 | ~PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n8985 = ~n13334 | ~PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n12717 = ~n8872 ^ n10045;
  assign n8871 = ~n10937 | ~INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n8960 = ~REIP_REG_15__SCAN_IN | ~n12029;
  assign n12670 = ~n12669 | ~n12668;
  assign n12669 = ~n12667 | ~REIP_REG_16__SCAN_IN;
  assign n12607 = ~n12030 | ~n12029;
  assign n11969 = ~n11968 | ~n11967;
  assign n12448 = ~n12417 | ~n12926;
  assign n12644 = ~n12643 | ~n12642;
  assign n12587 = ~n11717;
  assign n12585 = ~n12584 | ~n12583;
  assign n11948 = ~n10215 | ~n10214;
  assign n9300 = ~n9302;
  assign n8885 = ~n8884 ^ n10045;
  assign n8883 = ~n10937 | ~INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n8966 = n8881 ^ n10045;
  assign n8880 = ~n10937 | ~INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n11584 = n8863 ^ n10045;
  assign n11590 = ~n8860 ^ n10045;
  assign n10986 = n8851 ^ n10045;
  assign n10856 = n8833 ^ n10045;
  assign n8820 = ~n8818;
  assign n10932 = ~n9723 | ~n8810;
  assign n9494 = ~n9493 | ~n9492;
  assign n11752 = ~n11940;
  assign n11647 = ~n7601;
  assign n8487 = ~n9101;
  assign n8131 = ~n8130;
  assign n10297 = ~n8498 | ~n8791;
  assign n13471 = ~n8988;
  assign n9692 = ~n9691 | ~n9690;
  assign n13453 = PHYADDRPOINTER_REG_30__SCAN_IN ^ n9598;
  assign n13332 = PHYADDRPOINTER_REG_29__SCAN_IN ^ n9704;
  assign n13234 = PHYADDRPOINTER_REG_27__SCAN_IN ^ n9496;
  assign n9408 = ~n9407;
  assign n9405 = ~n9404;
  assign n13161 = PHYADDRPOINTER_REG_26__SCAN_IN ^ n9416;
  assign n12951 = PHYADDRPOINTER_REG_25__SCAN_IN ^ n9297;
  assign n13352 = PHYADDRPOINTER_REG_24__SCAN_IN ^ n9208;
  assign n13315 = PHYADDRPOINTER_REG_23__SCAN_IN ^ n9070;
  assign n9077 = ~n9079;
  assign n13224 = PHYADDRPOINTER_REG_22__SCAN_IN ^ n8968;
  assign n9383 = ~n13076;
  assign n13227 = n8934 ^ n8998;
  assign n13150 = n8973 ^ n8932;
  assign n8710 = ~PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n12601 = ~n8500 ^ n8499;
  assign n7671 = ~PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n8382 = ~PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n12463 = ~PHYADDRPOINTER_REG_11__SCAN_IN ^ n8343;
  assign n7670 = ~PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n12390 = ~PHYADDRPOINTER_REG_9__SCAN_IN ^ n8261;
  assign n11645 = PHYADDRPOINTER_REG_4__SCAN_IN ^ n8146;
  assign n10927 = ~n11948;
  assign n13468 = ~n13491 | ~REIP_REG_31__SCAN_IN;
  assign n13400 = n13191 ^ n13190;
  assign n9765 = ~n13131;
  assign n9773 = ~INSTADDRPOINTER_REG_25__SCAN_IN | ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n9366 = ~n13484 | ~n9555;
  assign n9201 = ~n12875;
  assign n13419 = ~n9316 ^ n9315;
  assign n13059 = ~n12696 ^ n12695;
  assign n9375 = ~INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n12844 = ~n9143 ^ n8482;
  assign n12755 = ~n12774 | ~n12520;
  assign n12761 = ~n8478 ^ n8477;
  assign n11237 = n8857 ^ n10045;
  assign n12776 = ~n12746 ^ n12745;
  assign n12509 = n11087 ^ n11086;
  assign n12770 = ~INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n12512 = ~n12469 ^ n12468;
  assign n12468 = ~n12467 | ~n12466;
  assign n12491 = n12438 ^ n12437;
  assign n12437 = ~n12436 | ~n12435;
  assign n8089 = ~n8088;
  assign n7316 = ~n8574;
  assign n7624 = ~n7623;
  assign n11921 = ~REIP_REG_9__SCAN_IN | ~n13491;
  assign n11919 = ~n12514;
  assign n11558 = ~n9119 | ~n11407;
  assign n13374 = ~n13045;
  assign n11397 = ~n11030 | ~n11029;
  assign n11432 = ~INSTADDRPOINTER_REG_4__SCAN_IN | ~INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n11325 = ~INSTADDRPOINTER_REG_2__SCAN_IN | ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n11330 = ~n11329 | ~n11328;
  assign n9126 = ~n11324;
  assign n10582 = ~n10581;
  assign n10372 = ~n10488;
  assign n11638 = n7591 ^ INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n11458 = ~n11457;
  assign n11607 = ~n11496;
  assign n10679 = ~n10692 | ~n10690;
  assign n11376 = ~n10684;
  assign n10902 = ~n10901 | ~n11851;
  assign n10629 = ~n10887;
  assign n10628 = ~n10618 | ~n10617;
  assign n10617 = ~n10677 | ~n7936;
  assign n10057 = ~n10063;
  assign n7648 = ~n12692;
  assign n7449 = n7393 ^ STATE_REG_1__SCAN_IN;
  assign n10039 = ~n10033 | ~n7601;
  assign n13037 = ~n13197 | ~n13161;
  assign n13022 = ~n9714 ^ n9713;
  assign n13506 = n12883 ^ n12882;
  assign n12928 = ~n12931;
  assign n9190 = ~n9189 | ~n9188;
  assign n8962 = ~REIP_REG_20__SCAN_IN | ~n9171;
  assign n12811 = ~REIP_REG_19__SCAN_IN | ~n12810;
  assign n12735 = ~n12944 | ~n13521;
  assign n12725 = ~n12724 | ~n12723;
  assign n13527 = ~n12718 ^ n12717;
  assign n12711 = ~n12710 | ~n12709;
  assign n12035 = ~n12034 | ~n12033;
  assign n12613 = PHYADDRPOINTER_REG_14__SCAN_IN ^ n8501;
  assign n12598 = ~n12597 | ~n12596;
  assign n11942 = ~n11939 | ~n13197;
  assign n11934 = ~n11933 | ~n11932;
  assign n12410 = ~n13330 | ~n12473;
  assign n12406 = ~n12405 | ~n12404;
  assign n11909 = ~n11908 | ~n11907;
  assign n11912 = ~n11911 | ~n12631;
  assign n12379 = ~n12926 | ~n11900;
  assign n12394 = ~n12393 | ~n12392;
  assign n12389 = ~REIP_REG_8__SCAN_IN | ~n12631;
  assign n12387 = ~n12386 | ~n12385;
  assign n12425 = ~n12424 | ~n12423;
  assign n13440 = ~n9731 ^ n9730;
  assign n13264 = ~n8967 ^ n8966;
  assign n9343 = ~n9342 | ~n9341;
  assign n9342 = ~n9339;
  assign n12045 = ~n12040;
  assign n12841 = ~n11589 ^ n11584;
  assign n13548 = ~n13559 | ~n13546;
  assign n10352 = ~n10351 | ~n10350;
  assign n13554 = ~n13559 | ~n13552;
  assign n13562 = ~n13559 | ~n13558;
  assign n13181 = ~n13180 | ~n13179;
  assign n13097 = ~n13096 | ~n13095;
  assign n13014 = ~n13013 | ~n13012;
  assign n12966 = ~n12965 | ~n12964;
  assign n12905 = ~n12904 | ~n12903;
  assign n12798 = ~n7008 | ~DATAI_20_;
  assign n10206 = ~n10203 & ~n10202;
  assign n10283 = ~n13566 | ~DATAI_2_;
  assign n10446 = ~n13566;
  assign n10293 = ~n13566 | ~DATAI_9_;
  assign n10273 = ~n13566 | ~DATAI_11_;
  assign n13473 = ~n13472 | ~n13471;
  assign n13457 = ~n13456 | ~n13455;
  assign n13455 = ~n13467 | ~PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n13168 = ~n13161 | ~n13472;
  assign n13353 = ~n13472 | ~n13352;
  assign n9578 = ~n9741;
  assign n13225 = ~n13472 | ~n13224;
  assign n13154 = ~PHYADDRPOINTER_REG_21__SCAN_IN ^ n8892;
  assign n13086 = PHYADDRPOINTER_REG_20__SCAN_IN ^ n8751;
  assign n12917 = ~PHYADDRPOINTER_REG_19__SCAN_IN ^ n8711;
  assign n13056 = ~n12912 ^ n12911;
  assign n12993 = ~PHYADDRPOINTER_REG_18__SCAN_IN ^ n8670;
  assign n12985 = ~n13288 | ~INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n12990 = ~n13467 | ~PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n12894 = PHYADDRPOINTER_REG_17__SCAN_IN ^ n8663;
  assign n13005 = ~n12980 ^ n12890;
  assign n12868 = n8540 ^ n8624;
  assign n9334 = n12888 & n9333;
  assign n12827 = PHYADDRPOINTER_REG_15__SCAN_IN ^ n8539;
  assign n9151 = ~n9150;
  assign n11939 = ~PHYADDRPOINTER_REG_13__SCAN_IN ^ n8435;
  assign n12741 = n8382 ^ n8381;
  assign n12465 = ~n12463 | ~n13472;
  assign n12441 = ~n13467 | ~PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n12433 = n8269 ^ n8267;
  assign n12495 = ~n13491 | ~REIP_REG_10__SCAN_IN;
  assign n11764 = ~n13467 | ~PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n12616 = ~PHYADDRPOINTER_REG_8__SCAN_IN ^ n8184;
  assign n11419 = ~n13467 | ~PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n12428 = PHYADDRPOINTER_REG_7__SCAN_IN ^ n8176;
  assign n11344 = ~n13467 | ~PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n12449 = ~PHYADDRPOINTER_REG_6__SCAN_IN ^ n8167;
  assign n12634 = PHYADDRPOINTER_REG_5__SCAN_IN ^ n8159;
  assign n12575 = PHYADDRPOINTER_REG_3__SCAN_IN ^ n8134;
  assign n10325 = ~n10324 | ~n10323;
  assign n13480 = ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n9349 = ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n12838 = ~n12836 | ~n12835;
  assign n12769 = ~n11238 ^ n11237;
  assign n12501 = ~INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n11928 = n11839 ^ n11838;
  assign n11926 = ~n11925 | ~n11924;
  assign n11436 = ~n11435 | ~n11434;
  assign n12003 = ~n12002 | ~n12001;
  assign n12001 = ~INSTQUEUE_REG_0__3__SCAN_IN | ~n12136;
  assign n12011 = ~n12010 | ~n12009;
  assign n12009 = ~INSTQUEUE_REG_0__4__SCAN_IN | ~n12136;
  assign n11989 = ~n11988 | ~n11987;
  assign n11987 = ~INSTQUEUE_REG_0__5__SCAN_IN | ~n12136;
  assign n12019 = ~n12018 | ~n12017;
  assign n12017 = ~INSTQUEUE_REG_0__7__SCAN_IN | ~n12136;
  assign n11167 = ~n11166 | ~n11165;
  assign n12550 = ~INSTQUEUE_REG_2__2__SCAN_IN | ~n12563;
  assign n12539 = ~INSTQUEUE_REG_2__5__SCAN_IN | ~n12563;
  assign n12566 = ~n12565 | ~n12564;
  assign n12564 = ~INSTQUEUE_REG_2__6__SCAN_IN | ~n12563;
  assign n11185 = ~n11184 | ~n11183;
  assign n11659 = ~INSTQUEUE_REG_4__1__SCAN_IN | ~n11701;
  assign n11677 = ~n11676 | ~n11675;
  assign n11675 = ~INSTQUEUE_REG_4__3__SCAN_IN | ~n11701;
  assign n11683 = ~INSTQUEUE_REG_4__4__SCAN_IN | ~n11701;
  assign n11667 = ~INSTQUEUE_REG_4__5__SCAN_IN | ~n11701;
  assign n11704 = ~n11703 | ~n11702;
  assign n11702 = ~INSTQUEUE_REG_4__6__SCAN_IN | ~n11701;
  assign n11693 = ~n11692 | ~n11691;
  assign n11691 = ~INSTQUEUE_REG_4__7__SCAN_IN | ~n11701;
  assign n11159 = ~n11158 | ~n11157;
  assign n12181 = ~n12180 | ~n12179;
  assign n12179 = ~INSTQUEUE_REG_6__2__SCAN_IN | ~n12276;
  assign n12165 = ~n12164 | ~n12163;
  assign n12163 = ~INSTQUEUE_REG_6__3__SCAN_IN | ~n12276;
  assign n12173 = ~n12172 | ~n12171;
  assign n12171 = ~INSTQUEUE_REG_6__4__SCAN_IN | ~n12276;
  assign n12152 = ~n12151 | ~n12150;
  assign n12150 = ~INSTQUEUE_REG_6__5__SCAN_IN | ~n12276;
  assign n12190 = ~n12189 | ~n12188;
  assign n11361 = ~n11360 | ~n11359;
  assign n11492 = ~n11491 | ~n11490;
  assign n11542 = ~n11541 | ~n11540;
  assign n11534 = ~n11533 | ~n11532;
  assign n11526 = ~n11525 | ~n11524;
  assign n11518 = ~n11517 | ~n11516;
  assign n11510 = ~n11509 | ~n11508;
  assign n10693 = ~n10692 | ~n10691;
  assign n11007 = ~n11006 | ~n11005;
  assign n10999 = ~n10998 | ~n10997;
  assign n11795 = ~n11794 | ~n11793;
  assign n11771 = ~n11770 | ~n11769;
  assign n11769 = ~INSTQUEUE_REG_12__3__SCAN_IN | ~n11882;
  assign n11779 = ~n11778 | ~n11777;
  assign n11741 = ~n11740 | ~n11739;
  assign n11739 = ~INSTQUEUE_REG_12__5__SCAN_IN | ~n11882;
  assign n11803 = ~n11802 | ~n11801;
  assign n11874 = n10621 | n10886;
  assign n11787 = ~n11786 | ~n11785;
  assign n12061 = ~n12060 | ~n12059;
  assign n12059 = ~INSTQUEUE_REG_14__1__SCAN_IN | ~n12248;
  assign n12074 = ~n12073 | ~n12072;
  assign n12072 = ~INSTQUEUE_REG_14__5__SCAN_IN | ~n12248;
  assign n12090 = ~n12089 | ~n12088;
  assign n12082 = ~n12081 | ~n12080;
  assign n12650 = ~REIP_REG_5__SCAN_IN;
  assign n12418 = ~REIP_REG_7__SCAN_IN;
  assign n9956 = ~REIP_REG_23__SCAN_IN;
  assign n12632 = ~n12631 | ~n12630;
  assign n12462 = ~n12446 | ~n12651;
  assign n12652 = ~n12651 | ~n12650;
  assign n11657 = ~REIP_REG_4__SCAN_IN | ~n12593;
  assign n11652 = ~n11651 | ~n11650;
  assign n12594 = ~REIP_REG_3__SCAN_IN | ~n12593;
  assign n12299 = ~n12298 | ~n12297;
  assign n12296 = ~n12283 | ~n12282;
  assign n11729 = ~n11727 & ~n11726;
  assign n11960 = ~n11947 | ~PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n12702 = n12698 & n12697;
  assign n13522 = ~EBX_REG_18__SCAN_IN | ~n13560;
  assign n11090 = ~n13185 | ~n12473;
  assign n10868 = ~n13185 | ~n12391;
  assign n13537 = ~n13536 | ~n13535;
  assign n13543 = ~n13542 | ~n13541;
  assign n10471 = ~n13185 | ~n12297;
  assign n10935 = ~n13559 | ~n11954;
  assign n13394 = ~n7008 | ~DATAI_31_;
  assign n9309 = ~n9308 | ~n9307;
  assign n9257 = ~n9256 | ~n9255;
  assign n9086 = ~n9085 | ~n9084;
  assign n8939 = ~n8938 | ~n8937;
  assign n8799 = ~n8798 | ~n8797;
  assign n12659 = ~n12658 | ~n12657;
  assign n12532 = ~n12531 | ~n12530;
  assign n12486 = ~n12485 | ~n12484;
  assign n11025 = ~n13176 | ~n12473;
  assign n10822 = ~n13176 | ~n12391;
  assign n10360 = ~n13176 | ~n12297;
  assign n10172 = ~n10206 | ~DATAO_REG_30__SCAN_IN;
  assign n10163 = ~n10206 | ~DATAO_REG_29__SCAN_IN;
  assign n10127 = ~n10206 | ~DATAO_REG_28__SCAN_IN;
  assign n10119 = ~n10206 | ~DATAO_REG_27__SCAN_IN;
  assign n10107 = ~n10206 | ~DATAO_REG_26__SCAN_IN;
  assign n10103 = ~n10206 | ~DATAO_REG_25__SCAN_IN;
  assign n10099 = ~n10206 | ~DATAO_REG_24__SCAN_IN;
  assign n10095 = ~n10206 | ~DATAO_REG_23__SCAN_IN;
  assign n10091 = ~n10206 | ~DATAO_REG_22__SCAN_IN;
  assign n10087 = ~n10206 | ~DATAO_REG_21__SCAN_IN;
  assign n10123 = ~n10206 | ~DATAO_REG_20__SCAN_IN;
  assign n10083 = ~n10206 | ~DATAO_REG_19__SCAN_IN;
  assign n10115 = ~n10206 | ~DATAO_REG_18__SCAN_IN;
  assign n10111 = ~n10206 | ~DATAO_REG_17__SCAN_IN;
  assign n10167 = ~n10206 | ~DATAO_REG_16__SCAN_IN;
  assign n10143 = ~n10206 | ~DATAO_REG_15__SCAN_IN;
  assign n10200 = ~n10206 | ~DATAO_REG_14__SCAN_IN;
  assign n10155 = ~n10206 | ~DATAO_REG_13__SCAN_IN;
  assign n10151 = ~n10206 | ~DATAO_REG_12__SCAN_IN;
  assign n10180 = ~n10206 | ~DATAO_REG_11__SCAN_IN;
  assign n10184 = ~n10206 | ~DATAO_REG_10__SCAN_IN;
  assign n10135 = ~n10206 | ~DATAO_REG_9__SCAN_IN;
  assign n10192 = ~n10206 | ~DATAO_REG_8__SCAN_IN;
  assign n10131 = ~n10206 | ~DATAO_REG_7__SCAN_IN;
  assign n10147 = ~n10206 | ~DATAO_REG_6__SCAN_IN;
  assign n10139 = ~n10206 | ~DATAO_REG_5__SCAN_IN;
  assign n10207 = ~n10206 | ~DATAO_REG_4__SCAN_IN;
  assign n10176 = ~n10206 | ~DATAO_REG_3__SCAN_IN;
  assign n10196 = ~n10206 | ~DATAO_REG_2__SCAN_IN;
  assign n10188 = ~n10206 | ~DATAO_REG_1__SCAN_IN;
  assign n10159 = ~n10206 | ~DATAO_REG_0__SCAN_IN;
  assign n13570 = ~n13569 | ~n13568;
  assign n13155 = n13472 & n13154;
  assign n13087 = n13472 & n13086;
  assign n8429 = ~n12762 | ~n7672;
  assign n7672 = ~n13472 | ~n11939;
  assign n11843 = ~n12391 | ~n13463;
  assign n11842 = ~n11837 | ~n11836;
  assign n10569 = ~n10564 | ~n10563;
  assign n10481 = ~n10480 | ~n10479;
  assign n13360 = ~n13359 | ~INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n13503 = ~n13500 | ~INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n13499 = ~n13479 | ~INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n13379 = ~n13415 | ~INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n13260 = ~n13255 | ~n13254;
  assign n13055 = ~n13249 & ~n13053;
  assign n13003 = ~n13114 | ~n13002;
  assign n12759 = ~n12837 | ~INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n12784 = ~INSTADDRPOINTER_REG_12__SCAN_IN | ~n12783;
  assign n12525 = ~INSTADDRPOINTER_REG_11__SCAN_IN | ~n12783;
  assign n12518 = ~n12511 | ~n12510;
  assign n12505 = ~n12504 | ~n12503;
  assign n11898 = ~n11897 | ~n11896;
  assign n11897 = ~n11893 | ~n11892;
  assign n11562 = ~INSTADDRPOINTER_REG_7__SCAN_IN | ~n11917;
  assign n12214 = ~n12198 | ~n12197;
  assign n11411 = ~INSTADDRPOINTER_REG_5__SCAN_IN | ~n12201;
  assign n11405 = ~n11404 | ~n11403;
  assign n11582 = ~n11581 | ~n11580;
  assign n11104 = ~n11092 | ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n11103 = ~n11102 & ~n11101;
  assign n11092 = ~n11326 | ~n11395;
  assign n11396 = ~n11394 & ~n11393;
  assign n11835 = ~n11859 | ~n11833;
  assign n11833 = ~n11832 | ~n11831;
  assign n11818 = ~n11859 | ~n11816;
  assign n11827 = ~n11859 | ~n11825;
  assign n11863 = ~n11860 | ~n11859;
  assign n12116 = ~INSTQUEUE_REG_0__0__SCAN_IN | ~n12136;
  assign n12108 = ~INSTQUEUE_REG_0__1__SCAN_IN | ~n12136;
  assign n12124 = ~INSTQUEUE_REG_0__2__SCAN_IN | ~n12136;
  assign n12137 = ~INSTQUEUE_REG_0__6__SCAN_IN | ~n12136;
  assign n12331 = ~INSTQUEUE_REG_2__0__SCAN_IN | ~n12563;
  assign n12343 = ~INSTQUEUE_REG_2__1__SCAN_IN | ~n12563;
  assign n12355 = ~INSTQUEUE_REG_2__3__SCAN_IN | ~n12563;
  assign n12366 = ~INSTQUEUE_REG_2__4__SCAN_IN | ~n12563;
  assign n12377 = ~INSTQUEUE_REG_2__7__SCAN_IN | ~n12563;
  assign n11464 = ~INSTQUEUE_REG_4__0__SCAN_IN | ~n11701;
  assign n11472 = ~INSTQUEUE_REG_4__2__SCAN_IN | ~n11701;
  assign n12257 = ~INSTQUEUE_REG_6__0__SCAN_IN | ~n12276;
  assign n12265 = ~INSTQUEUE_REG_6__1__SCAN_IN | ~n12276;
  assign n12277 = ~INSTQUEUE_REG_6__7__SCAN_IN | ~n12276;
  assign n11870 = ~INSTQUEUE_REG_12__0__SCAN_IN | ~n11882;
  assign n11883 = ~INSTQUEUE_REG_12__1__SCAN_IN | ~n11882;
  assign n12221 = ~INSTQUEUE_REG_14__0__SCAN_IN | ~n12248;
  assign n12249 = ~INSTQUEUE_REG_14__2__SCAN_IN | ~n12248;
  assign n12229 = ~INSTQUEUE_REG_14__3__SCAN_IN | ~n12248;
  assign n12237 = ~INSTQUEUE_REG_14__4__SCAN_IN | ~n12248;
  assign n7004 = ~n11156 & ~n11155;
  assign n7005 = ~n13567 & ~n10515;
  assign n11852 = n8018 ^ n10635;
  assign n8018 = ~n7949 | ~n7948;
  assign n7008 = ~n13178 & ~n8796;
  assign n10027 = ~n10025;
  assign n13481 = ~INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n7009 = n8265 | n8264;
  assign n12415 = ~PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n7010 = ~n9102 & ~n11155;
  assign n7011 = ~n13389 & ~n11155;
  assign n7597 = ~FLUSH_REG_SCAN_IN;
  assign n9883 = ~REIP_REG_31__SCAN_IN;
  assign n9102 = ~n7261 & ~n7260;
  assign n8970 = ~PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n8148 = ~EAX_REG_4__SCAN_IN;
  assign n8533 = ~EAX_REG_15__SCAN_IN;
  assign n8268 = ~EAX_REG_10__SCAN_IN;
  assign n8377 = ~EAX_REG_12__SCAN_IN;
  assign n8971 = ~PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n7012 = n11481 | n12307;
  assign n9169 = ~REIP_REG_21__SCAN_IN;
  assign n12638 = ~PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n8001 = ~INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n8067 = ~n8090;
  assign n8177 = ~EAX_REG_7__SCAN_IN;
  assign n8185 = ~EAX_REG_8__SCAN_IN;
  assign n7013 = n8535 | n8534;
  assign n7014 = n8470 | n8469;
  assign n7015 = n8379 | n8378;
  assign n7016 = n8193 | n8418;
  assign n9657 = ~n9057;
  assign n13491 = ~n10034 & ~STATE2_REG_0__SCAN_IN;
  assign n13222 = ~n13491;
  assign n7017 = n10211 | n8125;
  assign n7292 = ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n7373 = ~n7388;
  assign n7855 = ~n8004;
  assign n7329 = ~n7328;
  assign n7045 = ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n7183 = ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n8119 = ~EAX_REG_0__SCAN_IN;
  assign n8783 = ~EAX_REG_21__SCAN_IN;
  assign n8467 = ~EAX_REG_14__SCAN_IN;
  assign n7148 = ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n8924 = ~EAX_REG_22__SCAN_IN;
  assign n8186 = ~PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n7487 = ~n7484 & ~n7483;
  assign n7546 = ~n7545;
  assign n7959 = ~n7928 & ~n7335;
  assign n9572 = ~n13144;
  assign n10780 = ~n10779;
  assign n7398 = ~n7408;
  assign n9726 = ~n13103;
  assign n13163 = ~PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n9080 = ~n8999 & ~n8998;
  assign n12309 = ~n12322;
  assign n11483 = ~n11495;
  assign n10534 = ~n10533;
  assign n7601 = ~n9092 | ~n10245;
  assign n8796 = ~n8101 | ~n8791;
  assign n12477 = ~n12026 | ~n12025;
  assign n10076 = ~n10515 & ~n9092;
  assign n12961 = ~n12900 & ~n12899;
  assign n9301 = ~n9303;
  assign n8540 = ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n7669 = ~n10209;
  assign n11593 = ~n11589;
  assign n10787 = ~n11847;
  assign n7657 = ~n8943;
  assign n12963 = ~n9543;
  assign n12790 = ~EAX_REG_19__SCAN_IN;
  assign n10441 = ~EAX_REG_30__SCAN_IN;
  assign n10432 = ~EAX_REG_5__SCAN_IN;
  assign n10826 = ~n10825 | ~n10824;
  assign n11578 = ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n9918 = ~REIP_REG_18__SCAN_IN;
  assign n12676 = ~REIP_REG_16__SCAN_IN;
  assign n9648 = ~n7299;
  assign n9501 = ~n8195;
  assign n7018 = ~n9501 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n9053 = ~n7032 | ~n7521;
  assign n9636 = ~n9053;
  assign n9051 = ~n7526 | ~n10374;
  assign n7267 = ~n7043 | ~n7048;
  assign n9640 = ~n7032 | ~n7631;
  assign n9522 = ~n9640;
  assign n8587 = ~n7043 | ~n7631;
  assign n7026 = ~n9657 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n9642 = ~n7631 | ~n7637;
  assign n8591 = ~n7048 | ~n10374;
  assign n7056 = ~n7055 & ~n7054;
  assign n9665 = ~n7288;
  assign n9602 = ~n8196;
  assign n9599 = ~n7286;
  assign n9656 = ~n8585;
  assign n7087 = ~n7071 | ~n7070;
  assign n9662 = ~n8551;
  assign n9607 = ~n9642;
  assign n9610 = ~n9051;
  assign n7086 = ~n7085 | ~n7084;
  assign n7614 = ~n10499 & ~n11156;
  assign n7094 = ~n9665 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n7097 = ~n9602 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n7096 = ~n9610 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n7105 = ~n9599 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n7116 = ~n7115 | ~n7114;
  assign n13389 = ~n7117 & ~n7116;
  assign n7465 = ~n7614 & ~n13389;
  assign n8498 = ~n10499 | ~n11156;
  assign n7159 = ~n7137 & ~n7136;
  assign n7158 = ~n7157 & ~n7156;
  assign n7191 = ~n8551 & ~n9058;
  assign n9092 = ~n10574;
  assign n7229 = ~n7213 | ~n7212;
  assign n7228 = ~n7227 | ~n7226;
  assign n7441 = ~n7413 & ~n7231;
  assign n7394 = ~n9132 & ~n8792;
  assign n7411 = ~n7518 & ~n7508;
  assign n8574 = ~n7513 | ~n7411;
  assign n8791 = ~n13389;
  assign n7326 = ~n10341 & ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n7349 = ~n7325 & ~n7324;
  assign n7328 = ~n7327 & ~n7326;
  assign n7334 = ~INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~n7332;
  assign n7382 = ~n7334 & ~n7333;
  assign n7383 = INSTQUEUERD_ADDR_REG_4__SCAN_IN | n7382;
  assign n7401 = ~n7383 & ~n11628;
  assign n8082 = ~n10499 | ~n10515;
  assign n7340 = ~n7339 | ~n7338;
  assign n7365 = n7352 | n7351;
  assign n7353 = n7400 | n10490;
  assign n7363 = n7365 | n7364;
  assign n7375 = n7371 | n7370;
  assign n7380 = ~n7379 & ~n7378;
  assign n7387 = ~n7381 & ~n7380;
  assign n7390 = ~n7389 & ~n7388;
  assign n7397 = ~n7396 & ~n7395;
  assign n8946 = ~n7398 | ~n9092;
  assign n10075 = ~n9100 | ~n7399;
  assign n8948 = ~n7407 & ~n7406;
  assign n7516 = ~n10391;
  assign n9107 = ~n7650 & ~n7412;
  assign n8804 = ~n9107 | ~n7464;
  assign n7414 = ~n7436 & ~n7613;
  assign n7415 = ~n7425 & ~n10574;
  assign n9099 = n7419 | n7418;
  assign n7420 = n11637 & n9102;
  assign n7424 = n7423 | n7422;
  assign n7592 = ~n8496 & ~n7424;
  assign n7426 = ~n7425 & ~n10748;
  assign n7434 = ~n7426 & ~n13389;
  assign n7506 = ~n7434 | ~n7433;
  assign n7447 = ~n7458 | ~n7435;
  assign n9111 = ~n8796 & ~n9723;
  assign n7440 = ~n9111 & ~n7436;
  assign n7437 = ~n10240 & ~n7231;
  assign n7453 = ~n7447 | ~n7446;
  assign n7457 = ~n7495 | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n9787 = ~n11497 & ~STATE2_REG_1__SCAN_IN;
  assign n7568 = ~n7457 | ~n7456;
  assign n7567 = ~n7475 | ~n7474;
  assign n7559 = ~n7568 | ~n7567;
  assign n7479 = ~n7495 | ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7558 = ~n7485 | ~n7487;
  assign n7490 = ~n7486 | ~n7558;
  assign n7494 = ~n7495 | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n11440 = n11357 | n7499;
  assign n11854 = ~n12588;
  assign n7512 = n7506 & n11647;
  assign n7510 = ~n7507 | ~n10045;
  assign n7509 = ~n8796 | ~n7508;
  assign n7511 = ~n7510 | ~n7509;
  assign n7514 = ~n7512 & ~n7511;
  assign n7515 = ~n9111 & ~n8792;
  assign n7517 = ~n7516 | ~n7515;
  assign n7519 = ~n8801 | ~n8008;
  assign n7520 = ~n9117;
  assign n7544 = ~n9139 | ~n7520;
  assign n7523 = ~n10374 & ~n7521;
  assign n7522 = ~n10341 & ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n7524 = ~n7523 & ~n7522;
  assign n7525 = ~n7524 & ~n7631;
  assign n7534 = ~n7544 | ~n7525;
  assign n7545 = ~n8814 & ~n8574;
  assign n7527 = ~n10374 & ~n8135;
  assign n7528 = ~n7527 & ~n7526;
  assign n10363 = ~n7528 | ~n8591;
  assign n7532 = n7545 & n10363;
  assign n7529 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7530 = n7529 ^ INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n7531 = ~n7530 & ~n7570;
  assign n7533 = ~n7532 & ~n7531;
  assign n7535 = ~n7534 | ~n7533;
  assign n10362 = n7536 | n7535;
  assign n7587 = n12145 | n7627;
  assign n7554 = ~n10616 & ~n7561;
  assign n7547 = n10341 ^ INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n7552 = ~n7544 | ~n7547;
  assign n7550 = ~n7547 & ~n7546;
  assign n7548 = ~INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7549 = ~n7570 & ~n7548;
  assign n7551 = ~n7550 & ~n7549;
  assign n7553 = ~n7552 | ~n7551;
  assign n10338 = n7554 | n7553;
  assign n7581 = ~n10637 & ~n7628;
  assign n7569 = ~n7561;
  assign n7566 = ~n7936 | ~n7569;
  assign n10373 = ~n7637;
  assign n7562 = ~n10373 | ~n10341;
  assign n7564 = ~n8574 & ~n7562;
  assign n7563 = ~n7570 & ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n7565 = ~n7564 & ~n7563;
  assign n10369 = ~n7566 | ~n7565;
  assign n7575 = ~n7577 & ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n11949 = n7568 ^ n7567;
  assign n7574 = ~n11949 | ~n7569;
  assign n7572 = ~n8574 | ~n8118;
  assign n7571 = ~n7570 | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n7573 = ~n7572 | ~n7571;
  assign n10383 = ~n7574 | ~n7573;
  assign n7576 = ~n7575 & ~n10383;
  assign n7578 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n7577;
  assign n7596 = ~INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n7598 = ~n7596 & ~n11813;
  assign n7599 = ~n7598 | ~n7597;
  assign n7609 = ~FLUSH_REG_SCAN_IN & ~MORE_REG_SCAN_IN;
  assign n7604 = ~n7602 & ~n8946;
  assign n7603 = ~n8949 & ~n9092;
  assign n7607 = ~n7604 & ~n7603;
  assign n7605 = ~n10937 | ~n7641;
  assign n10055 = ~n7605 & ~n11647;
  assign n7606 = ~n10055 & ~READY_N;
  assign n7608 = ~n7607 & ~n7606;
  assign n7610 = ~n7609 & ~n10043;
  assign n7617 = ~n7623 | ~n9139;
  assign n7619 = ~n7617 | ~n10033;
  assign n7618 = ~n9117 | ~n7650;
  assign n7621 = ~n7619 | ~n7618;
  assign n7620 = ~n8948 & ~n8946;
  assign n7622 = ~n7621 & ~n7620;
  assign n10071 = ~n7622 & ~n13389;
  assign n7625 = ~n10071 & ~n7664;
  assign n7630 = ~n11813 & ~FLUSH_REG_SCAN_IN;
  assign n7632 = ~n7631 | ~n7630;
  assign n8978 = ~n8980 & ~n7641;
  assign n7647 = ~n9156 | ~n8978;
  assign n7642 = ~STATE2_REG_1__SCAN_IN & ~n10490;
  assign n10063 = ~n11813 & ~STATE2_REG_0__SCAN_IN;
  assign n7644 = ~n10063 | ~READY_N;
  assign n10056 = ~n10490 | ~STATE2_REG_2__SCAN_IN;
  assign n7651 = ~n10490 | ~n10488;
  assign n7652 = ~n10056 | ~n7651;
  assign n7653 = ~n7652 & ~n10063;
  assign n7655 = ~STATE2_REG_0__SCAN_IN | ~STATE2_REG_3__SCAN_IN;
  assign n7656 = ~STATE2_REG_2__SCAN_IN & ~n12680;
  assign n12684 = ~n7656 | ~STATE2_REG_0__SCAN_IN;
  assign n7658 = ~n7657 | ~n12684;
  assign U3148 = n7663 | n7662;
  assign n12305 = ~STATE2_REG_3__SCAN_IN & ~STATE2_REG_2__SCAN_IN;
  assign n10060 = ~n7665 | ~n11480;
  assign n7666 = ~n10060 | ~n10490;
  assign n7668 = ~n10056;
  assign n7667 = ~n11813 & ~STATEBS16_REG_SCAN_IN;
  assign n10209 = ~n7668 & ~n7667;
  assign n7730 = n7729 | n7728;
  assign n7943 = n7793 | n7792;
  assign n7854 = ~n8003;
  assign n7920 = ~n11949 | ~n10490;
  assign n8079 = ~n7918 & ~n7917;
  assign n7927 = ~n7920 | ~n7992;
  assign n8090 = ~n7928 | ~n7929;
  assign n7942 = ~n7935 | ~n7986;
  assign n7975 = ~n7942 | ~n7987;
  assign n7974 = ~n7947 & ~n7946;
  assign n7965 = ~n7964 & ~n8046;
  assign n8063 = ~n7968 | ~n7967;
  assign n11820 = n7975 ^ n7974;
  assign n7982 = ~n11820 | ~n8092;
  assign n7978 = ~n8019;
  assign n7977 = ~n7976 & ~n8002;
  assign n7979 = ~n7978 & ~n7977;
  assign n7980 = ~n7979 & ~n10240;
  assign n7981 = ~n7980 & ~n7996;
  assign n8016 = ~n7983 | ~INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n7985 = ~n8016;
  assign n10327 = ~n7985 & ~n7984;
  assign n7989 = ~n7987 | ~n7986;
  assign n10886 = ~n7995 | ~n7994;
  assign n8000 = ~n10886 & ~n8082;
  assign n7998 = ~n7996;
  assign n7997 = ~n10076 | ~n8004;
  assign n7999 = ~n7998 | ~n7997;
  assign n10216 = ~n8000 & ~n7999;
  assign n10224 = ~n10216 & ~n8001;
  assign n8007 = ~n8002;
  assign n8005 = ~n8004 | ~n8003;
  assign n8006 = ~n10076 | ~n8005;
  assign n8010 = ~n8007 & ~n8006;
  assign n8009 = ~n8008 | ~n10499;
  assign n10222 = ~n8010 & ~n8009;
  assign n8012 = ~n8011 | ~n10222;
  assign n8015 = ~n8013 & ~n8012;
  assign n10328 = ~n8015 & ~n8014;
  assign n10474 = ~n8017 | ~n8016;
  assign n11845 = ~n11852;
  assign n8024 = ~n11845 | ~n8092;
  assign n8021 = ~n8020 & ~n8019;
  assign n8022 = ~n8021 & ~n10240;
  assign n8023 = ~n8022 | ~n8032;
  assign n8025 = ~n8024 | ~n8023;
  assign n11332 = ~INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n8028 = ~n8026 & ~n11332;
  assign n10473 = ~n8027 & ~n8028;
  assign n10476 = ~n10474 | ~n10473;
  assign n10565 = ~n10476 | ~n8029;
  assign n8033 = ~n8032 ^ n8031;
  assign n10566 = ~n8038 & ~n8037;
  assign n11027 = ~n8040 | ~n8039;
  assign n8050 = ~n8043 & ~n10240;
  assign n12196 = ~INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n8054 = ~n8051 & ~n12196;
  assign n11029 = ~n11027 | ~n11028;
  assign n11338 = ~n11029 | ~n8055;
  assign n11340 = ~n11339 | ~n11338;
  assign n11413 = ~n11340 | ~n8057;
  assign n11415 = ~n11413 | ~n11414;
  assign n11759 = ~n11415 | ~n8078;
  assign n11761 = ~n11759 | ~n11758;
  assign n8096 = ~n11838 | ~n11839;
  assign n8097 = ~n12438 | ~n12436;
  assign n8098 = ~n12469;
  assign n8099 = ~n8098 | ~n12467;
  assign n12746 = ~n8099 | ~n12466;
  assign n8100 = ~n12746 | ~n12744;
  assign n8478 = ~n8100 | ~n12743;
  assign n9633 = ~n8101 & ~n11497;
  assign n9708 = ~n11478 & ~STATE2_REG_2__SCAN_IN;
  assign n8103 = ~EAX_REG_2__SCAN_IN;
  assign n12292 = PHYADDRPOINTER_REG_1__SCAN_IN ^ PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n8104 = ~n12292;
  assign n8106 = ~n9698 | ~n8104;
  assign n8105 = ~n9708 | ~PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n8115 = ~n8136 & ~n8111;
  assign n8112 = ~n11497 | ~PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n10213 = ~n10886 | ~n11156;
  assign n8124 = ~PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n8125 = ~n8124 & ~STATE2_REG_2__SCAN_IN;
  assign n10313 = ~n10305 & ~n10304;
  assign n8149 = ~PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n8150 = ~n9535 & ~n8149;
  assign n10461 = ~n10351 & ~n10350;
  assign n10666 = ~n10461 | ~n10460;
  assign n8198 = ~n8195 & ~n8194;
  assign n8197 = ~n8196 & ~n9056;
  assign n8203 = ~n8198 & ~n8197;
  assign n8201 = ~n9640 & ~n9058;
  assign n8200 = ~n9053 & ~n8199;
  assign n8202 = ~n8201 & ~n8200;
  assign n8205 = ~n9599 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n8204 = ~n9662 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n8209 = ~n9672 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n8208 = ~n9673 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n8213 = ~n8209 | ~n8208;
  assign n8211 = ~n9648 | ~INSTQUEUE_REG_6__0__SCAN_IN;
  assign n8210 = ~n9653 | ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n8212 = ~n8211 | ~n8210;
  assign n8221 = ~n8213 & ~n8212;
  assign n8215 = ~n9656 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n8214 = ~n9665 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n8219 = ~n8215 | ~n8214;
  assign n8217 = ~n9647 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n8216 = ~n9610 | ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n8218 = ~n8217 | ~n8216;
  assign n8220 = ~n8219 & ~n8218;
  assign n8223 = ~n9657 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n8222 = ~n9607 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n8231 = ~n9656 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n8230 = ~n9610 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n8233 = ~n9672 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n8232 = ~n7003 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n8234 = ~n8233 | ~n8232;
  assign n8237 = ~n9665 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n8236 = ~n9636 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n8239 = ~n9599 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n8238 = ~n9602 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n8245 = ~n9522 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n8244 = ~n9607 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n8247 = ~n9501 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n8246 = ~n9648 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n8251 = ~n9673 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n8250 = ~n9653 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n8253 = ~n9647 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n8252 = ~n9662 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n8276 = ~n9599 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n8275 = ~n9665 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n8280 = ~n8276 | ~n8275;
  assign n8278 = ~n9607 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n8277 = ~n9653 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n8279 = ~n8278 | ~n8277;
  assign n8288 = ~n8280 & ~n8279;
  assign n8282 = ~n9656 | ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n8281 = ~n9522 | ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n8286 = ~n8282 | ~n8281;
  assign n8284 = ~n9647 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n8283 = ~n9673 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n8285 = ~n8284 | ~n8283;
  assign n8287 = ~n8286 & ~n8285;
  assign n8290 = ~n9501 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n8289 = ~n9602 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n8294 = ~n8290 | ~n8289;
  assign n8292 = ~n9610 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n8291 = ~n9662 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n8293 = ~n8292 | ~n8291;
  assign n8302 = ~n8294 & ~n8293;
  assign n8296 = ~n9657 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n8295 = ~n9636 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n8298 = ~n9672 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n8297 = ~n9648 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n8299 = ~n8298 | ~n8297;
  assign n8301 = ~n8300 & ~n8299;
  assign n8305 = n8304 | n8303;
  assign n8311 = ~n9672 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n8310 = ~n9607 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n8315 = ~n8311 | ~n8310;
  assign n8313 = ~n9501 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n8312 = ~n9665 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n8314 = ~n8313 | ~n8312;
  assign n8323 = ~n8315 & ~n8314;
  assign n8317 = ~n9656 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n8316 = ~n9673 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n8321 = ~n8317 | ~n8316;
  assign n8319 = ~n9647 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n8318 = ~n9522 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n8320 = ~n8319 | ~n8318;
  assign n8322 = ~n8321 & ~n8320;
  assign n8325 = ~n9610 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n8324 = ~n9653 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n8329 = ~n8325 | ~n8324;
  assign n8327 = ~n9636 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n8326 = ~n9648 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n8328 = ~n8327 | ~n8326;
  assign n8337 = ~n8329 & ~n8328;
  assign n8331 = ~n7003 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n8330 = ~n9602 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n8335 = ~n8331 | ~n8330;
  assign n8333 = ~n9599 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n8332 = ~n9662 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n8334 = ~n8333 | ~n8332;
  assign n8336 = ~n8335 & ~n8334;
  assign n8340 = n8339 | n8338;
  assign n8347 = ~n9647 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n8346 = ~n9662 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n8351 = ~n8347 | ~n8346;
  assign n8349 = ~n9602 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n8348 = ~n9607 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n8350 = ~n8349 | ~n8348;
  assign n8359 = ~n8351 & ~n8350;
  assign n8353 = ~n9672 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n8352 = ~n9665 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n8357 = ~n8353 | ~n8352;
  assign n8355 = ~n9673 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n8354 = ~n9648 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n8356 = ~n8355 | ~n8354;
  assign n8358 = ~n8357 & ~n8356;
  assign n8361 = ~n9656 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n8360 = ~n9522 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n8365 = ~n8361 | ~n8360;
  assign n8363 = ~n9657 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n8362 = ~n9653 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n8364 = ~n8363 | ~n8362;
  assign n8373 = ~n8365 & ~n8364;
  assign n8367 = ~n9501 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n8366 = ~n9599 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n8371 = ~n8367 | ~n8366;
  assign n8369 = ~n9610 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n8368 = ~n9636 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n8370 = ~n8369 | ~n8368;
  assign n8372 = ~n8371 & ~n8370;
  assign n8386 = ~n9656 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n8385 = ~n9636 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n8390 = ~n8386 | ~n8385;
  assign n8388 = ~n9672 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n8387 = ~n9610 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n8389 = ~n8388 | ~n8387;
  assign n8398 = ~n8390 & ~n8389;
  assign n8392 = ~n9665 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n8391 = ~n9607 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n8396 = ~n8392 | ~n8391;
  assign n8394 = ~n9599 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n8393 = ~n9653 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n8395 = ~n8394 | ~n8393;
  assign n8397 = ~n8396 & ~n8395;
  assign n8400 = ~n9501 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n8399 = ~n9602 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n8404 = ~n8400 | ~n8399;
  assign n8402 = ~n7003 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n8401 = ~n9648 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n8412 = ~n8404 & ~n8403;
  assign n8406 = ~n9647 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n8405 = ~n9522 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n8410 = ~n8406 | ~n8405;
  assign n8408 = ~n9673 | ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n8407 = ~n9662 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n8409 = ~n8408 | ~n8407;
  assign n8411 = ~n8410 & ~n8409;
  assign n8415 = ~n8418;
  assign n8420 = ~n9535 & ~n8434;
  assign U2973 = n8429 | n8428;
  assign n8468 = ~PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n8475 = ~n13164 & ~n8468;
  assign n8473 = n12613 | n9789;
  assign n8437 = ~n9672 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n8436 = ~n9522 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n8441 = ~n8437 | ~n8436;
  assign n8439 = ~n9647 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n8438 = ~n9648 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n8440 = ~n8439 | ~n8438;
  assign n8449 = ~n8441 & ~n8440;
  assign n8443 = ~n9501 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n8442 = ~n9657 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n8447 = ~n8443 | ~n8442;
  assign n8445 = ~n9610 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n8444 = ~n9607 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n8446 = ~n8445 | ~n8444;
  assign n8448 = ~n8447 & ~n8446;
  assign n8451 = ~n9656 | ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n8450 = ~n9673 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n8455 = ~n8451 | ~n8450;
  assign n8453 = ~n9602 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n8452 = ~n9636 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n8454 = ~n8453 | ~n8452;
  assign n8463 = ~n8455 & ~n8454;
  assign n8457 = ~n9599 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n8456 = ~n9665 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n8461 = ~n8457 | ~n8456;
  assign n8459 = ~n9653 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n8458 = ~n9662 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n8460 = ~n8459 | ~n8458;
  assign n8462 = ~n8461 & ~n8460;
  assign n8464 = ~n8463 | ~n8462;
  assign n8466 = ~n8465 & ~n8464;
  assign n8469 = ~n9535 & ~n8468;
  assign n8480 = ~n8478 | ~n8477;
  assign n8481 = ~INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n8483 = n12844 | n13465;
  assign U2972 = n8486 | n8485;
  assign n8494 = ~n10391 | ~n8487;
  assign n8497 = n8496 | n8495;
  assign n8503 = ~n9672 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n8502 = ~n7003 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n8507 = ~n8503 | ~n8502;
  assign n8505 = ~n9656 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n8504 = ~n9673 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n8506 = ~n8505 | ~n8504;
  assign n8515 = ~n8507 & ~n8506;
  assign n8509 = ~n9501 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n8508 = ~n9648 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n8513 = ~n8509 | ~n8508;
  assign n8511 = ~n9607 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n8510 = ~n9653 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n8512 = ~n8511 | ~n8510;
  assign n8514 = ~n8513 & ~n8512;
  assign n8531 = ~n8515 | ~n8514;
  assign n8517 = ~n9647 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n8516 = ~n9602 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n8521 = ~n8517 | ~n8516;
  assign n8519 = ~n9522 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n8518 = ~n9610 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n8520 = ~n8519 | ~n8518;
  assign n8529 = ~n8521 & ~n8520;
  assign n8523 = ~n9665 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n8522 = ~n9636 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n8527 = ~n8523 | ~n8522;
  assign n8525 = ~n9599 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n8524 = ~n9662 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n8526 = ~n8525 | ~n8524;
  assign n8528 = ~n8527 & ~n8526;
  assign n8530 = ~n8529 | ~n8528;
  assign n8532 = ~n8531 & ~n8530;
  assign n8534 = ~n9535 & ~n12821;
  assign n8543 = ~n9656 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n8542 = ~n9607 | ~INSTQUEUE_REG_15__0__SCAN_IN;
  assign n8547 = ~n8543 | ~n8542;
  assign n8545 = ~n9610 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n8544 = ~n9602 | ~INSTQUEUE_REG_4__0__SCAN_IN;
  assign n8546 = ~n8545 | ~n8544;
  assign n8573 = ~n8547 & ~n8546;
  assign n8550 = ~n8587 & ~n9058;
  assign n8549 = ~n9053 & ~n8548;
  assign n8555 = ~n8550 & ~n8549;
  assign n8553 = ~n8593 & ~n9052;
  assign n8552 = ~n8551 & ~n9056;
  assign n8554 = ~n8553 & ~n8552;
  assign n8571 = ~n8555 | ~n8554;
  assign n8557 = ~n9501 | ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n8556 = ~n9673 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n8561 = ~n8557 | ~n8556;
  assign n8559 = ~n9522 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n8558 = ~n9665 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n8560 = ~n8559 | ~n8558;
  assign n8569 = ~n8561 & ~n8560;
  assign n8563 = ~n9599 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n8562 = ~n9648 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n8567 = ~n8563 | ~n8562;
  assign n8565 = ~n9672 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n8564 = ~n9657 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n8566 = ~n8565 | ~n8564;
  assign n8568 = ~n8567 & ~n8566;
  assign n8570 = ~n8569 | ~n8568;
  assign n8572 = ~n8571 & ~n8570;
  assign n9696 = ~n8574 & ~n10490;
  assign n8576 = ~EAX_REG_16__SCAN_IN;
  assign n8577 = ~n11497 | ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n8589 = ~n8585 & ~n8584;
  assign n8588 = ~n8587 & ~n8586;
  assign n8597 = ~n8589 & ~n8588;
  assign n8595 = ~n8591 & ~n8590;
  assign n8594 = ~n8593 & ~n8592;
  assign n8596 = ~n8595 & ~n8594;
  assign n8601 = ~n8597 | ~n8596;
  assign n8599 = ~n9599 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n8598 = ~n9602 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n8600 = ~n8599 | ~n8598;
  assign n8621 = ~n8601 & ~n8600;
  assign n8603 = ~n9501 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n8602 = ~n9662 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n8607 = ~n8603 | ~n8602;
  assign n8605 = ~n9610 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n8604 = ~n9607 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n8606 = ~n8605 | ~n8604;
  assign n8615 = ~n8607 & ~n8606;
  assign n8609 = ~n9672 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n8608 = ~n9665 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n8613 = ~n8609 | ~n8608;
  assign n8611 = ~n9636 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n8610 = ~n9648 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n8612 = ~n8611 | ~n8610;
  assign n8614 = ~n8613 & ~n8612;
  assign n8619 = ~n8615 | ~n8614;
  assign n8617 = ~n9522 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n8616 = ~n9657 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n8618 = ~n8617 | ~n8616;
  assign n8620 = ~n8619 & ~n8618;
  assign n8623 = ~EAX_REG_17__SCAN_IN;
  assign n8625 = ~n9708 | ~PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n8632 = ~n7003 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n8631 = ~n9653 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n8636 = ~n8632 | ~n8631;
  assign n8634 = ~n9607 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n8633 = ~n9662 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n8635 = ~n8634 | ~n8633;
  assign n8644 = ~n8636 & ~n8635;
  assign n8638 = ~n9656 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n8637 = ~n9665 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n8642 = ~n8638 | ~n8637;
  assign n8640 = ~n9647 | ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n8639 = ~n9522 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n8641 = ~n8640 | ~n8639;
  assign n8643 = ~n8642 & ~n8641;
  assign n8646 = ~n9599 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n8645 = ~n9636 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n8650 = ~n8646 | ~n8645;
  assign n8648 = ~n9610 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n8647 = ~n9602 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n8649 = ~n8648 | ~n8647;
  assign n8658 = ~n8650 & ~n8649;
  assign n8652 = ~n9673 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n8651 = ~n9648 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n8656 = ~n8652 | ~n8651;
  assign n8654 = ~n9501 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n8653 = ~n9672 | ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n8655 = ~n8654 | ~n8653;
  assign n8657 = ~n8656 & ~n8655;
  assign n8661 = ~n8660 & ~n8659;
  assign n8669 = n8661 | n9067;
  assign n8662 = ~EAX_REG_18__SCAN_IN;
  assign n8665 = ~n9708 | ~PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n8672 = ~n9501 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n8671 = ~n9610 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n8676 = ~n8672 | ~n8671;
  assign n8674 = ~n9673 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n8673 = ~n9636 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n8675 = ~n8674 | ~n8673;
  assign n8684 = ~n8676 & ~n8675;
  assign n8678 = ~n9672 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n8677 = ~n9607 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n8682 = ~n8678 | ~n8677;
  assign n8680 = ~n9522 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n8679 = ~n9653 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n8681 = ~n8680 | ~n8679;
  assign n8683 = ~n8682 & ~n8681;
  assign n8700 = ~n8684 | ~n8683;
  assign n8686 = ~n9656 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n8685 = ~n9599 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n8690 = ~n8686 | ~n8685;
  assign n8688 = ~n9647 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n8687 = ~n9657 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n8689 = ~n8688 | ~n8687;
  assign n8698 = ~n8690 & ~n8689;
  assign n8692 = ~n9602 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n8691 = ~n9662 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n8696 = ~n8692 | ~n8691;
  assign n8694 = ~n9665 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n8693 = ~n9648 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n8695 = ~n8694 | ~n8693;
  assign n8697 = ~n8696 & ~n8695;
  assign n8699 = ~n8698 | ~n8697;
  assign n8701 = ~n8700 & ~n8699;
  assign n8706 = n8701 | n9067;
  assign n8702 = ~n11478 & ~PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n8704 = ~STATE2_REG_2__SCAN_IN & ~n8702;
  assign n8713 = ~n9501 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n8712 = ~n9610 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n8717 = ~n8713 | ~n8712;
  assign n8715 = ~n9647 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n8714 = ~n9607 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n8716 = ~n8715 | ~n8714;
  assign n8725 = ~n8717 & ~n8716;
  assign n8719 = ~n7003 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n8718 = ~n9662 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n8723 = ~n8719 | ~n8718;
  assign n8721 = ~n9599 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n8720 = ~n9636 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n8722 = ~n8721 | ~n8720;
  assign n8724 = ~n8723 & ~n8722;
  assign n8741 = ~n8725 | ~n8724;
  assign n8727 = ~n9673 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n8726 = ~n9665 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n8731 = ~n8727 | ~n8726;
  assign n8729 = ~n9656 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n8728 = ~n9522 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n8730 = ~n8729 | ~n8728;
  assign n8739 = ~n8731 & ~n8730;
  assign n8733 = ~n9672 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n8732 = ~n9648 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n8737 = ~n8733 | ~n8732;
  assign n8735 = ~n9602 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n8734 = ~n9653 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n8736 = ~n8735 | ~n8734;
  assign n8738 = ~n8737 & ~n8736;
  assign n8740 = ~n8739 | ~n8738;
  assign n8742 = ~n8741 & ~n8740;
  assign n8748 = n8742 | n9067;
  assign n8743 = ~EAX_REG_20__SCAN_IN;
  assign n8744 = ~n11497 | ~PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n8753 = ~n9673 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n8752 = ~n9665 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n8757 = ~n8753 | ~n8752;
  assign n8755 = ~n9599 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n8754 = ~n9610 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n8756 = ~n8755 | ~n8754;
  assign n8765 = ~n8757 & ~n8756;
  assign n8759 = ~n9636 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n8758 = ~n9662 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n8763 = ~n8759 | ~n8758;
  assign n8761 = ~n9501 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n8760 = ~n9656 | ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n8762 = ~n8761 | ~n8760;
  assign n8764 = ~n8763 & ~n8762;
  assign n8781 = ~n8765 | ~n8764;
  assign n8767 = ~n9602 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n8766 = ~n9648 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n8771 = ~n8767 | ~n8766;
  assign n8769 = ~n7003 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n8768 = ~n9607 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n8770 = ~n8769 | ~n8768;
  assign n8779 = ~n8771 & ~n8770;
  assign n8773 = ~n9672 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n8772 = ~n9647 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n8777 = ~n8773 | ~n8772;
  assign n8775 = ~n9522 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n8774 = ~n9653 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n8776 = ~n8775 | ~n8774;
  assign n8778 = ~n8777 & ~n8776;
  assign n8780 = ~n8779 | ~n8778;
  assign n8782 = ~n8781 & ~n8780;
  assign n8788 = n8782 | n9067;
  assign n8784 = ~n11497 | ~PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n8785 = ~n9789 | ~n8784;
  assign n8793 = ~n8792 | ~n8791;
  assign n13177 = ~n13178 & ~n8793;
  assign n8797 = ~n13178 | ~EAX_REG_21__SCAN_IN;
  assign U2870 = n8800 | n8799;
  assign n8805 = ~n8804 | ~n8803;
  assign n12208 = ~n11402 & ~n11401;
  assign n11887 = ~n11553 & ~n11552;
  assign n10987 = ~n10865 & ~n10864;
  assign n11238 = ~n11087 & ~n11086;
  assign n8967 = ~n12696 & ~n12695;
  assign n8886 = ~n8967 | ~n8966;
  assign U2838 = n8890 | n8889;
  assign n8894 = ~n9636 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n8893 = ~n9662 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n8898 = ~n8894 | ~n8893;
  assign n8896 = ~n9647 | ~INSTQUEUE_REG_0__6__SCAN_IN;
  assign n8895 = ~n9653 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n8897 = ~n8896 | ~n8895;
  assign n8906 = ~n8898 & ~n8897;
  assign n8900 = ~n9501 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n8899 = ~n9602 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n8904 = ~n8900 | ~n8899;
  assign n8902 = ~n9656 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n8901 = ~n9648 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n8903 = ~n8902 | ~n8901;
  assign n8905 = ~n8904 & ~n8903;
  assign n8922 = ~n8906 | ~n8905;
  assign n8908 = ~n9610 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n8907 = ~n9607 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n8912 = ~n8908 | ~n8907;
  assign n8910 = ~n9672 | ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n8909 = ~n9522 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n8911 = ~n8910 | ~n8909;
  assign n8920 = ~n8912 & ~n8911;
  assign n8914 = ~n7003 | ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n8913 = ~n9665 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n8918 = ~n8914 | ~n8913;
  assign n8916 = ~n9599 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n8915 = ~n9673 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n8917 = ~n8916 | ~n8915;
  assign n8919 = ~n8918 & ~n8917;
  assign n8921 = ~n8920 | ~n8919;
  assign n8923 = ~n8922 & ~n8921;
  assign n8929 = n8923 | n9067;
  assign n8927 = ~n9686 & ~n8924;
  assign n8925 = ~n11497 | ~PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n8926 = ~n9789 | ~n8925;
  assign n8934 = ~n8999;
  assign n8937 = ~n13178 | ~EAX_REG_22__SCAN_IN;
  assign U2869 = n8940 | n8939;
  assign n8961 = ~REIP_REG_18__SCAN_IN | ~REIP_REG_17__SCAN_IN;
  assign n9951 = ~REIP_REG_14__SCAN_IN;
  assign n12603 = ~REIP_REG_13__SCAN_IN;
  assign n12029 = ~n9951 & ~n12603;
  assign n12380 = ~REIP_REG_9__SCAN_IN;
  assign n12630 = ~REIP_REG_8__SCAN_IN;
  assign n11911 = ~n12380 & ~n12630;
  assign n11975 = ~REIP_REG_10__SCAN_IN | ~n11911;
  assign n8941 = ~REIP_REG_12__SCAN_IN | ~REIP_REG_11__SCAN_IN;
  assign n12447 = ~REIP_REG_6__SCAN_IN;
  assign n9994 = ~REIP_REG_4__SCAN_IN;
  assign n11654 = ~REIP_REG_3__SCAN_IN | ~REIP_REG_2__SCAN_IN;
  assign n8942 = ~n10574 | ~n9855;
  assign n8955 = ~n10937 | ~n8942;
  assign n9091 = ~n8949;
  assign n10061 = n8951 & n10038;
  assign n8952 = ~n13491 & ~n10061;
  assign n11630 = n11654 | n12577;
  assign n12651 = ~n9994 & ~n11630;
  assign n12631 = ~n12418 & ~n12427;
  assign n9984 = ~REIP_REG_1__SCAN_IN;
  assign n8956 = ~n9984 & ~n11654;
  assign n8957 = ~REIP_REG_4__SCAN_IN | ~n8956;
  assign n8995 = n8962 | n12721;
  assign n13330 = ~n8989 & ~n8988;
  assign n8977 = ~n8973;
  assign n8982 = ~n8978 & ~n10240;
  assign n8979 = ~n9092 & ~EBX_REG_31__SCAN_IN;
  assign n8981 = n8980 & n8979;
  assign n8983 = ~n8982 & ~n8981;
  assign n13197 = ~n8989 & ~n13471;
  assign U2807 = n8997 | n8996;
  assign n9078 = ~n9080;
  assign n9001 = ~n9673 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n9000 = ~n9607 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n9005 = ~n9001 | ~n9000;
  assign n9003 = ~n9599 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n9002 = ~n9636 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n9004 = ~n9003 | ~n9002;
  assign n9029 = ~n9005 & ~n9004;
  assign n9007 = ~n9522 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n9006 = ~n9602 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n9011 = ~n9007 | ~n9006;
  assign n9009 = ~n9501 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n9008 = ~n9653 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n9010 = ~n9009 | ~n9008;
  assign n9019 = ~n9011 & ~n9010;
  assign n9013 = ~n9656 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n9012 = ~n7003 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n9017 = ~n9013 | ~n9012;
  assign n9015 = ~n9665 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n9014 = ~n9662 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n9016 = ~n9015 | ~n9014;
  assign n9018 = ~n9017 & ~n9016;
  assign n9027 = ~n9019 | ~n9018;
  assign n9021 = ~n9672 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n9020 = ~n9647 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n9025 = ~n9021 | ~n9020;
  assign n9023 = ~n9610 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n9022 = ~n9648 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n9024 = ~n9023 | ~n9022;
  assign n9026 = n9025 | n9024;
  assign n9028 = ~n9027 & ~n9026;
  assign n9031 = ~n9673 | ~INSTQUEUE_REG_11__0__SCAN_IN;
  assign n9030 = ~n9662 | ~INSTQUEUE_REG_4__0__SCAN_IN;
  assign n9035 = ~n9031 | ~n9030;
  assign n9033 = ~n9602 | ~INSTQUEUE_REG_5__0__SCAN_IN;
  assign n9032 = ~n9665 | ~INSTQUEUE_REG_12__0__SCAN_IN;
  assign n9034 = ~n9033 | ~n9032;
  assign n9066 = ~n9035 & ~n9034;
  assign n9037 = ~n9599 | ~INSTQUEUE_REG_13__0__SCAN_IN;
  assign n9036 = ~n9653 | ~INSTQUEUE_REG_7__0__SCAN_IN;
  assign n9041 = ~n9037 | ~n9036;
  assign n9039 = ~n9656 | ~INSTQUEUE_REG_10__0__SCAN_IN;
  assign n9038 = ~n9648 | ~INSTQUEUE_REG_8__0__SCAN_IN;
  assign n9040 = ~n9039 | ~n9038;
  assign n9049 = ~n9041 & ~n9040;
  assign n9043 = ~n9647 | ~INSTQUEUE_REG_1__0__SCAN_IN;
  assign n9042 = ~n9522 | ~INSTQUEUE_REG_2__0__SCAN_IN;
  assign n9047 = ~n9043 | ~n9042;
  assign n9045 = ~n9501 | ~INSTQUEUE_REG_14__0__SCAN_IN;
  assign n9044 = ~n9672 | ~INSTQUEUE_REG_9__0__SCAN_IN;
  assign n9046 = ~n9045 | ~n9044;
  assign n9048 = ~n9047 & ~n9046;
  assign n9064 = ~n9049 | ~n9048;
  assign n9055 = ~n9051 & ~n9050;
  assign n9054 = ~n9053 & ~n9052;
  assign n9062 = ~n9055 & ~n9054;
  assign n9060 = ~n9057 & ~n9056;
  assign n9059 = ~n9642 & ~n9058;
  assign n9061 = ~n9060 & ~n9059;
  assign n9063 = ~n9062 | ~n9061;
  assign n9065 = ~n9064 & ~n9063;
  assign n9068 = ~n9210 ^ n9209;
  assign n9076 = n9068 | n9067;
  assign n9069 = ~EAX_REG_23__SCAN_IN;
  assign n9072 = ~n9708 | ~PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n9084 = ~n13178 | ~EAX_REG_23__SCAN_IN;
  assign U2868 = n9087 | n9086;
  assign n11406 = ~n11325 & ~n11432;
  assign n9119 = ~n12202 & ~n12196;
  assign n11557 = ~n11406 | ~n9119;
  assign n11920 = ~n11893 & ~n9088;
  assign n12500 = ~n12501 & ~n12502;
  assign n12513 = ~n11920 | ~n12500;
  assign n12519 = ~n11557 & ~n12513;
  assign n12774 = ~n12771 & ~n12770;
  assign n9089 = ~n10515 & ~n9855;
  assign n9090 = ~n9089 & ~READY_N;
  assign n9104 = n9100 | n10245;
  assign n9109 = n9108 | n9107;
  assign n9125 = ~n9109 | ~n12691;
  assign n13043 = ~n9161 | ~n10077;
  assign n9112 = ~n9111 & ~n9110;
  assign n9113 = ~n9112 & ~n10574;
  assign n9115 = n9114 | n9113;
  assign n11324 = ~n9161 | ~n9115;
  assign n11579 = ~n9116 & ~n13250;
  assign n9118 = ~n8001 & ~n11578;
  assign n11569 = ~n9118 & ~INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n11407 = ~n11569 & ~n11432;
  assign n12520 = ~n12513 & ~n11558;
  assign n12836 = n9121 | n9120;
  assign n9348 = ~INSTADDRPOINTER_REG_14__SCAN_IN | ~INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n9357 = ~n12754 & ~n9348;
  assign n9360 = ~n9348 & ~n12755;
  assign n9123 = ~n13045 & ~n9360;
  assign n13377 = ~n11326 | ~n9127;
  assign n9157 = ~n9131;
  assign n9133 = ~n9157 | ~n9132;
  assign n9137 = ~n9134 | ~n9133;
  assign n9136 = ~n9135;
  assign n9141 = n9161 & n9140;
  assign n9145 = ~n9143 | ~n9142;
  assign n9152 = ~n9145 | ~n9144;
  assign n9149 = ~n9152;
  assign n12830 = ~n9331 | ~n9153;
  assign n9154 = ~n12826;
  assign n9159 = ~n9156;
  assign n9158 = ~n9157 | ~n7231;
  assign n9164 = n9163 & n9162;
  assign U3003 = n9168 | n9167;
  assign n9170 = ~n9169 | ~REIP_REG_20__SCAN_IN;
  assign n9311 = ~REIP_REG_21__SCAN_IN | ~REIP_REG_20__SCAN_IN;
  assign U2806 = n9183 | n9182;
  assign n9189 = ~n13335 | ~EBX_REG_23__SCAN_IN;
  assign n9188 = ~n13334 | ~PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n9193 = ~n10937 | ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n9199 = ~n9316 | ~n9315;
  assign n9196 = ~n10937 | ~INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n12875 = ~n9199 & ~n9198;
  assign U2804 = n9207 | n9206;
  assign n9212 = ~n9636 | ~INSTQUEUE_REG_6__1__SCAN_IN;
  assign n9211 = ~n9607 | ~INSTQUEUE_REG_0__1__SCAN_IN;
  assign n9216 = ~n9212 | ~n9211;
  assign n9214 = ~n9672 | ~INSTQUEUE_REG_9__1__SCAN_IN;
  assign n9213 = ~n9610 | ~INSTQUEUE_REG_15__1__SCAN_IN;
  assign n9215 = ~n9214 | ~n9213;
  assign n9224 = ~n9216 & ~n9215;
  assign n9218 = ~n9647 | ~INSTQUEUE_REG_1__1__SCAN_IN;
  assign n9217 = ~n9602 | ~INSTQUEUE_REG_5__1__SCAN_IN;
  assign n9222 = ~n9218 | ~n9217;
  assign n9220 = ~n9656 | ~INSTQUEUE_REG_10__1__SCAN_IN;
  assign n9219 = ~n9522 | ~INSTQUEUE_REG_2__1__SCAN_IN;
  assign n9221 = ~n9220 | ~n9219;
  assign n9223 = ~n9222 & ~n9221;
  assign n9240 = ~n9224 | ~n9223;
  assign n9226 = ~n9501 | ~INSTQUEUE_REG_14__1__SCAN_IN;
  assign n9225 = ~n9599 | ~INSTQUEUE_REG_13__1__SCAN_IN;
  assign n9230 = ~n9226 | ~n9225;
  assign n9228 = ~n9657 | ~INSTQUEUE_REG_3__1__SCAN_IN;
  assign n9227 = ~n9653 | ~INSTQUEUE_REG_7__1__SCAN_IN;
  assign n9229 = ~n9228 | ~n9227;
  assign n9238 = ~n9230 & ~n9229;
  assign n9232 = ~n9665 | ~INSTQUEUE_REG_12__1__SCAN_IN;
  assign n9231 = ~n9648 | ~INSTQUEUE_REG_8__1__SCAN_IN;
  assign n9236 = ~n9232 | ~n9231;
  assign n9234 = ~n9673 | ~INSTQUEUE_REG_11__1__SCAN_IN;
  assign n9233 = ~n9662 | ~INSTQUEUE_REG_4__1__SCAN_IN;
  assign n9235 = ~n9234 | ~n9233;
  assign n9237 = ~n9236 & ~n9235;
  assign n9239 = ~n9238 | ~n9237;
  assign n9260 = ~n9240 & ~n9239;
  assign n9241 = n9259 ^ n9260;
  assign n9242 = ~EAX_REG_24__SCAN_IN;
  assign n9245 = ~n9686 & ~n9242;
  assign n9243 = ~PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n9244 = ~n9535 & ~n9243;
  assign n9246 = ~n9245 & ~n9244;
  assign n9255 = ~n13178 | ~EAX_REG_24__SCAN_IN;
  assign U2867 = n9258 | n9257;
  assign n9262 = ~n9673 | ~INSTQUEUE_REG_11__2__SCAN_IN;
  assign n9261 = ~n9647 | ~INSTQUEUE_REG_1__2__SCAN_IN;
  assign n9266 = ~n9262 | ~n9261;
  assign n9264 = ~n9501 | ~INSTQUEUE_REG_14__2__SCAN_IN;
  assign n9263 = ~n9607 | ~INSTQUEUE_REG_0__2__SCAN_IN;
  assign n9265 = ~n9264 | ~n9263;
  assign n9270 = n9266 | n9265;
  assign n9268 = ~n9656 | ~INSTQUEUE_REG_10__2__SCAN_IN;
  assign n9267 = ~n9610 | ~INSTQUEUE_REG_15__2__SCAN_IN;
  assign n9269 = ~n9268 | ~n9267;
  assign n9290 = ~n9270 & ~n9269;
  assign n9272 = ~n9599 | ~INSTQUEUE_REG_13__2__SCAN_IN;
  assign n9271 = ~n9653 | ~INSTQUEUE_REG_7__2__SCAN_IN;
  assign n9276 = ~n9272 | ~n9271;
  assign n9274 = ~n9636 | ~INSTQUEUE_REG_6__2__SCAN_IN;
  assign n9273 = ~n9662 | ~INSTQUEUE_REG_4__2__SCAN_IN;
  assign n9275 = ~n9274 | ~n9273;
  assign n9284 = ~n9276 & ~n9275;
  assign n9278 = ~n9522 | ~INSTQUEUE_REG_2__2__SCAN_IN;
  assign n9277 = ~n9648 | ~INSTQUEUE_REG_8__2__SCAN_IN;
  assign n9282 = ~n9278 | ~n9277;
  assign n9280 = ~n9672 | ~INSTQUEUE_REG_9__2__SCAN_IN;
  assign n9279 = ~n9602 | ~INSTQUEUE_REG_5__2__SCAN_IN;
  assign n9281 = ~n9280 | ~n9279;
  assign n9283 = ~n9282 & ~n9281;
  assign n9288 = ~n9284 | ~n9283;
  assign n9286 = ~n9657 | ~INSTQUEUE_REG_3__2__SCAN_IN;
  assign n9285 = ~n9665 | ~INSTQUEUE_REG_12__2__SCAN_IN;
  assign n9287 = ~n9286 | ~n9285;
  assign n9289 = ~n9288 & ~n9287;
  assign n9291 = n9418 ^ n9417;
  assign n9294 = ~n9707 | ~EAX_REG_25__SCAN_IN;
  assign n9292 = ~n8970 & ~STATE2_REG_2__SCAN_IN;
  assign n9293 = ~n9292 & ~n9698;
  assign n9307 = ~n13178 | ~EAX_REG_25__SCAN_IN;
  assign U2866 = n9310 | n9309;
  assign n9312 = REIP_REG_22__SCAN_IN | n9311;
  assign U2805 = n9328 | n9327;
  assign n9335 = ~n9331 | ~n9330;
  assign n12889 = ~n9335 | ~n9333;
  assign n9336 = ~n9335 & ~n9334;
  assign n9341 = ~n9340;
  assign n9356 = ~INSTADDRPOINTER_REG_16__SCAN_IN | ~INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n9351 = ~n9348;
  assign n9350 = ~n9375 | ~n9349;
  assign n9352 = n9351 & n9350;
  assign n9353 = ~n9356 | ~n9352;
  assign U3002 = n9355 | n9354;
  assign n13272 = ~INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n13484 = ~n13481 & ~n13480;
  assign n12998 = ~n9356;
  assign n9558 = ~n9357 | ~n12998;
  assign n13048 = ~n9558 & ~n13112;
  assign n13053 = ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n9561 = ~n13257 & ~n13053;
  assign n13372 = ~n13048 | ~n9561;
  assign n13410 = ~INSTADDRPOINTER_REG_22__SCAN_IN | ~INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n9555 = ~n13372 & ~n13410;
  assign n9776 = ~n13272 & ~n9366;
  assign n9359 = ~n13043 & ~n9776;
  assign n9358 = ~n11324 & ~n9555;
  assign n9362 = ~n9359 & ~n9358;
  assign n9559 = ~n12998 | ~n9360;
  assign n13044 = ~n13112 & ~n9559;
  assign n13373 = ~n9561 | ~n13044;
  assign n9367 = ~n13410 & ~n13373;
  assign n13274 = ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n9772 = ~n13484 | ~n9367;
  assign n13501 = n9369 | n9368;
  assign n9371 = ~n9773;
  assign n9370 = ~INSTADDRPOINTER_REG_25__SCAN_IN & ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n9372 = ~n9371 & ~n9370;
  assign n13109 = ~INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n13002 = ~INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n9567 = ~n12889 & ~n9373;
  assign n9379 = ~n9567 | ~n9374;
  assign n13111 = ~n13002 | ~n13109;
  assign n9376 = ~INSTADDRPOINTER_REG_19__SCAN_IN & ~n13111;
  assign n9377 = ~n9376 | ~n9375;
  assign n13270 = ~n9379 | ~n9378;
  assign n9380 = ~n13484 | ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n13283 = ~n13257 & ~n9380;
  assign n13370 = ~INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n9406 = ~n9386 | ~n9385;
  assign n9390 = ~n10937 | ~INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n12883 = ~n12875 | ~n12874;
  assign n9393 = ~n10937 | ~INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n9714 = ~n12883 & ~n12882;
  assign n9396 = ~n10937 | ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n9395 = ~n10932 | ~EBX_REG_26__SCAN_IN;
  assign U2992 = n9403 | n9402;
  assign n13244 = ~n9409 | ~n9408;
  assign n9410 = ~INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n13239 = ~n13244 | ~n13240;
  assign n9415 = ~n13239 | ~n9411;
  assign n9780 = ~INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n9412 = ~n13434 & ~n9780;
  assign n9420 = ~n9501 | ~INSTQUEUE_REG_14__3__SCAN_IN;
  assign n9419 = ~n9672 | ~INSTQUEUE_REG_9__3__SCAN_IN;
  assign n9424 = ~n9420 | ~n9419;
  assign n9422 = ~n9599 | ~INSTQUEUE_REG_13__3__SCAN_IN;
  assign n9421 = ~n9665 | ~INSTQUEUE_REG_12__3__SCAN_IN;
  assign n9423 = ~n9422 | ~n9421;
  assign n9432 = ~n9424 & ~n9423;
  assign n9426 = ~n9522 | ~INSTQUEUE_REG_2__3__SCAN_IN;
  assign n9425 = ~n9607 | ~INSTQUEUE_REG_0__3__SCAN_IN;
  assign n9430 = ~n9426 | ~n9425;
  assign n9428 = ~n9636 | ~INSTQUEUE_REG_6__3__SCAN_IN;
  assign n9427 = ~n9648 | ~INSTQUEUE_REG_8__3__SCAN_IN;
  assign n9429 = ~n9428 | ~n9427;
  assign n9431 = ~n9430 & ~n9429;
  assign n9448 = ~n9432 | ~n9431;
  assign n9434 = ~n9656 | ~INSTQUEUE_REG_10__3__SCAN_IN;
  assign n9433 = ~n9673 | ~INSTQUEUE_REG_11__3__SCAN_IN;
  assign n9438 = ~n9434 | ~n9433;
  assign n9436 = ~n9657 | ~INSTQUEUE_REG_3__3__SCAN_IN;
  assign n9435 = ~n9662 | ~INSTQUEUE_REG_4__3__SCAN_IN;
  assign n9437 = ~n9436 | ~n9435;
  assign n9446 = ~n9438 & ~n9437;
  assign n9440 = ~n9647 | ~INSTQUEUE_REG_1__3__SCAN_IN;
  assign n9439 = ~n9610 | ~INSTQUEUE_REG_15__3__SCAN_IN;
  assign n9444 = ~n9440 | ~n9439;
  assign n9442 = ~n9602 | ~INSTQUEUE_REG_5__3__SCAN_IN;
  assign n9441 = ~n9653 | ~INSTQUEUE_REG_7__3__SCAN_IN;
  assign n9443 = ~n9442 | ~n9441;
  assign n9445 = ~n9444 & ~n9443;
  assign n9447 = ~n9446 | ~n9445;
  assign n9458 = ~n9448 & ~n9447;
  assign n9449 = n9457 ^ n9458;
  assign n9450 = ~EAX_REG_26__SCAN_IN;
  assign n9452 = ~n9686 & ~n9450;
  assign n9451 = ~n9535 & ~n13163;
  assign n9453 = ~n9452 & ~n9451;
  assign n9460 = ~n9501 | ~INSTQUEUE_REG_14__4__SCAN_IN;
  assign n9459 = ~n9665 | ~INSTQUEUE_REG_12__4__SCAN_IN;
  assign n9464 = ~n9460 | ~n9459;
  assign n9462 = ~n9672 | ~INSTQUEUE_REG_9__4__SCAN_IN;
  assign n9461 = ~n9648 | ~INSTQUEUE_REG_8__4__SCAN_IN;
  assign n9463 = ~n9462 | ~n9461;
  assign n9488 = ~n9464 & ~n9463;
  assign n9466 = ~n7003 | ~INSTQUEUE_REG_3__4__SCAN_IN;
  assign n9465 = ~n9662 | ~INSTQUEUE_REG_4__4__SCAN_IN;
  assign n9470 = ~n9466 | ~n9465;
  assign n9468 = ~n9599 | ~INSTQUEUE_REG_13__4__SCAN_IN;
  assign n9467 = ~n9653 | ~INSTQUEUE_REG_7__4__SCAN_IN;
  assign n9469 = ~n9468 | ~n9467;
  assign n9478 = ~n9470 & ~n9469;
  assign n9472 = ~n9602 | ~INSTQUEUE_REG_5__4__SCAN_IN;
  assign n9471 = ~n9636 | ~INSTQUEUE_REG_6__4__SCAN_IN;
  assign n9476 = ~n9472 | ~n9471;
  assign n9474 = ~n9647 | ~INSTQUEUE_REG_1__4__SCAN_IN;
  assign n9473 = ~n9522 | ~INSTQUEUE_REG_2__4__SCAN_IN;
  assign n9475 = ~n9474 | ~n9473;
  assign n9477 = ~n9476 & ~n9475;
  assign n9486 = ~n9478 | ~n9477;
  assign n9480 = ~n9610 | ~INSTQUEUE_REG_15__4__SCAN_IN;
  assign n9479 = ~n9673 | ~INSTQUEUE_REG_11__4__SCAN_IN;
  assign n9484 = ~n9480 | ~n9479;
  assign n9482 = ~n9656 | ~INSTQUEUE_REG_10__4__SCAN_IN;
  assign n9481 = ~n9607 | ~INSTQUEUE_REG_0__4__SCAN_IN;
  assign n9483 = ~n9482 | ~n9481;
  assign n9485 = n9484 | n9483;
  assign n9487 = ~n9486 & ~n9485;
  assign n9499 = ~n9488 | ~n9487;
  assign n9489 = n9500 ^ n9499;
  assign n9495 = n9489 & n9696;
  assign n9493 = ~n9707 | ~EAX_REG_27__SCAN_IN;
  assign n9491 = ~n9490 & ~STATE2_REG_2__SCAN_IN;
  assign n9492 = ~n9491 & ~n9698;
  assign n9503 = ~n9501 | ~INSTQUEUE_REG_14__5__SCAN_IN;
  assign n9502 = ~n9665 | ~INSTQUEUE_REG_12__5__SCAN_IN;
  assign n9507 = ~n9503 | ~n9502;
  assign n9505 = ~n9647 | ~INSTQUEUE_REG_1__5__SCAN_IN;
  assign n9504 = ~n9662 | ~INSTQUEUE_REG_4__5__SCAN_IN;
  assign n9506 = ~n9505 | ~n9504;
  assign n9515 = ~n9507 & ~n9506;
  assign n9509 = ~n9657 | ~INSTQUEUE_REG_3__5__SCAN_IN;
  assign n9508 = ~n9602 | ~INSTQUEUE_REG_5__5__SCAN_IN;
  assign n9513 = ~n9509 | ~n9508;
  assign n9511 = ~n9607 | ~INSTQUEUE_REG_0__5__SCAN_IN;
  assign n9510 = ~n9653 | ~INSTQUEUE_REG_7__5__SCAN_IN;
  assign n9512 = ~n9511 | ~n9510;
  assign n9514 = ~n9513 & ~n9512;
  assign n9532 = ~n9515 | ~n9514;
  assign n9517 = ~n9672 | ~INSTQUEUE_REG_9__5__SCAN_IN;
  assign n9516 = ~n9648 | ~INSTQUEUE_REG_8__5__SCAN_IN;
  assign n9521 = ~n9517 | ~n9516;
  assign n9519 = ~n9599 | ~INSTQUEUE_REG_13__5__SCAN_IN;
  assign n9518 = ~n9636 | ~INSTQUEUE_REG_6__5__SCAN_IN;
  assign n9520 = ~n9519 | ~n9518;
  assign n9530 = ~n9521 & ~n9520;
  assign n9524 = ~n9522 | ~INSTQUEUE_REG_2__5__SCAN_IN;
  assign n9523 = ~n9673 | ~INSTQUEUE_REG_11__5__SCAN_IN;
  assign n9528 = ~n9524 | ~n9523;
  assign n9526 = ~n9656 | ~INSTQUEUE_REG_10__5__SCAN_IN;
  assign n9525 = ~n9610 | ~INSTQUEUE_REG_15__5__SCAN_IN;
  assign n9527 = ~n9526 | ~n9525;
  assign n9529 = ~n9528 & ~n9527;
  assign n9531 = ~n9530 | ~n9529;
  assign n9635 = ~n9532 & ~n9531;
  assign n9533 = n9634 ^ n9635;
  assign n9542 = n9533 & n9696;
  assign n9534 = ~PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n9538 = ~n9535 & ~n9534;
  assign n13132 = ~n13092 & ~n9546;
  assign n9547 = ~n13467 | ~PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n9550 = ~n9766 | ~n9547;
  assign n13133 = ~n9548;
  assign n9549 = ~n13316 & ~n13133;
  assign U2958 = n9554 | n9553;
  assign n9556 = n13049 | n9555;
  assign n9565 = ~INSTADDRPOINTER_REG_16__SCAN_IN & ~n13111;
  assign n9571 = ~n9569 | ~n9568;
  assign n13077 = ~n9571 | ~n9570;
  assign n13414 = ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n9740 = ~n9574 | ~n13217;
  assign n13314 = ~n13491 | ~REIP_REG_23__SCAN_IN;
  assign n9581 = ~n13314;
  assign U2995 = n9586 | n9585;
  assign n13026 = ~REIP_REG_25__SCAN_IN | ~REIP_REG_26__SCAN_IN;
  assign n13126 = ~REIP_REG_27__SCAN_IN;
  assign n9587 = n13026 | n13126;
  assign n9888 = ~REIP_REG_30__SCAN_IN;
  assign n13200 = ~REIP_REG_29__SCAN_IN;
  assign n9594 = ~n9888 & ~n13200;
  assign n9590 = n12929 | n9594;
  assign n9592 = ~n13026;
  assign n9593 = ~REIP_REG_28__SCAN_IN | ~REIP_REG_27__SCAN_IN;
  assign n9601 = ~n9599 | ~INSTQUEUE_REG_13__7__SCAN_IN;
  assign n9600 = ~n9636 | ~INSTQUEUE_REG_6__7__SCAN_IN;
  assign n9606 = ~n9601 | ~n9600;
  assign n9604 = ~n9602 | ~INSTQUEUE_REG_5__7__SCAN_IN;
  assign n9603 = ~n9653 | ~INSTQUEUE_REG_7__7__SCAN_IN;
  assign n9605 = ~n9604 | ~n9603;
  assign n9616 = ~n9606 & ~n9605;
  assign n9609 = ~n9656 | ~INSTQUEUE_REG_10__7__SCAN_IN;
  assign n9608 = ~n9607 | ~INSTQUEUE_REG_0__7__SCAN_IN;
  assign n9614 = ~n9609 | ~n9608;
  assign n9612 = ~n9501 | ~INSTQUEUE_REG_14__7__SCAN_IN;
  assign n9611 = ~n9610 | ~INSTQUEUE_REG_15__7__SCAN_IN;
  assign n9613 = ~n9612 | ~n9611;
  assign n9615 = ~n9614 & ~n9613;
  assign n9632 = ~n9616 | ~n9615;
  assign n9618 = ~n9672 | ~INSTQUEUE_REG_9__7__SCAN_IN;
  assign n9617 = ~n9647 | ~INSTQUEUE_REG_1__7__SCAN_IN;
  assign n9622 = ~n9618 | ~n9617;
  assign n9620 = ~n9522 | ~INSTQUEUE_REG_2__7__SCAN_IN;
  assign n9619 = ~n9673 | ~INSTQUEUE_REG_11__7__SCAN_IN;
  assign n9621 = ~n9620 | ~n9619;
  assign n9630 = ~n9622 & ~n9621;
  assign n9624 = ~n9665 | ~INSTQUEUE_REG_12__7__SCAN_IN;
  assign n9623 = ~n9662 | ~INSTQUEUE_REG_4__7__SCAN_IN;
  assign n9628 = ~n9624 | ~n9623;
  assign n9626 = ~n7003 | ~INSTQUEUE_REG_3__7__SCAN_IN;
  assign n9625 = ~n9648 | ~INSTQUEUE_REG_8__7__SCAN_IN;
  assign n9627 = ~n9626 | ~n9625;
  assign n9629 = ~n9628 & ~n9627;
  assign n9631 = ~n9630 | ~n9629;
  assign n9682 = ~n9632 & ~n9631;
  assign n9681 = ~n9682 | ~n9633;
  assign n9695 = ~n9635 & ~n9634;
  assign n9638 = ~n9610 | ~INSTQUEUE_REG_15__6__SCAN_IN;
  assign n9637 = ~n9636 | ~INSTQUEUE_REG_6__6__SCAN_IN;
  assign n9646 = n9638 & n9637;
  assign n9639 = ~INSTQUEUE_REG_2__6__SCAN_IN;
  assign n9644 = ~n9640 & ~n9639;
  assign n9643 = ~n9642 & ~n9641;
  assign n9645 = ~n9644 & ~n9643;
  assign n9652 = ~n9646 | ~n9645;
  assign n9650 = ~n9647 | ~INSTQUEUE_REG_1__6__SCAN_IN;
  assign n9649 = ~n9648 | ~INSTQUEUE_REG_8__6__SCAN_IN;
  assign n9651 = ~n9650 | ~n9649;
  assign n9679 = ~n9652 & ~n9651;
  assign n9655 = ~n9602 | ~INSTQUEUE_REG_5__6__SCAN_IN;
  assign n9654 = ~n9653 | ~INSTQUEUE_REG_7__6__SCAN_IN;
  assign n9661 = ~n9655 | ~n9654;
  assign n9659 = ~n9656 | ~INSTQUEUE_REG_10__6__SCAN_IN;
  assign n9658 = ~n7003 | ~INSTQUEUE_REG_3__6__SCAN_IN;
  assign n9660 = ~n9659 | ~n9658;
  assign n9671 = ~n9661 & ~n9660;
  assign n9664 = ~n9501 | ~INSTQUEUE_REG_14__6__SCAN_IN;
  assign n9663 = ~n9662 | ~INSTQUEUE_REG_4__6__SCAN_IN;
  assign n9669 = ~n9664 | ~n9663;
  assign n9667 = ~n9599 | ~INSTQUEUE_REG_13__6__SCAN_IN;
  assign n9666 = ~n9665 | ~INSTQUEUE_REG_12__6__SCAN_IN;
  assign n9668 = ~n9667 | ~n9666;
  assign n9670 = ~n9669 & ~n9668;
  assign n9677 = ~n9671 | ~n9670;
  assign n9675 = ~n9672 | ~INSTQUEUE_REG_9__6__SCAN_IN;
  assign n9674 = ~n9673 | ~INSTQUEUE_REG_11__6__SCAN_IN;
  assign n9676 = ~n9675 | ~n9674;
  assign n9678 = ~n9677 & ~n9676;
  assign n9694 = ~n9679 | ~n9678;
  assign n9683 = ~n9695 | ~n9694;
  assign n9680 = ~n9683 | ~n9696;
  assign n9685 = ~n9681 | ~n9680;
  assign n9684 = ~n9683 | ~n9682;
  assign n9691 = ~n9685 | ~n9684;
  assign n9689 = ~n9686 & ~n10441;
  assign n9687 = ~n11497 | ~PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n9688 = ~n9789 | ~n9687;
  assign n9690 = ~n9689 & ~n9688;
  assign n9697 = n9695 ^ n9694;
  assign n9703 = n9697 & n9696;
  assign n9701 = ~n9707 | ~EAX_REG_29__SCAN_IN;
  assign n9699 = ~n8971 & ~STATE2_REG_2__SCAN_IN;
  assign n9700 = ~n9699 & ~n9698;
  assign n9702 = ~n9701 | ~n9700;
  assign n9706 = ~n9703 & ~n9702;
  assign n13174 = ~n13092 | ~n13091;
  assign n9712 = ~n13175 & ~n13174;
  assign n9710 = ~n9707 | ~EAX_REG_31__SCAN_IN;
  assign n9709 = ~n9708 | ~PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n13464 = n9712 ^ n9711;
  assign n12971 = ~n9714 | ~n9713;
  assign n9716 = ~n10937 | ~INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n9715 = ~n10932 | ~EBX_REG_27__SCAN_IN;
  assign n9761 = ~n12971 & ~n12970;
  assign n9719 = ~n10937 | ~INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n9718 = ~n10932 | ~EBX_REG_28__SCAN_IN;
  assign n9720 = ~n9719 | ~n9718;
  assign n13187 = ~n9761 | ~n9762;
  assign n9722 = ~n10937 | ~INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n9721 = ~n10932 | ~EBX_REG_29__SCAN_IN;
  assign n13103 = ~n13102 | ~n13101;
  assign n9725 = ~n10937 | ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n9724 = ~n10932 | ~EBX_REG_30__SCAN_IN;
  assign n9729 = ~n10937 | ~INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n9728 = ~n10932 | ~EBX_REG_31__SCAN_IN;
  assign n9730 = ~n9729 | ~n9728;
  assign n9733 = ~n13334 | ~PHYADDRPOINTER_REG_31__SCAN_IN;
  assign U2796 = n9739 | n9738;
  assign n9742 = ~n9740 | ~n13271;
  assign n9746 = ~n13347 | ~n13346;
  assign n9750 = ~n9746 | ~n9745;
  assign n9751 = ~n13467 | ~PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n9753 = ~n13508 | ~n9751;
  assign n9752 = ~n13316 & ~n12951;
  assign U2961 = n9757 | n9756;
  assign n13297 = ~INSTADDRPOINTER_REG_28__SCAN_IN | ~INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n13301 = ~n13297;
  assign n13273 = ~INSTADDRPOINTER_REG_27__SCAN_IN & ~INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n9759 = ~n13301 & ~n13273;
  assign n9763 = ~n9762;
  assign n9770 = ~n9769 & ~n9768;
  assign n9774 = ~n9773 & ~n9772;
  assign n9777 = ~n9776 | ~INSTADDRPOINTER_REG_26__SCAN_IN;
  assign U2990 = n9782 | n9781;
  assign n9783 = ~STATE_REG_1__SCAN_IN | ~n7393;
  assign n10023 = ~STATE_REG_0__SCAN_IN | ~n9783;
  assign n9784 = ~ADS_N_REG_SCAN_IN & ~n10023;
  assign n9861 = ~STATE_REG_0__SCAN_IN;
  assign U2789 = ~n9784 & ~n13515;
  assign n9786 = ~n11497 | ~n12680;
  assign n9785 = ~STATE2_REG_0__SCAN_IN | ~STATE2_REG_1__SCAN_IN;
  assign n9788 = ~n9786 & ~n9785;
  assign n9791 = ~n9788 & ~n9787;
  assign n9790 = ~n9789 | ~n10063;
  assign U3150 = ~n9791 | ~n9790;
  assign n13517 = ~n13515;
  assign n9793 = ~BE_N_REG_3__SCAN_IN | ~n13517;
  assign n9792 = ~BYTEENABLE_REG_3__SCAN_IN | ~n13515;
  assign U3445 = ~n9793 | ~n9792;
  assign n9795 = ~BE_N_REG_0__SCAN_IN | ~n13517;
  assign n9794 = ~BYTEENABLE_REG_0__SCAN_IN | ~n13515;
  assign U3448 = ~n9795 | ~n9794;
  assign n9797 = ~M_IO_N_REG_SCAN_IN | ~n13517;
  assign n9796 = ~MEMORYFETCH_REG_SCAN_IN | ~n13515;
  assign U3473 = ~n9797 | ~n9796;
  assign n9799 = ~BE_N_REG_2__SCAN_IN | ~n13517;
  assign n9798 = ~BYTEENABLE_REG_2__SCAN_IN | ~n13515;
  assign U3446 = ~n9799 | ~n9798;
  assign n9801 = ~BE_N_REG_1__SCAN_IN | ~n13517;
  assign n9800 = ~BYTEENABLE_REG_1__SCAN_IN | ~n13515;
  assign U3447 = ~n9801 | ~n9800;
  assign n9803 = ~DATAWIDTH_REG_30__SCAN_IN & ~DATAWIDTH_REG_31__SCAN_IN;
  assign n9802 = ~DATAWIDTH_REG_28__SCAN_IN & ~DATAWIDTH_REG_29__SCAN_IN;
  assign n9807 = ~n9803 | ~n9802;
  assign n9805 = ~DATAWIDTH_REG_18__SCAN_IN & ~DATAWIDTH_REG_19__SCAN_IN;
  assign n9804 = ~DATAWIDTH_REG_16__SCAN_IN & ~DATAWIDTH_REG_17__SCAN_IN;
  assign n9806 = ~n9805 | ~n9804;
  assign n9815 = ~n9807 & ~n9806;
  assign n9809 = ~DATAWIDTH_REG_26__SCAN_IN & ~DATAWIDTH_REG_27__SCAN_IN;
  assign n9808 = ~DATAWIDTH_REG_24__SCAN_IN & ~DATAWIDTH_REG_25__SCAN_IN;
  assign n9813 = ~n9809 | ~n9808;
  assign n9811 = ~DATAWIDTH_REG_22__SCAN_IN & ~DATAWIDTH_REG_23__SCAN_IN;
  assign n9810 = ~DATAWIDTH_REG_20__SCAN_IN & ~DATAWIDTH_REG_21__SCAN_IN;
  assign n9812 = ~n9811 | ~n9810;
  assign n9814 = ~n9813 & ~n9812;
  assign n9831 = ~n9815 | ~n9814;
  assign n9817 = ~DATAWIDTH_REG_14__SCAN_IN & ~DATAWIDTH_REG_15__SCAN_IN;
  assign n9816 = ~DATAWIDTH_REG_12__SCAN_IN & ~DATAWIDTH_REG_13__SCAN_IN;
  assign n9821 = ~n9817 | ~n9816;
  assign n9819 = ~DATAWIDTH_REG_3__SCAN_IN & ~DATAWIDTH_REG_2__SCAN_IN;
  assign n9818 = ~DATAWIDTH_REG_0__SCAN_IN | ~DATAWIDTH_REG_1__SCAN_IN;
  assign n9820 = ~n9819 | ~n9818;
  assign n9829 = ~n9821 & ~n9820;
  assign n9823 = ~DATAWIDTH_REG_10__SCAN_IN & ~DATAWIDTH_REG_11__SCAN_IN;
  assign n9822 = ~DATAWIDTH_REG_8__SCAN_IN & ~DATAWIDTH_REG_9__SCAN_IN;
  assign n9827 = ~n9823 | ~n9822;
  assign n9825 = ~DATAWIDTH_REG_6__SCAN_IN & ~DATAWIDTH_REG_7__SCAN_IN;
  assign n9824 = ~DATAWIDTH_REG_4__SCAN_IN & ~DATAWIDTH_REG_5__SCAN_IN;
  assign n9826 = ~n9825 | ~n9824;
  assign n9828 = ~n9827 & ~n9826;
  assign n9830 = ~n9829 | ~n9828;
  assign n9850 = ~n9831 & ~n9830;
  assign n9852 = ~n9850;
  assign n9839 = ~BYTEENABLE_REG_2__SCAN_IN | ~n9852;
  assign n9836 = ~REIP_REG_0__SCAN_IN | ~REIP_REG_1__SCAN_IN;
  assign n9849 = ~REIP_REG_0__SCAN_IN;
  assign n9833 = ~DATAWIDTH_REG_0__SCAN_IN | ~n9849;
  assign n9840 = ~DATAWIDTH_REG_1__SCAN_IN & ~DATAWIDTH_REG_0__SCAN_IN;
  assign n9832 = ~n9840;
  assign n9834 = ~n9833 | ~n9832;
  assign n9835 = ~n9834 | ~n9984;
  assign n9837 = ~n9836 | ~n9835;
  assign n9838 = ~n9837 | ~n9850;
  assign U3468 = ~n9839 | ~n9838;
  assign n9844 = ~BYTEENABLE_REG_3__SCAN_IN | ~n9852;
  assign n9841 = REIP_REG_1__SCAN_IN | DATAWIDTH_REG_1__SCAN_IN;
  assign n9845 = ~n9840 | ~n9849;
  assign n9842 = ~n9841 | ~n9845;
  assign n9843 = ~n9842 | ~n9850;
  assign U2795 = ~n9844 | ~n9843;
  assign n9846 = ~n9984 | ~n9845;
  assign n9848 = ~n9846 | ~n9850;
  assign n9847 = ~BYTEENABLE_REG_1__SCAN_IN | ~n9852;
  assign U2794 = ~n9848 | ~n9847;
  assign n9851 = ~n9984 | ~n9849;
  assign n9854 = ~n9851 | ~n9850;
  assign n9853 = ~BYTEENABLE_REG_0__SCAN_IN | ~n9852;
  assign U3469 = ~n9854 | ~n9853;
  assign n10018 = ~STATE_REG_1__SCAN_IN;
  assign n10011 = ~n10018 & ~n12680;
  assign n9858 = ~n10011 & ~n9855;
  assign n9863 = ~STATE_REG_1__SCAN_IN | ~HOLD;
  assign n10012 = ~STATE_REG_0__SCAN_IN | ~REQUESTPENDING_REG_SCAN_IN;
  assign n9856 = ~n9863 | ~n10012;
  assign n9864 = ~STATE_REG_2__SCAN_IN | ~HOLD;
  assign n9857 = ~n9856 | ~n9864;
  assign U3182 = ~n9858 | ~n9857;
  assign n9860 = ~W_R_N_REG_SCAN_IN | ~n13517;
  assign n9859 = READREQUEST_REG_SCAN_IN | n13517;
  assign U3470 = ~n9860 | ~n9859;
  assign n9862 = ~NA_N | ~n9861;
  assign n9866 = ~n9863 | ~n9862;
  assign n9865 = ~REQUESTPENDING_REG_SCAN_IN | ~n9864;
  assign n9867 = ~n9866 & ~n9865;
  assign n9868 = ~n9867 & ~n13515;
  assign n13514 = ~STATE_REG_2__SCAN_IN & ~STATE_REG_0__SCAN_IN;
  assign n9870 = ~n9868 & ~n13514;
  assign n9869 = ~n10011 | ~n7393;
  assign U3181 = ~n9870 | ~n9869;
  assign n12031 = ~REIP_REG_15__SCAN_IN;
  assign n10001 = ~STATE_REG_2__SCAN_IN | ~n13515;
  assign n9872 = ~n12031 & ~n10001;
  assign n9999 = ~n13515 | ~n7393;
  assign n9871 = ~n12676 & ~n9999;
  assign n9874 = ~n9872 & ~n9871;
  assign n9873 = ~ADDRESS_REG_14__SCAN_IN | ~n13517;
  assign U3198 = ~n9874 | ~n9873;
  assign n9876 = ~n12676 & ~n10001;
  assign n9897 = ~REIP_REG_17__SCAN_IN;
  assign n9875 = ~n9897 & ~n9999;
  assign n9878 = ~n9876 & ~n9875;
  assign n9877 = ~ADDRESS_REG_15__SCAN_IN | ~n13517;
  assign U3199 = ~n9878 | ~n9877;
  assign n9880 = ~n9169 & ~n10001;
  assign n13221 = ~REIP_REG_22__SCAN_IN;
  assign n9879 = ~n13221 & ~n9999;
  assign n9882 = ~n9880 & ~n9879;
  assign n9881 = ~ADDRESS_REG_20__SCAN_IN | ~n13517;
  assign U3204 = ~n9882 | ~n9881;
  assign n9885 = ~n9888 & ~n10001;
  assign n9884 = ~n9883 & ~n9999;
  assign n9887 = ~n9885 & ~n9884;
  assign n9886 = ~ADDRESS_REG_29__SCAN_IN | ~n13517;
  assign U3213 = ~n9887 | ~n9886;
  assign n9890 = ~n13200 & ~n10001;
  assign n9889 = ~n9888 & ~n9999;
  assign n9892 = ~n9890 & ~n9889;
  assign n9891 = ~ADDRESS_REG_28__SCAN_IN | ~n13517;
  assign U3212 = ~n9892 | ~n9891;
  assign n9894 = ~n12630 & ~n10001;
  assign n9893 = ~n12380 & ~n9999;
  assign n9896 = ~n9894 & ~n9893;
  assign n9895 = ~ADDRESS_REG_7__SCAN_IN | ~n13517;
  assign U3191 = ~n9896 | ~n9895;
  assign n9899 = ~n9897 & ~n10001;
  assign n9898 = ~n9918 & ~n9999;
  assign n9901 = ~n9899 & ~n9898;
  assign n9900 = ~ADDRESS_REG_16__SCAN_IN | ~n13517;
  assign U3200 = ~n9901 | ~n9900;
  assign n13035 = ~REIP_REG_26__SCAN_IN;
  assign n9903 = ~n13035 & ~n10001;
  assign n9902 = ~n13126 & ~n9999;
  assign n9905 = ~n9903 & ~n9902;
  assign n9904 = ~ADDRESS_REG_25__SCAN_IN | ~n13517;
  assign U3209 = ~n9905 | ~n9904;
  assign n9907 = ~n12650 & ~n10001;
  assign n9906 = ~n12447 & ~n9999;
  assign n9909 = ~n9907 & ~n9906;
  assign n9908 = ~ADDRESS_REG_4__SCAN_IN | ~n13517;
  assign U3188 = ~n9909 | ~n9908;
  assign n9957 = ~REIP_REG_24__SCAN_IN;
  assign n9911 = ~n9957 & ~n10001;
  assign n13024 = ~REIP_REG_25__SCAN_IN;
  assign n9910 = ~n13024 & ~n9999;
  assign n9913 = ~n9911 & ~n9910;
  assign n9912 = ~ADDRESS_REG_23__SCAN_IN | ~n13517;
  assign U3207 = ~n9913 | ~n9912;
  assign n9915 = ~n13126 & ~n10001;
  assign n13124 = ~REIP_REG_28__SCAN_IN;
  assign n9914 = ~n13124 & ~n9999;
  assign n9917 = ~n9915 & ~n9914;
  assign n9916 = ~ADDRESS_REG_26__SCAN_IN | ~n13517;
  assign U3210 = ~n9917 | ~n9916;
  assign n9920 = ~n9918 & ~n10001;
  assign n12817 = ~REIP_REG_19__SCAN_IN;
  assign n9919 = ~n12817 & ~n9999;
  assign n9922 = ~n9920 & ~n9919;
  assign n9921 = ~ADDRESS_REG_17__SCAN_IN | ~n13517;
  assign U3201 = ~n9922 | ~n9921;
  assign n9967 = ~REIP_REG_11__SCAN_IN;
  assign n9924 = ~n9967 & ~n10001;
  assign n9989 = ~REIP_REG_12__SCAN_IN;
  assign n9923 = ~n9989 & ~n9999;
  assign n9926 = ~n9924 & ~n9923;
  assign n9925 = ~ADDRESS_REG_10__SCAN_IN | ~n13517;
  assign U3194 = ~n9926 | ~n9925;
  assign n10000 = ~REIP_REG_20__SCAN_IN;
  assign n9928 = ~n10000 & ~n10001;
  assign n9927 = ~n9169 & ~n9999;
  assign n9930 = ~n9928 & ~n9927;
  assign n9929 = ~ADDRESS_REG_19__SCAN_IN | ~n13517;
  assign U3203 = ~n9930 | ~n9929;
  assign n9932 = ~n12380 & ~n10001;
  assign n11901 = ~REIP_REG_10__SCAN_IN;
  assign n9931 = ~n11901 & ~n9999;
  assign n9934 = ~n9932 & ~n9931;
  assign n9933 = ~ADDRESS_REG_8__SCAN_IN | ~n13517;
  assign U3192 = ~n9934 | ~n9933;
  assign n9936 = ~n13221 & ~n10001;
  assign n9935 = ~n9956 & ~n9999;
  assign n9938 = ~n9936 & ~n9935;
  assign n9937 = ~ADDRESS_REG_21__SCAN_IN | ~n13517;
  assign U3205 = ~n9938 | ~n9937;
  assign n9940 = ~n12603 & ~n10001;
  assign n9939 = ~n9951 & ~n9999;
  assign n9942 = ~n9940 & ~n9939;
  assign n9941 = ~ADDRESS_REG_12__SCAN_IN | ~n13517;
  assign U3196 = ~n9942 | ~n9941;
  assign n9944 = ~n12447 & ~n10001;
  assign n9943 = ~n12418 & ~n9999;
  assign n9946 = ~n9944 & ~n9943;
  assign n9945 = ~ADDRESS_REG_5__SCAN_IN | ~n13517;
  assign U3189 = ~n9946 | ~n9945;
  assign n9962 = ~REIP_REG_3__SCAN_IN;
  assign n9948 = ~n9962 & ~n10001;
  assign n9947 = ~n9994 & ~n9999;
  assign n9950 = ~n9948 & ~n9947;
  assign n9949 = ~ADDRESS_REG_2__SCAN_IN | ~n13517;
  assign U3186 = ~n9950 | ~n9949;
  assign n9953 = ~n9951 & ~n10001;
  assign n9952 = ~n12031 & ~n9999;
  assign n9955 = ~n9953 & ~n9952;
  assign n9954 = ~ADDRESS_REG_13__SCAN_IN | ~n13517;
  assign U3197 = ~n9955 | ~n9954;
  assign n9959 = ~n9956 & ~n10001;
  assign n9958 = ~n9957 & ~n9999;
  assign n9961 = ~n9959 & ~n9958;
  assign n9960 = ~ADDRESS_REG_22__SCAN_IN | ~n13517;
  assign U3206 = ~n9961 | ~n9960;
  assign n12284 = ~REIP_REG_2__SCAN_IN;
  assign n9964 = ~n12284 & ~n10001;
  assign n9963 = ~n9962 & ~n9999;
  assign n9966 = ~n9964 & ~n9963;
  assign n9965 = ~ADDRESS_REG_1__SCAN_IN | ~n13517;
  assign U3185 = ~n9966 | ~n9965;
  assign n9969 = ~n11901 & ~n10001;
  assign n9968 = ~n9967 & ~n9999;
  assign n9971 = ~n9969 & ~n9968;
  assign n9970 = ~ADDRESS_REG_9__SCAN_IN | ~n13517;
  assign U3193 = ~n9971 | ~n9970;
  assign n9973 = ~n13035 & ~n9999;
  assign n9972 = ~n13024 & ~n10001;
  assign n9975 = ~n9973 & ~n9972;
  assign n9974 = ~ADDRESS_REG_24__SCAN_IN | ~n13517;
  assign U3208 = ~n9975 | ~n9974;
  assign n9977 = ~n12630 & ~n9999;
  assign n9976 = ~n12418 & ~n10001;
  assign n9979 = ~n9977 & ~n9976;
  assign n9978 = ~ADDRESS_REG_6__SCAN_IN | ~n13517;
  assign U3190 = ~n9979 | ~n9978;
  assign n9981 = ~n13200 & ~n9999;
  assign n9980 = ~n13124 & ~n10001;
  assign n9983 = ~n9981 & ~n9980;
  assign n9982 = ~ADDRESS_REG_27__SCAN_IN | ~n13517;
  assign U3211 = ~n9983 | ~n9982;
  assign n9986 = ~n12284 & ~n9999;
  assign n9985 = ~n9984 & ~n10001;
  assign n9988 = ~n9986 & ~n9985;
  assign n9987 = ~ADDRESS_REG_0__SCAN_IN | ~n13517;
  assign U3184 = ~n9988 | ~n9987;
  assign n9991 = ~n12603 & ~n9999;
  assign n9990 = ~n9989 & ~n10001;
  assign n9993 = ~n9991 & ~n9990;
  assign n9992 = ~ADDRESS_REG_11__SCAN_IN | ~n13517;
  assign U3195 = ~n9993 | ~n9992;
  assign n9996 = ~n12650 & ~n9999;
  assign n9995 = ~n9994 & ~n10001;
  assign n9998 = ~n9996 & ~n9995;
  assign n9997 = ~ADDRESS_REG_3__SCAN_IN | ~n13517;
  assign U3187 = ~n9998 | ~n9997;
  assign n10003 = ~n10000 & ~n9999;
  assign n10002 = ~n12817 & ~n10001;
  assign n10005 = ~n10003 & ~n10002;
  assign n10004 = ~ADDRESS_REG_18__SCAN_IN | ~n13517;
  assign U3202 = ~n10005 | ~n10004;
  assign n10006 = ~NA_N & ~n12680;
  assign n10007 = ~n10018 & ~n10006;
  assign n10008 = ~REQUESTPENDING_REG_SCAN_IN & ~n10007;
  assign n10010 = ~STATE_REG_2__SCAN_IN & ~n10008;
  assign n10009 = ~STATE_REG_0__SCAN_IN | ~HOLD;
  assign n10017 = ~n10010 & ~n10009;
  assign n10015 = ~n10011;
  assign n10013 = ~NA_N & ~n10012;
  assign n10014 = ~STATE_REG_2__SCAN_IN & ~n10013;
  assign n10016 = ~n10015 & ~n10014;
  assign n10022 = ~n10017 & ~n10016;
  assign n10020 = ~STATE_REG_0__SCAN_IN & ~n7393;
  assign n10019 = ~NA_N | ~n10018;
  assign n10021 = ~n10020 | ~n10019;
  assign U3183 = ~n10022 | ~n10021;
  assign n10025 = ~n13517 | ~n10023;
  assign U3174 = DATAWIDTH_REG_8__SCAN_IN & n10025;
  assign U3172 = DATAWIDTH_REG_10__SCAN_IN & n10025;
  assign U3151 = DATAWIDTH_REG_31__SCAN_IN & n10025;
  assign U3171 = DATAWIDTH_REG_11__SCAN_IN & n10025;
  assign U3170 = DATAWIDTH_REG_12__SCAN_IN & n10025;
  assign U3175 = DATAWIDTH_REG_7__SCAN_IN & n10025;
  assign U3176 = DATAWIDTH_REG_6__SCAN_IN & n10025;
  assign U3177 = DATAWIDTH_REG_5__SCAN_IN & n10025;
  assign U3178 = DATAWIDTH_REG_4__SCAN_IN & n10025;
  assign U3180 = DATAWIDTH_REG_2__SCAN_IN & n10025;
  assign U3179 = DATAWIDTH_REG_3__SCAN_IN & n10025;
  assign n10024 = ~BS16_N & ~n13514;
  assign n10028 = ~n10024 & ~n10025;
  assign n10026 = ~DATAWIDTH_REG_0__SCAN_IN & ~n10027;
  assign U3451 = ~n10028 & ~n10026;
  assign U3153 = DATAWIDTH_REG_29__SCAN_IN & n10025;
  assign U3152 = DATAWIDTH_REG_30__SCAN_IN & n10025;
  assign U3173 = DATAWIDTH_REG_9__SCAN_IN & n10025;
  assign U3162 = DATAWIDTH_REG_20__SCAN_IN & n10025;
  assign U3161 = DATAWIDTH_REG_21__SCAN_IN & n10025;
  assign U3160 = DATAWIDTH_REG_22__SCAN_IN & n10025;
  assign U3169 = DATAWIDTH_REG_13__SCAN_IN & n10025;
  assign U3168 = DATAWIDTH_REG_14__SCAN_IN & n10025;
  assign U3167 = DATAWIDTH_REG_15__SCAN_IN & n10025;
  assign U3166 = DATAWIDTH_REG_16__SCAN_IN & n10025;
  assign U3165 = DATAWIDTH_REG_17__SCAN_IN & n10025;
  assign U3164 = DATAWIDTH_REG_18__SCAN_IN & n10025;
  assign U3163 = DATAWIDTH_REG_19__SCAN_IN & n10025;
  assign U3158 = DATAWIDTH_REG_24__SCAN_IN & n10025;
  assign U3157 = DATAWIDTH_REG_25__SCAN_IN & n10025;
  assign U3156 = DATAWIDTH_REG_26__SCAN_IN & n10025;
  assign U3159 = DATAWIDTH_REG_23__SCAN_IN & n10025;
  assign U3154 = DATAWIDTH_REG_28__SCAN_IN & n10025;
  assign U3155 = DATAWIDTH_REG_27__SCAN_IN & n10025;
  assign n10031 = ~n10028;
  assign n10029 = ~STATEBS16_REG_SCAN_IN | ~n10025;
  assign U2792 = ~n10031 | ~n10029;
  assign n10030 = ~DATAWIDTH_REG_1__SCAN_IN | ~n10025;
  assign U3452 = ~n10031 | ~n10030;
  assign n11631 = ~n10034;
  assign n10037 = ~n10242 & ~n11631;
  assign n10036 = ~MEMORYFETCH_REG_SCAN_IN | ~n10035;
  assign U2788 = ~n10037 | ~n10036;
  assign n10042 = ~n11631 | ~STATE2_REG_0__SCAN_IN;
  assign n10040 = ~n10039 | ~n10038;
  assign n10041 = ~CODEFETCH_REG_SCAN_IN | ~n10040;
  assign U2790 = ~n10042 | ~n10041;
  assign n10069 = ~n10043 | ~n12691;
  assign n10044 = ~FLUSH_REG_SCAN_IN | ~n10069;
  assign U2793 = ~n13465 | ~n10044;
  assign n10049 = ~n10061 & ~n11631;
  assign n10048 = ~n10049;
  assign n10046 = ~n11647 & ~n11497;
  assign n10047 = ~n10046 | ~n9723;
  assign n10051 = ~n10048 | ~n10047;
  assign n10050 = ~n10049 | ~READREQUEST_REG_SCAN_IN;
  assign U3474 = ~n10051 | ~n10050;
  assign n10053 = ~n10076 | ~n11478;
  assign n10052 = ~n11497 & ~READY_N;
  assign n10054 = ~n10053 | ~n10052;
  assign n10059 = ~n10055 & ~n10054;
  assign n10058 = ~n10057 | ~n10056;
  assign n10062 = ~n10059 & ~n10058;
  assign n10064 = n10061 | n10060;
  assign n10068 = ~n10062 | ~n10064;
  assign n10202 = n10063 & STATE2_REG_2__SCAN_IN;
  assign n10065 = n10202 & n12680;
  assign n10066 = ~n10065 & ~n10064;
  assign n10067 = ~REQUESTPENDING_REG_SCAN_IN | ~n10066;
  assign U3472 = ~n10068 | ~n10067;
  assign n10073 = ~MORE_REG_SCAN_IN | ~n10069;
  assign n10070 = ~n10069;
  assign n10072 = ~n10071 | ~n10070;
  assign U3471 = ~n10073 | ~n10072;
  assign n10078 = ~n10075 & ~n10074;
  assign U2892 = n10206 & DATAO_REG_31__SCAN_IN;
  assign n10082 = ~n10169 | ~EAX_REG_19__SCAN_IN;
  assign n10081 = ~n10202 | ~UWORD_REG_3__SCAN_IN;
  assign n10084 = n10082 & n10081;
  assign U2904 = ~n10084 | ~n10083;
  assign n10086 = ~n10169 | ~EAX_REG_21__SCAN_IN;
  assign n10085 = ~n10202 | ~UWORD_REG_5__SCAN_IN;
  assign n10088 = n10086 & n10085;
  assign U2902 = ~n10088 | ~n10087;
  assign n10090 = ~n10169 | ~EAX_REG_22__SCAN_IN;
  assign n10089 = ~n10202 | ~UWORD_REG_6__SCAN_IN;
  assign n10092 = n10090 & n10089;
  assign U2901 = ~n10092 | ~n10091;
  assign n10094 = ~n10169 | ~EAX_REG_23__SCAN_IN;
  assign n10093 = ~n10202 | ~UWORD_REG_7__SCAN_IN;
  assign n10096 = n10094 & n10093;
  assign U2900 = ~n10096 | ~n10095;
  assign n10098 = ~n10169 | ~EAX_REG_24__SCAN_IN;
  assign n10097 = ~n10202 | ~UWORD_REG_8__SCAN_IN;
  assign n10100 = n10098 & n10097;
  assign U2899 = ~n10100 | ~n10099;
  assign n10102 = ~n10169 | ~EAX_REG_25__SCAN_IN;
  assign n10101 = ~n10202 | ~UWORD_REG_9__SCAN_IN;
  assign n10104 = n10102 & n10101;
  assign U2898 = ~n10104 | ~n10103;
  assign n10106 = ~n10169 | ~EAX_REG_26__SCAN_IN;
  assign n10105 = ~n10202 | ~UWORD_REG_10__SCAN_IN;
  assign n10108 = n10106 & n10105;
  assign U2897 = ~n10108 | ~n10107;
  assign n10110 = ~n10169 | ~EAX_REG_17__SCAN_IN;
  assign n10109 = ~n10202 | ~UWORD_REG_1__SCAN_IN;
  assign n10112 = n10110 & n10109;
  assign U2906 = ~n10112 | ~n10111;
  assign n10114 = ~n10169 | ~EAX_REG_18__SCAN_IN;
  assign n10113 = ~n10202 | ~UWORD_REG_2__SCAN_IN;
  assign n10116 = n10114 & n10113;
  assign U2905 = ~n10116 | ~n10115;
  assign n10118 = ~n10169 | ~EAX_REG_27__SCAN_IN;
  assign n10117 = ~n10202 | ~UWORD_REG_11__SCAN_IN;
  assign n10120 = n10118 & n10117;
  assign U2896 = ~n10120 | ~n10119;
  assign n10122 = ~n10169 | ~EAX_REG_20__SCAN_IN;
  assign n10121 = ~n10202 | ~UWORD_REG_4__SCAN_IN;
  assign n10124 = n10122 & n10121;
  assign U2903 = ~n10124 | ~n10123;
  assign n10126 = ~n10169 | ~EAX_REG_28__SCAN_IN;
  assign n10125 = ~n10202 | ~UWORD_REG_12__SCAN_IN;
  assign n10128 = n10126 & n10125;
  assign U2895 = ~n10128 | ~n10127;
  assign n10130 = ~EAX_REG_7__SCAN_IN | ~n10203;
  assign n10129 = ~n10202 | ~LWORD_REG_7__SCAN_IN;
  assign n10132 = n10130 & n10129;
  assign U2916 = ~n10132 | ~n10131;
  assign n10134 = ~EAX_REG_9__SCAN_IN | ~n10203;
  assign n10133 = ~n10202 | ~LWORD_REG_9__SCAN_IN;
  assign n10136 = n10134 & n10133;
  assign U2914 = ~n10136 | ~n10135;
  assign n10138 = ~EAX_REG_5__SCAN_IN | ~n10203;
  assign n10137 = ~n10202 | ~LWORD_REG_5__SCAN_IN;
  assign n10140 = n10138 & n10137;
  assign U2918 = ~n10140 | ~n10139;
  assign n10142 = ~EAX_REG_15__SCAN_IN | ~n10203;
  assign n10141 = ~n10202 | ~LWORD_REG_15__SCAN_IN;
  assign n10144 = n10142 & n10141;
  assign U2908 = ~n10144 | ~n10143;
  assign n10146 = ~EAX_REG_6__SCAN_IN | ~n10203;
  assign n10145 = ~n10202 | ~LWORD_REG_6__SCAN_IN;
  assign n10148 = n10146 & n10145;
  assign U2917 = ~n10148 | ~n10147;
  assign n10150 = ~EAX_REG_12__SCAN_IN | ~n10203;
  assign n10149 = ~n10202 | ~LWORD_REG_12__SCAN_IN;
  assign n10152 = n10150 & n10149;
  assign U2911 = ~n10152 | ~n10151;
  assign n10154 = ~EAX_REG_13__SCAN_IN | ~n10203;
  assign n10153 = ~n10202 | ~LWORD_REG_13__SCAN_IN;
  assign n10156 = n10154 & n10153;
  assign U2910 = ~n10156 | ~n10155;
  assign n10158 = ~EAX_REG_0__SCAN_IN | ~n10203;
  assign n10157 = ~n10202 | ~LWORD_REG_0__SCAN_IN;
  assign n10160 = n10158 & n10157;
  assign U2923 = ~n10160 | ~n10159;
  assign n10162 = ~n10202 | ~UWORD_REG_13__SCAN_IN;
  assign n10161 = ~n10169 | ~EAX_REG_29__SCAN_IN;
  assign n10164 = n10162 & n10161;
  assign U2894 = ~n10164 | ~n10163;
  assign n10166 = ~n10202 | ~UWORD_REG_0__SCAN_IN;
  assign n10165 = ~n10169 | ~EAX_REG_16__SCAN_IN;
  assign n10168 = n10166 & n10165;
  assign U2907 = ~n10168 | ~n10167;
  assign n10171 = ~n10202 | ~UWORD_REG_14__SCAN_IN;
  assign n10170 = ~n10169 | ~EAX_REG_30__SCAN_IN;
  assign n10173 = n10171 & n10170;
  assign U2893 = ~n10173 | ~n10172;
  assign n10175 = ~n10202 | ~LWORD_REG_3__SCAN_IN;
  assign n10174 = ~EAX_REG_3__SCAN_IN | ~n10203;
  assign n10177 = n10175 & n10174;
  assign U2920 = ~n10177 | ~n10176;
  assign n10179 = ~n10202 | ~LWORD_REG_11__SCAN_IN;
  assign n10178 = ~EAX_REG_11__SCAN_IN | ~n10203;
  assign n10181 = n10179 & n10178;
  assign U2912 = ~n10181 | ~n10180;
  assign n10183 = ~n10202 | ~LWORD_REG_10__SCAN_IN;
  assign n10182 = ~EAX_REG_10__SCAN_IN | ~n10203;
  assign n10185 = n10183 & n10182;
  assign U2913 = ~n10185 | ~n10184;
  assign n10187 = ~n10202 | ~LWORD_REG_1__SCAN_IN;
  assign n10186 = ~EAX_REG_1__SCAN_IN | ~n10203;
  assign n10189 = n10187 & n10186;
  assign U2922 = ~n10189 | ~n10188;
  assign n10191 = ~n10202 | ~LWORD_REG_8__SCAN_IN;
  assign n10190 = ~EAX_REG_8__SCAN_IN | ~n10203;
  assign n10193 = n10191 & n10190;
  assign U2915 = ~n10193 | ~n10192;
  assign n10195 = ~n10202 | ~LWORD_REG_2__SCAN_IN;
  assign n10194 = ~EAX_REG_2__SCAN_IN | ~n10203;
  assign n10197 = n10195 & n10194;
  assign U2921 = ~n10197 | ~n10196;
  assign n10199 = ~n10202 | ~LWORD_REG_14__SCAN_IN;
  assign n10198 = ~EAX_REG_14__SCAN_IN | ~n10203;
  assign n10201 = n10199 & n10198;
  assign U2909 = ~n10201 | ~n10200;
  assign n10205 = ~n10202 | ~LWORD_REG_4__SCAN_IN;
  assign n10204 = ~EAX_REG_4__SCAN_IN | ~n10203;
  assign n10208 = n10205 & n10204;
  assign U2919 = ~n10208 | ~n10207;
  assign n10210 = ~n10209 | ~n13164;
  assign n10221 = ~n10210 | ~PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n10212 = ~n10211 & ~n11497;
  assign n10214 = ~n10213 | ~n10212;
  assign n10219 = ~n10927 & ~n13451;
  assign n11390 = ~REIP_REG_0__SCAN_IN | ~n13491;
  assign n11388 = n10216 ^ n8001;
  assign n10217 = ~n13348 | ~n11388;
  assign n10218 = ~n11390 | ~n10217;
  assign n10220 = ~n10219 & ~n10218;
  assign U2986 = ~n10221 | ~n10220;
  assign n10225 = ~n10223 | ~n10222;
  assign n10226 = ~n10225 ^ n10224;
  assign n10229 = ~n10226 | ~n11578;
  assign n10227 = ~n10226;
  assign n10228 = ~n10227 | ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n11093 = ~n10229 | ~n10228;
  assign n10232 = ~n13465 & ~n11093;
  assign n11094 = ~REIP_REG_1__SCAN_IN | ~n13491;
  assign n10230 = ~PHYADDRPOINTER_REG_1__SCAN_IN | ~n13467;
  assign n10231 = ~n11094 | ~n10230;
  assign n10239 = ~n10232 & ~n10231;
  assign n10237 = ~n13316 & ~PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n10235 = n10234 | n10233;
  assign n10236 = ~n11712 & ~n13451;
  assign n10238 = ~n10237 & ~n10236;
  assign U2985 = ~n10239 | ~n10238;
  assign n10244 = ~n7005 | ~EAX_REG_26__SCAN_IN;
  assign n10243 = ~UWORD_REG_10__SCAN_IN | ~n13567;
  assign n10246 = n10244 & n10243;
  assign n13566 = ~n13567 & ~n10245;
  assign U2934 = ~n10246 | ~n10439;
  assign n10248 = ~n7005 | ~EAX_REG_2__SCAN_IN;
  assign n10247 = ~LWORD_REG_2__SCAN_IN | ~n13567;
  assign n10249 = n10248 & n10247;
  assign U2941 = ~n10249 | ~n10283;
  assign n10251 = ~n7005 | ~EAX_REG_11__SCAN_IN;
  assign n10250 = ~LWORD_REG_11__SCAN_IN | ~n13567;
  assign n10252 = n10251 & n10250;
  assign U2950 = ~n10252 | ~n10273;
  assign n10254 = ~n7005 | ~EAX_REG_24__SCAN_IN;
  assign n10253 = ~UWORD_REG_8__SCAN_IN | ~n13567;
  assign n10255 = n10254 & n10253;
  assign U2932 = ~n10255 | ~n10410;
  assign n10257 = ~n7005 | ~EAX_REG_9__SCAN_IN;
  assign n10256 = ~LWORD_REG_9__SCAN_IN | ~n13567;
  assign n10258 = n10257 & n10256;
  assign U2948 = ~n10258 | ~n10293;
  assign n10260 = ~n7005 | ~EAX_REG_22__SCAN_IN;
  assign n10259 = ~UWORD_REG_6__SCAN_IN | ~n13567;
  assign n10261 = n10260 & n10259;
  assign U2930 = ~n10261 | ~n10426;
  assign n10263 = ~n7005 | ~EAX_REG_20__SCAN_IN;
  assign n10262 = ~UWORD_REG_4__SCAN_IN | ~n13567;
  assign n10264 = n10263 & n10262;
  assign U2928 = ~n10264 | ~n10418;
  assign n10266 = ~n7005 | ~EAX_REG_16__SCAN_IN;
  assign n10265 = ~UWORD_REG_0__SCAN_IN | ~n13567;
  assign n10267 = n10266 & n10265;
  assign U2924 = ~n10267 | ~n10430;
  assign n10269 = ~UWORD_REG_5__SCAN_IN | ~n13567;
  assign n10268 = ~n7005 | ~EAX_REG_21__SCAN_IN;
  assign n10270 = n10269 & n10268;
  assign U2929 = ~n10270 | ~n10435;
  assign n10272 = ~UWORD_REG_11__SCAN_IN | ~n13567;
  assign n10271 = ~n7005 | ~EAX_REG_27__SCAN_IN;
  assign n10274 = n10272 & n10271;
  assign U2935 = ~n10274 | ~n10273;
  assign n10276 = ~UWORD_REG_7__SCAN_IN | ~n13567;
  assign n10275 = ~n7005 | ~EAX_REG_23__SCAN_IN;
  assign n10277 = n10276 & n10275;
  assign U2931 = ~n10277 | ~n10414;
  assign n10279 = ~UWORD_REG_12__SCAN_IN | ~n13567;
  assign n10278 = ~n7005 | ~EAX_REG_28__SCAN_IN;
  assign n10280 = n10279 & n10278;
  assign U2936 = ~n10280 | ~n10406;
  assign n10282 = ~UWORD_REG_2__SCAN_IN | ~n13567;
  assign n10281 = ~n7005 | ~EAX_REG_18__SCAN_IN;
  assign n10284 = n10282 & n10281;
  assign U2926 = ~n10284 | ~n10283;
  assign n10286 = ~UWORD_REG_13__SCAN_IN | ~n13567;
  assign n10285 = ~n7005 | ~EAX_REG_29__SCAN_IN;
  assign n10287 = n10286 & n10285;
  assign U2937 = ~n10287 | ~n10422;
  assign n10289 = ~UWORD_REG_1__SCAN_IN | ~n13567;
  assign n10288 = ~n7005 | ~EAX_REG_17__SCAN_IN;
  assign n10290 = n10289 & n10288;
  assign U2925 = ~n10290 | ~n10402;
  assign n10292 = ~UWORD_REG_9__SCAN_IN | ~n13567;
  assign n10291 = ~n7005 | ~EAX_REG_25__SCAN_IN;
  assign n10294 = n10292 & n10291;
  assign U2933 = ~n10294 | ~n10293;
  assign n10296 = ~n12799 & ~n10927;
  assign n10295 = ~n8119 & ~n13391;
  assign n10299 = ~n10296 & ~n10295;
  assign n12099 = ~n13178 & ~n10297;
  assign n10298 = ~n12099 | ~DATAI_0_;
  assign U2891 = ~n10299 | ~n10298;
  assign n10399 = ~EAX_REG_1__SCAN_IN;
  assign n10301 = ~n10399 & ~n13391;
  assign n10300 = ~n12799 & ~n11712;
  assign n10303 = ~n10301 & ~n10300;
  assign n10302 = ~n12099 | ~DATAI_1_;
  assign U2890 = ~n10303 | ~n10302;
  assign n10454 = ~EAX_REG_3__SCAN_IN;
  assign n10309 = ~n10454 & ~n13391;
  assign n10307 = ~n10313;
  assign n10306 = ~n10305 | ~n10304;
  assign n10308 = ~n12799 & ~n13557;
  assign n10311 = ~n10309 & ~n10308;
  assign n10310 = ~n12099 | ~DATAI_3_;
  assign U2888 = ~n10311 | ~n10310;
  assign n10315 = ~n8148 & ~n13391;
  assign n10859 = ~n11649;
  assign n10314 = ~n12799 & ~n10859;
  assign n10317 = ~n10315 & ~n10314;
  assign n10316 = ~n12099 | ~DATAI_4_;
  assign U2887 = ~n10317 | ~n10316;
  assign n11567 = ~REIP_REG_2__SCAN_IN | ~n13491;
  assign n10318 = ~PHYADDRPOINTER_REG_2__SCAN_IN | ~n13467;
  assign n10326 = ~n11567 | ~n10318;
  assign n10324 = ~n12297 | ~n13463;
  assign n10323 = ~n12292 | ~n13472;
  assign n11573 = n10328 ^ n10327;
  assign n10329 = ~n13348 | ~n11573;
  assign U2984 = ~n10330 | ~n10329;
  assign n12507 = ~n10485 | ~STATE2_REG_0__SCAN_IN;
  assign n10333 = ~n12507 & ~n7597;
  assign n10332 = ~n12324 & ~STATE2_REG_0__SCAN_IN;
  assign n10334 = ~n10333 & ~n10332;
  assign n10336 = ~n10341 | ~n10372;
  assign n10337 = ~n10395 | ~n10336;
  assign n10349 = ~n10337 | ~INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n10346 = ~n10338 | ~n12681;
  assign n10370 = INSTADDRPOINTER_REG_31__SCAN_IN ^ INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n10339 = ~n10370;
  assign n10371 = ~STATE2_REG_1__SCAN_IN | ~INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n10344 = ~n10339 & ~n10371;
  assign n10342 = ~n10340 | ~n10372;
  assign n10343 = ~n10342 & ~n10341;
  assign n10345 = ~n10344 & ~n10343;
  assign n10347 = ~n10346 | ~n10345;
  assign n10348 = ~n10347 | ~n10395;
  assign U3459 = ~n10349 | ~n10348;
  assign n10355 = ~n10432 & ~n13391;
  assign n10353 = ~n10461;
  assign n10354 = ~n12799 & ~n13551;
  assign n10357 = ~n10355 & ~n10354;
  assign n10356 = ~n12099 | ~DATAI_5_;
  assign U2886 = ~n10357 | ~n10356;
  assign n10359 = ~EAX_REG_2__SCAN_IN | ~n13178;
  assign n10358 = ~n12099 | ~DATAI_2_;
  assign n10361 = n10359 & n10358;
  assign U2889 = ~n10361 | ~n10360;
  assign n10365 = ~n10362 | ~n12681;
  assign n10364 = ~n10363 | ~n10372;
  assign n10366 = ~n10365 | ~n10364;
  assign n10368 = ~n10395 | ~n10366;
  assign n10367 = ~n10396 | ~INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign U3456 = ~n10368 | ~n10367;
  assign n10379 = ~n10369 | ~n12681;
  assign n10377 = ~n10371 & ~n10370;
  assign n10375 = ~n10373 | ~n10372;
  assign n10376 = ~n10375 & ~n10374;
  assign n10378 = ~n10377 & ~n10376;
  assign n10380 = ~n10379 | ~n10378;
  assign n10382 = ~n10395 | ~n10380;
  assign n10381 = ~n10396 | ~INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign U3460 = ~n10382 | ~n10381;
  assign n10387 = ~n10383 | ~n12681;
  assign n10385 = ~n11813 & ~INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n10384 = ~n10488 & ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n10386 = ~n10385 & ~n10384;
  assign n10388 = ~n10387 | ~n10386;
  assign n10390 = ~n10395 | ~n10388;
  assign n10389 = ~n10396 | ~INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign U3461 = ~n10390 | ~n10389;
  assign n10393 = ~n11638;
  assign n10392 = ~n10391 | ~n12681;
  assign n10394 = ~n10393 & ~n10392;
  assign n10398 = ~n10395 | ~n10394;
  assign n10397 = ~n10396 | ~INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign U3455 = ~n10398 | ~n10397;
  assign n10400 = LWORD_REG_1__SCAN_IN & n13567;
  assign U2940 = ~n10403 | ~n10402;
  assign n10404 = LWORD_REG_12__SCAN_IN & n13567;
  assign U2951 = ~n10407 | ~n10406;
  assign n10408 = LWORD_REG_8__SCAN_IN & n13567;
  assign U2947 = ~n10411 | ~n10410;
  assign n10412 = LWORD_REG_7__SCAN_IN & n13567;
  assign U2946 = ~n10415 | ~n10414;
  assign n10416 = LWORD_REG_4__SCAN_IN & n13567;
  assign U2943 = ~n10419 | ~n10418;
  assign n11753 = ~EAX_REG_13__SCAN_IN;
  assign n10420 = LWORD_REG_13__SCAN_IN & n13567;
  assign U2952 = ~n10423 | ~n10422;
  assign n10459 = ~EAX_REG_6__SCAN_IN;
  assign n10424 = LWORD_REG_6__SCAN_IN & n13567;
  assign U2945 = ~n10427 | ~n10426;
  assign n10428 = LWORD_REG_0__SCAN_IN & n13567;
  assign U2939 = ~n10431 | ~n10430;
  assign n10433 = LWORD_REG_5__SCAN_IN & n13567;
  assign U2944 = ~n10436 | ~n10435;
  assign n10437 = LWORD_REG_10__SCAN_IN & n13567;
  assign U2949 = ~n10440 | ~n10439;
  assign n10443 = ~UWORD_REG_14__SCAN_IN | ~n13567;
  assign U2938 = ~n10444 | ~n10443;
  assign n10445 = ~DATAI_3_;
  assign n10448 = ~UWORD_REG_3__SCAN_IN | ~n13567;
  assign U2927 = ~n10449 | ~n10448;
  assign n10452 = ~LWORD_REG_14__SCAN_IN | ~n13567;
  assign U2953 = ~n10453 | ~n10452;
  assign n10457 = ~LWORD_REG_3__SCAN_IN | ~n13567;
  assign U2942 = ~n10458 | ~n10457;
  assign n10464 = ~n10459 & ~n13391;
  assign n10462 = n10461 | n10460;
  assign n10463 = ~n12799 & ~n13545;
  assign n10466 = ~n10464 & ~n10463;
  assign n10465 = ~n12099 | ~DATAI_6_;
  assign U2885 = ~n10466 | ~n10465;
  assign n12286 = n10468 ^ n10467;
  assign n10469 = ~EBX_REG_2__SCAN_IN | ~n13560;
  assign n10472 = n10470 & n10469;
  assign U2857 = ~n10472 | ~n10471;
  assign n10482 = ~n12575 & ~n13316;
  assign n10478 = ~n13557 & ~n13451;
  assign n10475 = n10474 | n10473;
  assign n11333 = ~n10476 | ~n10475;
  assign n10477 = ~n13465 & ~n11333;
  assign n10480 = ~n10478 & ~n10477;
  assign n10479 = ~n13467 | ~PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n10483 = ~n10482 & ~n10481;
  assign n11321 = ~n13491 | ~REIP_REG_3__SCAN_IN;
  assign U2983 = ~n10483 | ~n11321;
  assign n11699 = ~n10496 | ~n10674;
  assign n10503 = ~n11699 & ~n12536;
  assign n10487 = ~n10485;
  assign n10491 = ~n10489 | ~n10488;
  assign n10543 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n12316 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n10543;
  assign n11828 = ~n11949;
  assign n10542 = n12308 | n11828;
  assign n10494 = ~n12316 & ~n11497;
  assign n10498 = ~n12543 & ~n11253;
  assign n12537 = ~n10496 | ~n10886;
  assign n10497 = ~n12537 & ~n12544;
  assign n10501 = ~n10498 & ~n10497;
  assign n10747 = ~n11627 & ~n12324;
  assign n10500 = ~n12538 | ~n11247;
  assign n10502 = ~n10501 | ~n10500;
  assign n10512 = ~n10503 & ~n10502;
  assign n10505 = ~n10504;
  assign n10507 = ~STATE2_REG_3__SCAN_IN | ~n11488;
  assign n10509 = ~n12316 | ~n11480;
  assign n10511 = ~INSTQUEUE_REG_3__5__SCAN_IN | ~n11248;
  assign U3049 = ~n10512 | ~n10511;
  assign n10519 = ~n12537 & ~n12333;
  assign n10514 = ~n12334 & ~n11253;
  assign n10513 = ~n11699 & ~n12335;
  assign n10517 = ~n10514 & ~n10513;
  assign n10516 = ~n12338 | ~n11247;
  assign n10518 = ~n10517 | ~n10516;
  assign n10521 = ~n10519 & ~n10518;
  assign n10520 = ~INSTQUEUE_REG_3__1__SCAN_IN | ~n11248;
  assign U3045 = ~n10521 | ~n10520;
  assign n11872 = ~n10526 | ~n10886;
  assign n10532 = ~n11872 & ~n12333;
  assign n10584 = ~n12145 & ~n10637;
  assign n11730 = ~n10584 | ~n10638;
  assign n12287 = ~n10616;
  assign n10522 = ~n11743 & ~n11828;
  assign n10524 = ~n11730 & ~n11497;
  assign n10528 = ~n12334 & ~n11290;
  assign n12092 = ~n10526 | ~n10674;
  assign n10527 = ~n12092 & ~n12335;
  assign n10530 = ~n10528 & ~n10527;
  assign n10529 = ~n12338 | ~n11284;
  assign n10531 = ~n10530 | ~n10529;
  assign n10540 = ~n10532 & ~n10531;
  assign n10537 = ~n11730 | ~n11480;
  assign n10539 = ~INSTQUEUE_REG_13__1__SCAN_IN | ~n11285;
  assign U3125 = ~n10540 | ~n10539;
  assign n12561 = ~n10548 | ~n10674;
  assign n10554 = ~n12561 & ~n12335;
  assign n11979 = ~n10543 | ~n10638;
  assign n10546 = ~n11979 & ~n11497;
  assign n10550 = ~n12334 & ~n11264;
  assign n10549 = ~n12128 & ~n12333;
  assign n10552 = ~n10550 & ~n10549;
  assign n10551 = ~n12338 | ~n11258;
  assign n10553 = ~n10552 | ~n10551;
  assign n10562 = ~n10554 & ~n10553;
  assign n10556 = ~n10555;
  assign n10559 = ~n11979 | ~n11480;
  assign n10561 = ~INSTQUEUE_REG_1__1__SCAN_IN | ~n11259;
  assign U3029 = ~n10562 | ~n10561;
  assign n10564 = ~n11645 | ~n13472;
  assign n10563 = ~PHYADDRPOINTER_REG_4__SCAN_IN | ~n13467;
  assign n11424 = ~REIP_REG_4__SCAN_IN | ~n13491;
  assign n11429 = n10566 ^ n10565;
  assign n10567 = ~n13348 | ~n11429;
  assign n10568 = ~n11424 | ~n10567;
  assign n10570 = ~n11649 | ~n13463;
  assign U2982 = ~n10571 | ~n10570;
  assign n10578 = ~n12128 & ~n12301;
  assign n10573 = ~n12312 & ~n11264;
  assign n10572 = ~n12561 & ~n12313;
  assign n10576 = ~n10573 & ~n10572;
  assign n10575 = ~n12317 | ~n11258;
  assign n10577 = ~n10576 | ~n10575;
  assign n10580 = ~n10578 & ~n10577;
  assign n10579 = ~INSTQUEUE_REG_1__0__SCAN_IN | ~n11259;
  assign U3028 = ~n10580 | ~n10579;
  assign n12126 = ~n10590 | ~n10674;
  assign n10596 = ~n12126 & ~n12313;
  assign n12050 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n10584;
  assign n10587 = ~n12063 & ~n11828;
  assign n10589 = ~n10598 & ~n10597;
  assign n10588 = ~n12050 & ~n11497;
  assign n10592 = ~n12312 & ~n11311;
  assign n12239 = ~n10590 | ~n10886;
  assign n10591 = ~n12239 & ~n12301;
  assign n10594 = ~n10592 & ~n10591;
  assign n10593 = ~n12317 | ~n10585;
  assign n10595 = ~n10594 | ~n10593;
  assign n10604 = ~n10596 & ~n10595;
  assign n10599 = ~n10597;
  assign n10601 = ~n12050 | ~n11480;
  assign n10603 = ~INSTQUEUE_REG_15__0__SCAN_IN | ~n11306;
  assign U3140 = ~n10604 | ~n10603;
  assign n10610 = ~n12239 & ~n12333;
  assign n10606 = ~n12334 & ~n11311;
  assign n10605 = ~n12126 & ~n12335;
  assign n10608 = ~n10606 & ~n10605;
  assign n10607 = ~n12338 | ~n10585;
  assign n10609 = ~n10608 | ~n10607;
  assign n10612 = ~n10610 & ~n10609;
  assign n10611 = ~INSTQUEUE_REG_15__1__SCAN_IN | ~n11306;
  assign U3141 = ~n10612 | ~n10611;
  assign n10627 = ~n11874 & ~n12335;
  assign n10675 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n10637;
  assign n10892 = n10638 | n10675;
  assign n10618 = ~n10615;
  assign n10620 = n10887 & n10628;
  assign n10619 = ~n10892 & ~n11497;
  assign n10623 = ~n12334 & ~n11300;
  assign n11301 = n10621 | n10674;
  assign n10622 = ~n11301 & ~n12333;
  assign n10625 = ~n10623 & ~n10622;
  assign n10624 = ~n12338 | ~n10615;
  assign n10626 = ~n10625 | ~n10624;
  assign n10634 = ~n10627 & ~n10626;
  assign n10631 = ~n10892 | ~n11480;
  assign n10633 = ~INSTQUEUE_REG_11__1__SCAN_IN | ~n11295;
  assign U3109 = ~n10634 | ~n10633;
  assign n10636 = ~n10635;
  assign n12183 = ~n10642 | ~n10674;
  assign n10648 = ~n12183 & ~n12335;
  assign n10784 = ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~n10637;
  assign n11451 = ~n10784 | ~n10638;
  assign n11457 = n10781 | n7936;
  assign n10639 = ~n11457 & ~n11828;
  assign n10641 = ~n10651 & ~n10649;
  assign n10640 = ~n11451 & ~n11497;
  assign n10644 = ~n12334 & ~n11275;
  assign n10643 = ~n11707 & ~n12333;
  assign n10646 = ~n10644 & ~n10643;
  assign n10645 = ~n12338 | ~n11269;
  assign n10647 = ~n10646 | ~n10645;
  assign n10656 = ~n10648 & ~n10647;
  assign n10650 = ~n10649;
  assign n10653 = ~n11451 | ~n11480;
  assign n10655 = ~INSTQUEUE_REG_5__1__SCAN_IN | ~n11270;
  assign U3061 = ~n10656 | ~n10655;
  assign n10662 = ~n12183 & ~n12313;
  assign n10658 = ~n12312 & ~n11275;
  assign n10657 = ~n11707 & ~n12301;
  assign n10660 = ~n10658 & ~n10657;
  assign n10659 = ~n12317 | ~n11269;
  assign n10661 = ~n10660 | ~n10659;
  assign n10664 = ~n10662 & ~n10661;
  assign n10663 = ~INSTQUEUE_REG_5__0__SCAN_IN | ~n11270;
  assign U3060 = ~n10664 | ~n10663;
  assign n10670 = ~n8177 & ~n13391;
  assign n10669 = ~n12799 & ~n13539;
  assign n10671 = ~n12099 | ~DATAI_7_;
  assign U2884 = ~n10672 | ~n10671;
  assign n10688 = ~n11614 & ~n12544;
  assign n11489 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n10675;
  assign n10680 = ~STATE2_REG_2__SCAN_IN | ~n11489;
  assign n10684 = ~INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n11489;
  assign n10678 = ~n10677 | ~n12307;
  assign n10683 = ~n12543 & ~n11382;
  assign n10682 = ~n11383 & ~n12536;
  assign n10686 = ~n10683 & ~n10682;
  assign n10685 = ~n11376 | ~n12538;
  assign n10687 = ~n10686 | ~n10685;
  assign n10696 = ~n10688 & ~n10687;
  assign n10689 = ~n12305 & ~n11489;
  assign n10691 = ~n10690;
  assign n10695 = ~INSTQUEUE_REG_9__5__SCAN_IN | ~n11377;
  assign U3097 = ~n10696 | ~n10695;
  assign n10702 = ~n11614 & ~n12301;
  assign n10698 = ~n12312 & ~n11382;
  assign n10697 = ~n11383 & ~n12313;
  assign n10700 = ~n10698 & ~n10697;
  assign n10699 = ~n11376 | ~n12317;
  assign n10701 = ~n10700 | ~n10699;
  assign n10704 = ~n10702 & ~n10701;
  assign n10703 = ~INSTQUEUE_REG_9__0__SCAN_IN | ~n11377;
  assign U3092 = ~n10704 | ~n10703;
  assign n10710 = ~n11614 & ~n12333;
  assign n10706 = ~n12334 & ~n11382;
  assign n10705 = ~n11383 & ~n12335;
  assign n10708 = ~n10706 & ~n10705;
  assign n10707 = ~n11376 | ~n12338;
  assign n10709 = ~n10708 | ~n10707;
  assign n10712 = ~n10710 & ~n10709;
  assign n10711 = ~INSTQUEUE_REG_9__1__SCAN_IN | ~n11377;
  assign U3093 = ~n10712 | ~n10711;
  assign n10716 = ~n11872 & ~n12544;
  assign n10714 = ~n12538 | ~n11284;
  assign n10713 = ~INSTQUEUE_REG_13__5__SCAN_IN | ~n11285;
  assign n10715 = ~n10714 | ~n10713;
  assign n10720 = ~n10716 & ~n10715;
  assign n10718 = ~n12543 & ~n11290;
  assign n10717 = ~n12092 & ~n12536;
  assign n10719 = ~n10718 & ~n10717;
  assign U3129 = ~n10720 | ~n10719;
  assign n10724 = ~n11872 & ~n12301;
  assign n10722 = ~n12317 | ~n11284;
  assign n10721 = ~INSTQUEUE_REG_13__0__SCAN_IN | ~n11285;
  assign n10723 = ~n10722 | ~n10721;
  assign n10728 = ~n10724 & ~n10723;
  assign n10726 = ~n12312 & ~n11290;
  assign n10725 = ~n12092 & ~n12313;
  assign n10727 = ~n10726 & ~n10725;
  assign U3124 = ~n10728 | ~n10727;
  assign n10732 = ~n12561 & ~n12536;
  assign n10730 = ~n12538 | ~n11258;
  assign n10729 = ~INSTQUEUE_REG_1__5__SCAN_IN | ~n11259;
  assign n10731 = ~n10730 | ~n10729;
  assign n10736 = ~n10732 & ~n10731;
  assign n10734 = ~n12543 & ~n11264;
  assign n10733 = ~n12128 & ~n12544;
  assign n10735 = ~n10734 & ~n10733;
  assign U3033 = ~n10736 | ~n10735;
  assign n10740 = ~n12239 & ~n12544;
  assign n10738 = ~n12538 | ~n10585;
  assign n10737 = ~INSTQUEUE_REG_15__5__SCAN_IN | ~n11306;
  assign n10739 = ~n10738 | ~n10737;
  assign n10744 = ~n10740 & ~n10739;
  assign n10742 = ~n12543 & ~n11311;
  assign n10741 = ~n12126 & ~n12536;
  assign n10743 = ~n10742 & ~n10741;
  assign U3145 = ~n10744 | ~n10743;
  assign n10752 = ~n11874 & ~n12345;
  assign n10746 = ~n12346 & ~n11300;
  assign n10745 = ~n11301 & ~n12347;
  assign n10750 = ~n10746 & ~n10745;
  assign n12350 = ~n10748 & ~n11155;
  assign n10749 = ~n12350 | ~n10615;
  assign n10751 = ~n10750 | ~n10749;
  assign n10754 = ~n10752 & ~n10751;
  assign n10753 = ~INSTQUEUE_REG_11__3__SCAN_IN | ~n11295;
  assign U3111 = ~n10754 | ~n10753;
  assign n10760 = ~n12239 & ~n12347;
  assign n10756 = ~n12346 & ~n11311;
  assign n10755 = ~n12126 & ~n12345;
  assign n10758 = ~n10756 & ~n10755;
  assign n10757 = ~n12350 | ~n10585;
  assign n10759 = ~n10758 | ~n10757;
  assign n10762 = ~n10760 & ~n10759;
  assign n10761 = ~INSTQUEUE_REG_15__3__SCAN_IN | ~n11306;
  assign U3143 = ~n10762 | ~n10761;
  assign n10766 = ~n11699 & ~n12313;
  assign n10764 = ~n12317 | ~n11247;
  assign n10763 = ~INSTQUEUE_REG_3__0__SCAN_IN | ~n11248;
  assign n10765 = ~n10764 | ~n10763;
  assign n10770 = ~n10766 & ~n10765;
  assign n10768 = ~n12312 & ~n11253;
  assign n10767 = ~n12537 & ~n12301;
  assign n10769 = ~n10768 & ~n10767;
  assign U3044 = ~n10770 | ~n10769;
  assign n10776 = ~n12128 & ~n12347;
  assign n10772 = ~n12346 & ~n11264;
  assign n10771 = ~n12561 & ~n12345;
  assign n10774 = ~n10772 & ~n10771;
  assign n10773 = ~n12350 | ~n11258;
  assign n10775 = ~n10774 | ~n10773;
  assign n10778 = ~n10776 & ~n10775;
  assign n10777 = ~INSTQUEUE_REG_1__3__SCAN_IN | ~n11259;
  assign U3031 = ~n10778 | ~n10777;
  assign n10793 = ~n11606 & ~n12335;
  assign n10782 = ~n12154 & ~n11828;
  assign n12139 = ~INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n10784;
  assign n10785 = ~n12139 & ~n11497;
  assign n10789 = ~n12334 & ~n11363;
  assign n12267 = ~n10787 | ~n10886;
  assign n10788 = ~n12267 & ~n12333;
  assign n10791 = ~n10789 & ~n10788;
  assign n10790 = ~n11357 | ~n12338;
  assign n10792 = ~n10791 | ~n10790;
  assign n10802 = ~n10793 & ~n10792;
  assign n10795 = ~n10794;
  assign n10799 = ~n12139 | ~n11480;
  assign n10801 = ~INSTQUEUE_REG_7__1__SCAN_IN | ~n11358;
  assign U3077 = ~n10802 | ~n10801;
  assign n10808 = ~n12267 & ~n12301;
  assign n10804 = ~n12312 & ~n11363;
  assign n10803 = ~n11606 & ~n12313;
  assign n10806 = ~n10804 & ~n10803;
  assign n10805 = ~n11357 | ~n12317;
  assign n10807 = ~n10806 | ~n10805;
  assign n10810 = ~n10808 & ~n10807;
  assign n10809 = ~INSTQUEUE_REG_7__0__SCAN_IN | ~n11358;
  assign U3076 = ~n10810 | ~n10809;
  assign n10814 = ~n12183 & ~n12536;
  assign n10812 = ~n12538 | ~n11269;
  assign n10811 = ~INSTQUEUE_REG_5__5__SCAN_IN | ~n11270;
  assign n10813 = ~n10812 | ~n10811;
  assign n10818 = ~n10814 & ~n10813;
  assign n10816 = ~n12543 & ~n11275;
  assign n10815 = ~n11707 & ~n12544;
  assign n10817 = ~n10816 & ~n10815;
  assign U3065 = ~n10818 | ~n10817;
  assign n10820 = ~EAX_REG_9__SCAN_IN | ~n13178;
  assign n10819 = ~n12099 | ~DATAI_9_;
  assign n10823 = n10820 & n10819;
  assign U2882 = ~n10823 | ~n10822;
  assign n10829 = ~n8185 & ~n13391;
  assign n10827 = n10825 | n10824;
  assign n10830 = ~n12099 | ~DATAI_8_;
  assign U2883 = ~n10831 | ~n10830;
  assign n10837 = ~n11606 & ~n12345;
  assign n10833 = ~n12346 & ~n11363;
  assign n10832 = ~n12267 & ~n12347;
  assign n10835 = ~n10833 & ~n10832;
  assign n10834 = ~n11357 | ~n12350;
  assign n10836 = ~n10835 | ~n10834;
  assign n10839 = ~n10837 & ~n10836;
  assign n10838 = ~INSTQUEUE_REG_7__3__SCAN_IN | ~n11358;
  assign U3079 = ~n10839 | ~n10838;
  assign n10843 = ~n11874 & ~n12536;
  assign n10841 = ~n12538 | ~n10615;
  assign n10840 = ~INSTQUEUE_REG_11__5__SCAN_IN | ~n11295;
  assign n10842 = ~n10841 | ~n10840;
  assign n10847 = ~n10843 & ~n10842;
  assign n10845 = ~n12543 & ~n11300;
  assign n10844 = ~n11301 & ~n12544;
  assign n10846 = ~n10845 & ~n10844;
  assign U3113 = ~n10847 | ~n10846;
  assign n10851 = ~n11874 & ~n12313;
  assign n10849 = ~n12317 | ~n10615;
  assign n10848 = ~INSTQUEUE_REG_11__0__SCAN_IN | ~n11295;
  assign n10850 = ~n10849 | ~n10848;
  assign n10855 = ~n10851 & ~n10850;
  assign n10853 = ~n12312 & ~n11300;
  assign n10852 = ~n11301 & ~n12301;
  assign n10854 = ~n10853 & ~n10852;
  assign U3108 = ~n10855 | ~n10854;
  assign n10858 = n10857 | n10856;
  assign n11629 = ~n10858 | ~n11402;
  assign n10861 = ~n13528 & ~n11629;
  assign n10860 = ~n8806 & ~n10859;
  assign n10863 = ~n10861 & ~n10860;
  assign n10862 = ~EBX_REG_4__SCAN_IN | ~n13560;
  assign U2855 = ~n10863 | ~n10862;
  assign n12381 = n10865 ^ n10864;
  assign n10866 = ~EBX_REG_9__SCAN_IN | ~n13560;
  assign n10869 = n10867 & n10866;
  assign U2850 = ~n10869 | ~n10868;
  assign n10875 = ~n11614 & ~n12347;
  assign n10871 = ~n12346 & ~n11382;
  assign n10870 = ~n11383 & ~n12345;
  assign n10873 = ~n10871 & ~n10870;
  assign n10872 = ~n11376 | ~n12350;
  assign n10874 = ~n10873 | ~n10872;
  assign n10877 = ~n10875 & ~n10874;
  assign n10876 = ~INSTQUEUE_REG_9__3__SCAN_IN | ~n11377;
  assign U3095 = ~n10877 | ~n10876;
  assign n10881 = ~n11606 & ~n12536;
  assign n10879 = ~n11357 | ~n12538;
  assign n10878 = ~INSTQUEUE_REG_7__5__SCAN_IN | ~n11358;
  assign n10880 = ~n10879 | ~n10878;
  assign n10885 = ~n10881 & ~n10880;
  assign n10883 = ~n12543 & ~n11363;
  assign n10882 = ~n12267 & ~n12544;
  assign n10884 = ~n10883 & ~n10882;
  assign U3081 = ~n10885 | ~n10884;
  assign n10897 = ~n11301 & ~n12313;
  assign n12146 = ~n11441;
  assign n12065 = ~n12146 | ~INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n10888 = ~n12065 & ~n12302;
  assign n10891 = ~n12312 & ~n11171;
  assign n10890 = ~n11383 & ~n12301;
  assign n10895 = ~n10891 & ~n10890;
  assign n10894 = ~n12317 | ~n10893;
  assign n10896 = ~n10895 | ~n10894;
  assign n10910 = ~n10897 & ~n10896;
  assign n10899 = ~n10898;
  assign n12156 = ~n10899 | ~STATE2_REG_2__SCAN_IN;
  assign n10900 = ~n12156;
  assign n12056 = n12065 & STATE2_REG_2__SCAN_IN;
  assign n11851 = ~n11445;
  assign n10905 = ~n12324 & ~n10893;
  assign n10907 = n10906 | n10905;
  assign n10909 = ~INSTQUEUE_REG_10__0__SCAN_IN | ~n11178;
  assign U3100 = ~n10910 | ~n10909;
  assign n10916 = ~n11301 & ~n12345;
  assign n10912 = ~n12346 & ~n11171;
  assign n10911 = ~n11383 & ~n12347;
  assign n10914 = ~n10912 & ~n10911;
  assign n10913 = ~n12350 | ~n10893;
  assign n10915 = ~n10914 | ~n10913;
  assign n10918 = ~n10916 & ~n10915;
  assign n10917 = ~INSTQUEUE_REG_10__3__SCAN_IN | ~n11178;
  assign U3103 = ~n10918 | ~n10917;
  assign n10924 = ~n11301 & ~n12335;
  assign n10920 = ~n12334 & ~n11171;
  assign n10919 = ~n11383 & ~n12333;
  assign n10922 = ~n10920 & ~n10919;
  assign n10921 = ~n12338 | ~n10893;
  assign n10923 = ~n10922 | ~n10921;
  assign n10926 = ~n10924 & ~n10923;
  assign n10925 = ~INSTQUEUE_REG_10__1__SCAN_IN | ~n11178;
  assign U3101 = ~n10926 | ~n10925;
  assign n10931 = ~n8806 & ~n10927;
  assign n10929 = ~EBX_REG_0__SCAN_IN;
  assign n10930 = ~n10929 & ~n10928;
  assign n10936 = ~n10931 & ~n10930;
  assign n10933 = ~n10932 & ~INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n11954 = ~n10934 & ~n10933;
  assign U2859 = ~n10936 | ~n10935;
  assign n11713 = n10938 ^ n10937;
  assign n10940 = ~n13528 & ~n11713;
  assign n10939 = ~n8806 & ~n11712;
  assign n10942 = ~n10940 & ~n10939;
  assign n10941 = ~EBX_REG_1__SCAN_IN | ~n13560;
  assign U2858 = ~n10942 | ~n10941;
  assign n10946 = ~n12183 & ~n12345;
  assign n10944 = ~n12350 | ~n11269;
  assign n10943 = ~INSTQUEUE_REG_5__3__SCAN_IN | ~n11270;
  assign n10945 = ~n10944 | ~n10943;
  assign n10950 = ~n10946 & ~n10945;
  assign n10948 = ~n12346 & ~n11275;
  assign n10947 = ~n11707 & ~n12347;
  assign n10949 = ~n10948 & ~n10947;
  assign U3063 = ~n10950 | ~n10949;
  assign n10954 = ~n11872 & ~n12347;
  assign n10952 = ~n12350 | ~n11284;
  assign n10951 = ~INSTQUEUE_REG_13__3__SCAN_IN | ~n11285;
  assign n10953 = ~n10952 | ~n10951;
  assign n10958 = ~n10954 & ~n10953;
  assign n10956 = ~n12346 & ~n11290;
  assign n10955 = ~n12092 & ~n12345;
  assign n10957 = ~n10956 & ~n10955;
  assign U3127 = ~n10958 | ~n10957;
  assign n10962 = ~n11699 & ~n12345;
  assign n10960 = ~n12350 | ~n11247;
  assign n10959 = ~INSTQUEUE_REG_3__3__SCAN_IN | ~n11248;
  assign n10961 = ~n10960 | ~n10959;
  assign n10966 = ~n10962 & ~n10961;
  assign n10964 = ~n12346 & ~n11253;
  assign n10963 = ~n12537 & ~n12347;
  assign n10965 = ~n10964 & ~n10963;
  assign U3047 = ~n10966 | ~n10965;
  assign n10972 = ~n11874 & ~n12357;
  assign n10968 = ~n12358 & ~n11300;
  assign n10967 = ~n11301 & ~n12359;
  assign n10970 = ~n10968 & ~n10967;
  assign n10969 = ~n7006 | ~n10615;
  assign n10971 = ~n10970 | ~n10969;
  assign n10974 = ~n10972 & ~n10971;
  assign n10973 = ~INSTQUEUE_REG_11__4__SCAN_IN | ~n11295;
  assign U3112 = ~n10974 | ~n10973;
  assign n10980 = ~n12239 & ~n12359;
  assign n10976 = ~n12358 & ~n11311;
  assign n10975 = ~n12126 & ~n12357;
  assign n10978 = ~n10976 & ~n10975;
  assign n10977 = ~n7006 | ~n10585;
  assign n10979 = ~n10978 | ~n10977;
  assign n10982 = ~n10980 & ~n10979;
  assign n10981 = ~INSTQUEUE_REG_15__4__SCAN_IN | ~n11306;
  assign U3144 = ~n10982 | ~n10981;
  assign n10985 = n10984 | n10983;
  assign n10988 = n10987 | n10986;
  assign n10991 = ~EBX_REG_10__SCAN_IN | ~n13560;
  assign U2849 = ~n10992 | ~n10991;
  assign n10993 = ~n8268 & ~n13391;
  assign n10995 = ~n12099 | ~DATAI_10_;
  assign U2881 = ~n10996 | ~n10995;
  assign n11000 = ~n11301 & ~n12536;
  assign n10998 = ~n12538 | ~n10893;
  assign n10997 = ~INSTQUEUE_REG_10__5__SCAN_IN | ~n11178;
  assign n11004 = ~n11000 & ~n10999;
  assign n11002 = ~n12543 & ~n11171;
  assign n11001 = ~n11383 & ~n12544;
  assign n11003 = ~n11002 & ~n11001;
  assign U3105 = ~n11004 | ~n11003;
  assign n11008 = ~n11301 & ~n12357;
  assign n11006 = ~n7006 | ~n10893;
  assign n11005 = ~INSTQUEUE_REG_10__4__SCAN_IN | ~n11178;
  assign n11012 = ~n11008 & ~n11007;
  assign n11010 = ~n12358 & ~n11171;
  assign n11009 = ~n11383 & ~n12359;
  assign n11011 = ~n11010 & ~n11009;
  assign U3104 = ~n11012 | ~n11011;
  assign n11016 = ~n11301 & ~n12370;
  assign n11014 = ~n7011 | ~n10893;
  assign n11013 = ~INSTQUEUE_REG_10__7__SCAN_IN | ~n11178;
  assign n11015 = ~n11014 | ~n11013;
  assign n11020 = ~n11016 & ~n11015;
  assign n11018 = ~n12369 & ~n11171;
  assign n11017 = ~n11383 & ~n12368;
  assign n11019 = ~n11018 & ~n11017;
  assign U3107 = ~n11020 | ~n11019;
  assign n11022 = ~EAX_REG_11__SCAN_IN | ~n13178;
  assign n11021 = ~n12099 | ~DATAI_11_;
  assign n11026 = n11022 & n11021;
  assign U2880 = ~n11026 | ~n11025;
  assign n11036 = ~n12634 & ~n13316;
  assign n11032 = ~n13551 & ~n13451;
  assign n11030 = n11028 | n11027;
  assign n11031 = ~n13465 & ~n11397;
  assign n11034 = ~n11032 & ~n11031;
  assign n11033 = ~n13467 | ~PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n11398 = ~n13491 | ~REIP_REG_5__SCAN_IN;
  assign U2981 = ~n11037 | ~n11398;
  assign n11043 = ~n12183 & ~n12370;
  assign n11039 = ~n12369 & ~n11275;
  assign n11038 = ~n11707 & ~n12368;
  assign n11041 = ~n11039 & ~n11038;
  assign n11040 = ~n7011 | ~n11269;
  assign n11042 = ~n11041 | ~n11040;
  assign n11045 = ~n11043 & ~n11042;
  assign n11044 = ~INSTQUEUE_REG_5__7__SCAN_IN | ~n11270;
  assign U3067 = ~n11045 | ~n11044;
  assign n11049 = ~n12092 & ~n12357;
  assign n11047 = ~n7006 | ~n11284;
  assign n11046 = ~INSTQUEUE_REG_13__4__SCAN_IN | ~n11285;
  assign n11048 = ~n11047 | ~n11046;
  assign n11053 = ~n11049 & ~n11048;
  assign n11051 = ~n12358 & ~n11290;
  assign n11050 = ~n11872 & ~n12359;
  assign n11052 = ~n11051 & ~n11050;
  assign U3128 = ~n11053 | ~n11052;
  assign n11057 = ~n12183 & ~n12357;
  assign n11055 = ~n7006 | ~n11269;
  assign n11054 = ~INSTQUEUE_REG_5__4__SCAN_IN | ~n11270;
  assign n11056 = ~n11055 | ~n11054;
  assign n11061 = ~n11057 & ~n11056;
  assign n11059 = ~n12358 & ~n11275;
  assign n11058 = ~n11707 & ~n12359;
  assign n11060 = ~n11059 & ~n11058;
  assign U3064 = ~n11061 | ~n11060;
  assign n11065 = ~n12561 & ~n12357;
  assign n11063 = ~n7006 | ~n11258;
  assign n11062 = ~INSTQUEUE_REG_1__4__SCAN_IN | ~n11259;
  assign n11064 = ~n11063 | ~n11062;
  assign n11069 = ~n11065 & ~n11064;
  assign n11067 = ~n12358 & ~n11264;
  assign n11066 = ~n12128 & ~n12359;
  assign n11068 = ~n11067 & ~n11066;
  assign U3032 = ~n11069 | ~n11068;
  assign n11073 = ~n11699 & ~n12357;
  assign n11071 = ~n7006 | ~n11247;
  assign n11070 = ~INSTQUEUE_REG_3__4__SCAN_IN | ~n11248;
  assign n11072 = ~n11071 | ~n11070;
  assign n11077 = ~n11073 & ~n11072;
  assign n11075 = ~n12358 & ~n11253;
  assign n11074 = ~n12537 & ~n12359;
  assign n11076 = ~n11075 & ~n11074;
  assign U3048 = ~n11077 | ~n11076;
  assign n11081 = ~n12267 & ~n12359;
  assign n11079 = ~n11357 | ~n7006;
  assign n11078 = ~INSTQUEUE_REG_7__4__SCAN_IN | ~n11358;
  assign n11080 = ~n11079 | ~n11078;
  assign n11085 = ~n11081 & ~n11080;
  assign n11083 = ~n12358 & ~n11363;
  assign n11082 = ~n11606 & ~n12357;
  assign n11084 = ~n11083 & ~n11082;
  assign U3080 = ~n11085 | ~n11084;
  assign n11089 = ~EBX_REG_11__SCAN_IN | ~n13560;
  assign n11091 = n11089 & n11088;
  assign U2848 = ~n11091 | ~n11090;
  assign n11102 = ~n13504 & ~n11093;
  assign n11096 = ~n13490 & ~n11713;
  assign n11095 = ~n11094;
  assign n11100 = ~n11096 & ~n11095;
  assign n11097 = ~INSTADDRPOINTER_REG_0__SCAN_IN | ~n13299;
  assign n11098 = ~n11097 | ~n13043;
  assign n11099 = ~n11098 | ~n11578;
  assign n11101 = ~n11100 | ~n11099;
  assign U3017 = ~n11104 | ~n11103;
  assign n11110 = ~n11614 & ~n12368;
  assign n11106 = ~n12369 & ~n11382;
  assign n11105 = ~n11383 & ~n12370;
  assign n11108 = ~n11106 & ~n11105;
  assign n11107 = ~n11376 | ~n7011;
  assign n11109 = ~n11108 | ~n11107;
  assign n11112 = ~n11110 & ~n11109;
  assign n11111 = ~INSTQUEUE_REG_9__7__SCAN_IN | ~n11377;
  assign U3099 = ~n11112 | ~n11111;
  assign n11116 = ~n11614 & ~n12359;
  assign n11114 = ~n11376 | ~n7006;
  assign n11113 = ~INSTQUEUE_REG_9__4__SCAN_IN | ~n11377;
  assign n11115 = ~n11114 | ~n11113;
  assign n11120 = ~n11116 & ~n11115;
  assign n11118 = ~n12358 & ~n11382;
  assign n11117 = ~n11383 & ~n12357;
  assign n11119 = ~n11118 & ~n11117;
  assign U3096 = ~n11120 | ~n11119;
  assign n11124 = ~n11301 & ~n12549;
  assign n11122 = ~n7010 | ~n10893;
  assign n11121 = ~INSTQUEUE_REG_10__2__SCAN_IN | ~n11178;
  assign n11123 = ~n11122 | ~n11121;
  assign n11128 = ~n11124 & ~n11123;
  assign n11126 = ~n12554 & ~n11171;
  assign n11125 = ~n11383 & ~n12555;
  assign n11127 = ~n11126 & ~n11125;
  assign U3102 = ~n11128 | ~n11127;
  assign n11134 = ~n11874 & ~n12549;
  assign n11130 = ~n12554 & ~n11300;
  assign n11129 = ~n11301 & ~n12555;
  assign n11132 = ~n11130 & ~n11129;
  assign n11131 = ~n7010 | ~n10615;
  assign n11133 = ~n11132 | ~n11131;
  assign n11136 = ~n11134 & ~n11133;
  assign n11135 = ~INSTQUEUE_REG_11__2__SCAN_IN | ~n11295;
  assign U3110 = ~n11136 | ~n11135;
  assign n11142 = ~n12126 & ~n12549;
  assign n11138 = ~n12554 & ~n11311;
  assign n11137 = ~n12239 & ~n12555;
  assign n11140 = ~n11138 & ~n11137;
  assign n11139 = ~n7010 | ~n10585;
  assign n11141 = ~n11140 | ~n11139;
  assign n11144 = ~n11142 & ~n11141;
  assign n11143 = ~INSTQUEUE_REG_15__2__SCAN_IN | ~n11306;
  assign U3142 = ~n11144 | ~n11143;
  assign n11150 = ~n11872 & ~n12555;
  assign n11146 = ~n12554 & ~n11290;
  assign n11145 = ~n12092 & ~n12549;
  assign n11148 = ~n11146 & ~n11145;
  assign n11147 = ~n7010 | ~n11284;
  assign n11149 = ~n11148 | ~n11147;
  assign n11152 = ~n11150 & ~n11149;
  assign n11151 = ~INSTQUEUE_REG_13__2__SCAN_IN | ~n11285;
  assign U3126 = ~n11152 | ~n11151;
  assign n11160 = ~n12183 & ~n12570;
  assign n11154 = ~n12569 & ~n11275;
  assign n11153 = ~n11707 & ~n12560;
  assign n11158 = ~n11154 & ~n11153;
  assign n11157 = ~n7004 | ~n11269;
  assign n11162 = ~n11160 & ~n11159;
  assign n11161 = ~INSTQUEUE_REG_5__6__SCAN_IN | ~n11270;
  assign U3066 = ~n11162 | ~n11161;
  assign n11168 = ~n12561 & ~n12570;
  assign n11164 = ~n12569 & ~n11264;
  assign n11163 = ~n12128 & ~n12560;
  assign n11166 = ~n11164 & ~n11163;
  assign n11165 = ~n7004 | ~n11258;
  assign n11170 = ~n11168 & ~n11167;
  assign n11169 = ~INSTQUEUE_REG_1__6__SCAN_IN | ~n11259;
  assign U3034 = ~n11170 | ~n11169;
  assign n11177 = ~n11301 & ~n12570;
  assign n11173 = ~n12569 & ~n11171;
  assign n11172 = ~n11383 & ~n12560;
  assign n11175 = ~n11173 & ~n11172;
  assign n11174 = ~n7004 | ~n10893;
  assign n11176 = ~n11175 | ~n11174;
  assign n11180 = ~n11177 & ~n11176;
  assign n11179 = ~INSTQUEUE_REG_10__6__SCAN_IN | ~n11178;
  assign U3106 = ~n11180 | ~n11179;
  assign n11186 = ~n11699 & ~n12570;
  assign n11182 = ~n12569 & ~n11253;
  assign n11181 = ~n12537 & ~n12560;
  assign n11184 = ~n11182 & ~n11181;
  assign n11183 = ~n7004 | ~n11247;
  assign n11188 = ~n11186 & ~n11185;
  assign n11187 = ~INSTQUEUE_REG_3__6__SCAN_IN | ~n11248;
  assign U3050 = ~n11188 | ~n11187;
  assign n11192 = ~n12561 & ~n12370;
  assign n11190 = ~n7011 | ~n11258;
  assign n11189 = ~INSTQUEUE_REG_1__7__SCAN_IN | ~n11259;
  assign n11191 = ~n11190 | ~n11189;
  assign n11196 = ~n11192 & ~n11191;
  assign n11194 = ~n12369 & ~n11264;
  assign n11193 = ~n12128 & ~n12368;
  assign n11195 = ~n11194 & ~n11193;
  assign U3035 = ~n11196 | ~n11195;
  assign n11200 = ~n11874 & ~n12370;
  assign n11198 = ~n7011 | ~n10615;
  assign n11197 = ~INSTQUEUE_REG_11__7__SCAN_IN | ~n11295;
  assign n11199 = ~n11198 | ~n11197;
  assign n11204 = ~n11200 & ~n11199;
  assign n11202 = ~n12369 & ~n11300;
  assign n11201 = ~n11301 & ~n12368;
  assign n11203 = ~n11202 & ~n11201;
  assign U3115 = ~n11204 | ~n11203;
  assign n11208 = ~n11872 & ~n12368;
  assign n11206 = ~n7011 | ~n11284;
  assign n11205 = ~INSTQUEUE_REG_13__7__SCAN_IN | ~n11285;
  assign n11207 = ~n11206 | ~n11205;
  assign n11212 = ~n11208 & ~n11207;
  assign n11210 = ~n12369 & ~n11290;
  assign n11209 = ~n12092 & ~n12370;
  assign n11211 = ~n11210 & ~n11209;
  assign U3131 = ~n11212 | ~n11211;
  assign n11216 = ~n12239 & ~n12368;
  assign n11214 = ~n7011 | ~n10585;
  assign n11213 = ~INSTQUEUE_REG_15__7__SCAN_IN | ~n11306;
  assign n11215 = ~n11214 | ~n11213;
  assign n11220 = ~n11216 & ~n11215;
  assign n11218 = ~n12369 & ~n11311;
  assign n11217 = ~n12126 & ~n12370;
  assign n11219 = ~n11218 & ~n11217;
  assign U3147 = ~n11220 | ~n11219;
  assign n11224 = ~n11699 & ~n12370;
  assign n11222 = ~n7011 | ~n11247;
  assign n11221 = ~INSTQUEUE_REG_3__7__SCAN_IN | ~n11248;
  assign n11223 = ~n11222 | ~n11221;
  assign n11228 = ~n11224 & ~n11223;
  assign n11226 = ~n12369 & ~n11253;
  assign n11225 = ~n12537 & ~n12368;
  assign n11227 = ~n11226 & ~n11225;
  assign U3051 = ~n11228 | ~n11227;
  assign n11232 = ~n11606 & ~n12370;
  assign n11230 = ~n11357 | ~n7011;
  assign n11229 = ~INSTQUEUE_REG_7__7__SCAN_IN | ~n11358;
  assign n11231 = ~n11230 | ~n11229;
  assign n11236 = ~n11232 & ~n11231;
  assign n11234 = ~n12369 & ~n11363;
  assign n11233 = ~n12267 & ~n12368;
  assign n11235 = ~n11234 & ~n11233;
  assign U3083 = ~n11236 | ~n11235;
  assign n11242 = n11240 | n11239;
  assign n11245 = ~EBX_REG_12__SCAN_IN | ~n13560;
  assign U2847 = ~n11246 | ~n11245;
  assign n11252 = ~n12537 & ~n12555;
  assign n11250 = ~n7010 | ~n11247;
  assign n11249 = ~INSTQUEUE_REG_3__2__SCAN_IN | ~n11248;
  assign n11251 = ~n11250 | ~n11249;
  assign n11257 = ~n11252 & ~n11251;
  assign n11255 = ~n12554 & ~n11253;
  assign n11254 = ~n11699 & ~n12549;
  assign n11256 = ~n11255 & ~n11254;
  assign U3046 = ~n11257 | ~n11256;
  assign n11263 = ~n12561 & ~n12549;
  assign n11261 = ~n7010 | ~n11258;
  assign n11260 = ~INSTQUEUE_REG_1__2__SCAN_IN | ~n11259;
  assign n11262 = ~n11261 | ~n11260;
  assign n11268 = ~n11263 & ~n11262;
  assign n11266 = ~n12554 & ~n11264;
  assign n11265 = ~n12128 & ~n12555;
  assign n11267 = ~n11266 & ~n11265;
  assign U3030 = ~n11268 | ~n11267;
  assign n11274 = ~n12183 & ~n12549;
  assign n11272 = ~n7010 | ~n11269;
  assign n11271 = ~INSTQUEUE_REG_5__2__SCAN_IN | ~n11270;
  assign n11273 = ~n11272 | ~n11271;
  assign n11279 = ~n11274 & ~n11273;
  assign n11277 = ~n12554 & ~n11275;
  assign n11276 = ~n11707 & ~n12555;
  assign n11278 = ~n11277 & ~n11276;
  assign U3062 = ~n11279 | ~n11278;
  assign n11281 = ~n8377 & ~n13391;
  assign n11282 = ~n12099 | ~DATAI_12_;
  assign U2879 = ~n11283 | ~n11282;
  assign n11289 = ~n12092 & ~n12570;
  assign n11287 = ~n7004 | ~n11284;
  assign n11286 = ~INSTQUEUE_REG_13__6__SCAN_IN | ~n11285;
  assign n11288 = ~n11287 | ~n11286;
  assign n11294 = ~n11289 & ~n11288;
  assign n11292 = ~n12569 & ~n11290;
  assign n11291 = ~n11872 & ~n12560;
  assign n11293 = ~n11292 & ~n11291;
  assign U3130 = ~n11294 | ~n11293;
  assign n11299 = ~n11874 & ~n12570;
  assign n11297 = ~n7004 | ~n10615;
  assign n11296 = ~INSTQUEUE_REG_11__6__SCAN_IN | ~n11295;
  assign n11298 = ~n11297 | ~n11296;
  assign n11305 = ~n11299 & ~n11298;
  assign n11303 = ~n12569 & ~n11300;
  assign n11302 = ~n11301 & ~n12560;
  assign n11304 = ~n11303 & ~n11302;
  assign U3114 = ~n11305 | ~n11304;
  assign n11310 = ~n12239 & ~n12560;
  assign n11308 = ~n7004 | ~n10585;
  assign n11307 = ~INSTQUEUE_REG_15__6__SCAN_IN | ~n11306;
  assign n11309 = ~n11308 | ~n11307;
  assign n11315 = ~n11310 & ~n11309;
  assign n11313 = ~n12569 & ~n11311;
  assign n11312 = ~n12126 & ~n12570;
  assign n11314 = ~n11313 & ~n11312;
  assign U3146 = ~n11315 | ~n11314;
  assign n11323 = ~INSTADDRPOINTER_REG_3__SCAN_IN & ~n11430;
  assign n13558 = n11319 ^ n11318;
  assign n11320 = ~n13558 | ~n13507;
  assign n11322 = ~n11321 | ~n11320;
  assign n11337 = ~n11323 & ~n11322;
  assign n11568 = ~n8001 & ~n11325;
  assign n11331 = ~n11324 & ~n11568;
  assign n11327 = n13043 | n11325;
  assign n11329 = ~n11327 | ~n13298;
  assign n11328 = ~n13374 | ~n11569;
  assign n11335 = ~n11332 & ~n11427;
  assign n11334 = ~n13504 & ~n11333;
  assign n11336 = ~n11335 & ~n11334;
  assign U3015 = ~n11337 | ~n11336;
  assign n11343 = ~n13545 & ~n13451;
  assign n11341 = n11339 | n11338;
  assign n11342 = ~n13465 & ~n12199;
  assign n11345 = ~n11343 & ~n11342;
  assign n12204 = ~n13491 | ~REIP_REG_6__SCAN_IN;
  assign U2980 = ~n11348 | ~n12204;
  assign n11352 = ~n12267 & ~n12555;
  assign n11350 = ~n11357 | ~n7010;
  assign n11349 = ~INSTQUEUE_REG_7__2__SCAN_IN | ~n11358;
  assign n11351 = ~n11350 | ~n11349;
  assign n11356 = ~n11352 & ~n11351;
  assign n11354 = ~n12554 & ~n11363;
  assign n11353 = ~n11606 & ~n12549;
  assign n11355 = ~n11354 & ~n11353;
  assign U3078 = ~n11356 | ~n11355;
  assign n11362 = ~n11606 & ~n12570;
  assign n11360 = ~n11357 | ~n7004;
  assign n11359 = ~INSTQUEUE_REG_7__6__SCAN_IN | ~n11358;
  assign n11367 = ~n11362 & ~n11361;
  assign n11365 = ~n12569 & ~n11363;
  assign n11364 = ~n12267 & ~n12560;
  assign n11366 = ~n11365 & ~n11364;
  assign U3082 = ~n11367 | ~n11366;
  assign n11371 = ~n11614 & ~n12555;
  assign n11369 = ~n11376 | ~n7010;
  assign n11368 = ~INSTQUEUE_REG_9__2__SCAN_IN | ~n11377;
  assign n11370 = ~n11369 | ~n11368;
  assign n11375 = ~n11371 & ~n11370;
  assign n11373 = ~n12554 & ~n11382;
  assign n11372 = ~n11383 & ~n12549;
  assign n11374 = ~n11373 & ~n11372;
  assign U3094 = ~n11375 | ~n11374;
  assign n11381 = ~n11614 & ~n12560;
  assign n11379 = ~n11376 | ~n7004;
  assign n11378 = ~INSTQUEUE_REG_9__6__SCAN_IN | ~n11377;
  assign n11387 = ~n11381 & ~n11380;
  assign n11385 = ~n12569 & ~n11382;
  assign n11384 = ~n11383 & ~n12570;
  assign n11386 = ~n11385 & ~n11384;
  assign U3098 = ~n11387 | ~n11386;
  assign n11389 = ~n9141 | ~n11388;
  assign n11394 = ~n11390 | ~n11389;
  assign n11392 = ~n13507 | ~n11954;
  assign n11391 = ~INSTADDRPOINTER_REG_0__SCAN_IN | ~n13298;
  assign n11393 = ~n11392 | ~n11391;
  assign U3018 = ~n11396 | ~n11395;
  assign n11400 = ~n13504 & ~n11397;
  assign n11399 = ~n11398;
  assign n11404 = ~n11400 & ~n11399;
  assign n13552 = n11402 ^ n11401;
  assign n11403 = ~n13507 | ~n13552;
  assign n11409 = ~n13049 & ~n11406;
  assign n11408 = ~n13045 & ~n11407;
  assign n11410 = ~n11409 & ~n11408;
  assign U3013 = ~n11412 | ~n11411;
  assign n11418 = ~n13539 & ~n13451;
  assign n11416 = n11414 | n11413;
  assign n11549 = ~n13491 | ~REIP_REG_7__SCAN_IN;
  assign U2979 = ~n11423 | ~n11549;
  assign n11426 = ~n11424;
  assign n11425 = ~n13490 & ~n11629;
  assign n11439 = ~n11426 & ~n11425;
  assign n11428 = ~INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n11437 = ~n11428 & ~n11427;
  assign n11435 = ~n9141 | ~n11429;
  assign n11431 = ~INSTADDRPOINTER_REG_4__SCAN_IN & ~INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n11433 = ~n11431 & ~n11430;
  assign n11434 = ~n11433 | ~n11432;
  assign U3014 = ~n11439 | ~n11438;
  assign n11455 = ~n11699 & ~n12301;
  assign n11474 = ~n11440;
  assign n11991 = ~n11474 | ~n11441;
  assign n11448 = ~n11991 & ~n12156;
  assign n11450 = ~n12312 & ~n11706;
  assign n11449 = ~n11707 & ~n12313;
  assign n11453 = ~n11450 & ~n11449;
  assign n11452 = ~n12317 | ~n11700;
  assign n11465 = ~n11455 & ~n11454;
  assign n11460 = ~n12324 & ~n11700;
  assign n11462 = n11461 | n11460;
  assign n11983 = ~n11991 | ~STATE2_REG_2__SCAN_IN;
  assign U3052 = ~n11465 | ~n11464;
  assign n11471 = ~n11699 & ~n12555;
  assign n11467 = ~n12554 & ~n11706;
  assign n11466 = ~n11707 & ~n12549;
  assign n11469 = ~n11467 & ~n11466;
  assign n11468 = ~n7010 | ~n11700;
  assign n11473 = ~n11471 & ~n11470;
  assign U3054 = ~n11473 | ~n11472;
  assign n11493 = ~n11614 & ~n12313;
  assign n11487 = ~n11606 & ~n12301;
  assign n11498 = ~n11474 & ~n12146;
  assign n11745 = ~n11498;
  assign n11485 = ~n11745 & ~n12302;
  assign n11482 = ~n11481;
  assign n11486 = ~n11613 & ~n12312;
  assign n11491 = ~n11487 & ~n11486;
  assign n11496 = ~n11489 | ~n11488;
  assign n11490 = ~n11607 | ~n12317;
  assign n11505 = ~n11493 & ~n11492;
  assign n11500 = ~STATE2_REG_3__SCAN_IN | ~n11496;
  assign n11734 = ~n11498 & ~n11497;
  assign n11499 = ~n11734;
  assign n11501 = ~n11500 | ~n11499;
  assign n11504 = ~INSTQUEUE_REG_8__0__SCAN_IN | ~n11608;
  assign U3084 = ~n11505 | ~n11504;
  assign n11511 = ~n11606 & ~n12368;
  assign n11507 = ~n12369 & ~n11613;
  assign n11506 = ~n11614 & ~n12370;
  assign n11509 = ~n11507 & ~n11506;
  assign n11508 = ~n11607 | ~n7011;
  assign n11513 = ~n11511 & ~n11510;
  assign n11512 = ~INSTQUEUE_REG_8__7__SCAN_IN | ~n11608;
  assign U3091 = ~n11513 | ~n11512;
  assign n11519 = ~n11606 & ~n12560;
  assign n11515 = ~n12569 & ~n11613;
  assign n11514 = ~n11614 & ~n12570;
  assign n11517 = ~n11515 & ~n11514;
  assign n11516 = ~n11607 | ~n7004;
  assign n11521 = ~n11519 & ~n11518;
  assign n11520 = ~INSTQUEUE_REG_8__6__SCAN_IN | ~n11608;
  assign U3090 = ~n11521 | ~n11520;
  assign n11527 = ~n11606 & ~n12359;
  assign n11523 = ~n12358 & ~n11613;
  assign n11522 = ~n11614 & ~n12357;
  assign n11525 = ~n11523 & ~n11522;
  assign n11524 = ~n11607 | ~n7006;
  assign n11529 = ~n11527 & ~n11526;
  assign n11528 = ~INSTQUEUE_REG_8__4__SCAN_IN | ~n11608;
  assign U3088 = ~n11529 | ~n11528;
  assign n11535 = ~n11606 & ~n12347;
  assign n11531 = ~n12346 & ~n11613;
  assign n11530 = ~n11614 & ~n12345;
  assign n11533 = ~n11531 & ~n11530;
  assign n11532 = ~n11607 | ~n12350;
  assign n11537 = ~n11535 & ~n11534;
  assign n11536 = ~INSTQUEUE_REG_8__3__SCAN_IN | ~n11608;
  assign U3087 = ~n11537 | ~n11536;
  assign n11543 = ~n11606 & ~n12555;
  assign n11539 = ~n12554 & ~n11613;
  assign n11538 = ~n11614 & ~n12549;
  assign n11541 = ~n11539 & ~n11538;
  assign n11540 = ~n11607 | ~n7010;
  assign n11545 = ~n11543 & ~n11542;
  assign n11544 = ~INSTQUEUE_REG_8__2__SCAN_IN | ~n11608;
  assign U3086 = ~n11545 | ~n11544;
  assign n11551 = ~n13504 & ~n11548;
  assign n11550 = ~n11549;
  assign n11555 = ~n11551 & ~n11550;
  assign n13540 = n11553 ^ n11552;
  assign n11554 = ~n13507 | ~n13540;
  assign n11917 = n13377 | n11561;
  assign U3011 = ~n11563 | ~n11562;
  assign n11580 = ~INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n11564 = ~n13049 & ~INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n11565 = ~n13377 & ~n11564;
  assign n11577 = ~n11580 & ~n11565;
  assign n11566 = ~n12286 | ~n13507;
  assign n11572 = ~n11567 | ~n11566;
  assign n11570 = ~n11569 & ~n11568;
  assign n11571 = ~n11570 & ~n13045;
  assign n11575 = ~n11572 & ~n11571;
  assign n11574 = ~n9141 | ~n11573;
  assign n11581 = ~n11579 & ~n11578;
  assign U3016 = ~n11583 | ~n11582;
  assign n11587 = ~EBX_REG_14__SCAN_IN | ~n13560;
  assign U2845 = ~n11588 | ~n11587;
  assign n11592 = ~n11591 | ~n11590;
  assign n11596 = ~EBX_REG_13__SCAN_IN | ~n13560;
  assign U2846 = ~n11597 | ~n11596;
  assign n11601 = ~n11606 & ~n12333;
  assign n11599 = ~n11607 | ~n12338;
  assign n11598 = ~INSTQUEUE_REG_8__1__SCAN_IN | ~n11608;
  assign n11600 = ~n11599 | ~n11598;
  assign n11605 = ~n11601 & ~n11600;
  assign n11603 = ~n12334 & ~n11613;
  assign n11602 = ~n11614 & ~n12335;
  assign n11604 = ~n11603 & ~n11602;
  assign U3085 = ~n11605 | ~n11604;
  assign n11612 = ~n11606 & ~n12544;
  assign n11610 = ~n11607 | ~n12538;
  assign n11609 = ~INSTQUEUE_REG_8__5__SCAN_IN | ~n11608;
  assign n11611 = ~n11610 | ~n11609;
  assign n11618 = ~n11612 & ~n11611;
  assign n11616 = ~n12543 & ~n11613;
  assign n11615 = ~n11614 & ~n12536;
  assign n11617 = ~n11616 & ~n11615;
  assign U3089 = ~n11618 | ~n11617;
  assign n11621 = ~n12099 | ~DATAI_14_;
  assign U2877 = ~n11622 | ~n11621;
  assign n11625 = ~n12507;
  assign U3019 = ~n11628 & ~n11859;
  assign n11642 = ~n13329 & ~n11629;
  assign n11635 = ~REIP_REG_4__SCAN_IN & ~n11630;
  assign n11633 = ~n13334 | ~PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n11634 = ~n12805 | ~n11633;
  assign n11640 = ~n11635 & ~n11634;
  assign n11639 = ~n11638 | ~n12587;
  assign n11641 = ~n11640 | ~n11639;
  assign n11644 = ~n11642 & ~n11641;
  assign n11643 = ~EBX_REG_4__SCAN_IN | ~n13335;
  assign n11651 = ~n11645 | ~n13197;
  assign n11650 = ~n12298 | ~n11649;
  assign U2823 = ~n11658 | ~n11657;
  assign n11662 = ~n11699 & ~n12333;
  assign n11660 = ~n12338 | ~n11700;
  assign n11664 = ~n12334 & ~n11706;
  assign n11663 = ~n11707 & ~n12335;
  assign n11665 = ~n11664 & ~n11663;
  assign U3053 = ~n11666 | ~n11665;
  assign n11670 = ~n11699 & ~n12544;
  assign n11668 = ~n12538 | ~n11700;
  assign n11672 = ~n12543 & ~n11706;
  assign n11671 = ~n11707 & ~n12536;
  assign n11673 = ~n11672 & ~n11671;
  assign U3057 = ~n11674 | ~n11673;
  assign n11678 = ~n11699 & ~n12347;
  assign n11676 = ~n12350 | ~n11700;
  assign n11680 = ~n12346 & ~n11706;
  assign n11679 = ~n11707 & ~n12345;
  assign n11681 = ~n11680 & ~n11679;
  assign U3055 = ~n11682 | ~n11681;
  assign n11686 = ~n11699 & ~n12359;
  assign n11684 = ~n7006 | ~n11700;
  assign n11688 = ~n12358 & ~n11706;
  assign n11687 = ~n11707 & ~n12357;
  assign n11689 = ~n11688 & ~n11687;
  assign U3056 = ~n11690 | ~n11689;
  assign n11694 = ~n11699 & ~n12368;
  assign n11692 = ~n7011 | ~n11700;
  assign n11696 = ~n12369 & ~n11706;
  assign n11695 = ~n11707 & ~n12370;
  assign n11697 = ~n11696 & ~n11695;
  assign U3059 = ~n11698 | ~n11697;
  assign n11705 = ~n11699 & ~n12560;
  assign n11703 = ~n7004 | ~n11700;
  assign n11709 = ~n12569 & ~n11706;
  assign n11708 = ~n11707 & ~n12570;
  assign n11710 = ~n11709 & ~n11708;
  assign U3058 = ~n11711 | ~n11710;
  assign n11727 = ~n12635 & ~n11712;
  assign n11723 = ~n13329 & ~n11713;
  assign n11716 = ~REIP_REG_1__SCAN_IN | ~n11714;
  assign n11715 = ~n13334 | ~PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n11721 = ~n11716 | ~n11715;
  assign n11719 = ~n12307 & ~n11717;
  assign n11720 = n11719 | n11718;
  assign n11722 = n11721 | n11720;
  assign n11725 = ~n11723 & ~n11722;
  assign n11724 = ~n13335 | ~EBX_REG_1__SCAN_IN;
  assign n11726 = ~n11725 | ~n11724;
  assign n11728 = n13333 | PHYADDRPOINTER_REG_1__SCAN_IN;
  assign U2826 = ~n11729 | ~n11728;
  assign n11742 = ~n11872 & ~n12536;
  assign n11740 = ~n12538 | ~n11877;
  assign n11736 = ~n12324 & ~n11877;
  assign n11751 = ~n11742 & ~n11741;
  assign n11746 = ~n11745 & ~n12156;
  assign n11749 = ~n12543 & ~n11873;
  assign n11748 = ~n11874 & ~n12544;
  assign n11750 = ~n11749 & ~n11748;
  assign U3121 = ~n11751 | ~n11750;
  assign n11754 = ~n11753 & ~n13391;
  assign n11756 = ~n12099 | ~DATAI_13_;
  assign U2878 = ~n11757 | ~n11756;
  assign n11760 = n11759 | n11758;
  assign n11889 = ~n13491 | ~REIP_REG_8__SCAN_IN;
  assign U2978 = ~n11768 | ~n11889;
  assign n11772 = ~n11872 & ~n12345;
  assign n11770 = ~n12350 | ~n11877;
  assign n11776 = ~n11772 & ~n11771;
  assign n11774 = ~n12346 & ~n11873;
  assign n11773 = ~n11874 & ~n12347;
  assign n11775 = ~n11774 & ~n11773;
  assign U3119 = ~n11776 | ~n11775;
  assign n11780 = ~n11872 & ~n12357;
  assign n11778 = ~n7006 | ~n11877;
  assign n11777 = ~INSTQUEUE_REG_12__4__SCAN_IN | ~n11882;
  assign n11784 = ~n11780 & ~n11779;
  assign n11782 = ~n12358 & ~n11873;
  assign n11781 = ~n11874 & ~n12359;
  assign n11783 = ~n11782 & ~n11781;
  assign U3120 = ~n11784 | ~n11783;
  assign n11788 = ~n11872 & ~n12370;
  assign n11786 = ~n7011 | ~n11877;
  assign n11785 = ~INSTQUEUE_REG_12__7__SCAN_IN | ~n11882;
  assign n11792 = ~n11788 & ~n11787;
  assign n11790 = ~n12369 & ~n11873;
  assign n11789 = ~n11874 & ~n12368;
  assign n11791 = ~n11790 & ~n11789;
  assign U3123 = ~n11792 | ~n11791;
  assign n11796 = ~n11872 & ~n12549;
  assign n11794 = ~n7010 | ~n11877;
  assign n11793 = ~INSTQUEUE_REG_12__2__SCAN_IN | ~n11882;
  assign n11800 = ~n11796 & ~n11795;
  assign n11798 = ~n12554 & ~n11873;
  assign n11797 = ~n11874 & ~n12555;
  assign n11799 = ~n11798 & ~n11797;
  assign U3118 = ~n11800 | ~n11799;
  assign n11804 = ~n11872 & ~n12570;
  assign n11802 = ~n7004 | ~n11877;
  assign n11801 = ~INSTQUEUE_REG_12__6__SCAN_IN | ~n11882;
  assign n11808 = ~n11804 & ~n11803;
  assign n11806 = ~n12569 & ~n11873;
  assign n11805 = ~n11874 & ~n12560;
  assign n11807 = ~n11806 & ~n11805;
  assign U3122 = ~n11808 | ~n11807;
  assign n11812 = ~n11810 | ~n11809;
  assign n11811 = ~n7990 | ~n11851;
  assign n11815 = ~n11812 | ~n11811;
  assign n11853 = ~n11813 & ~STATE2_REG_3__SCAN_IN;
  assign n11822 = ~n11853;
  assign n11814 = ~n7936 | ~n11822;
  assign n11816 = ~n11815 | ~n11814;
  assign U3464 = ~n11818 | ~n11817;
  assign n11819 = ~n7990 | ~STATEBS16_REG_SCAN_IN;
  assign n11821 = ~n11820 ^ n11819;
  assign n11824 = ~n11821 | ~n12305;
  assign n11823 = ~n12287 | ~n11822;
  assign n11825 = ~n11824 | ~n11823;
  assign U3463 = ~n11827 | ~n11826;
  assign n11829 = ~n11828 & ~n11853;
  assign n11832 = ~n11830 & ~n11829;
  assign U3465 = ~n11835 | ~n11834;
  assign n11837 = ~n12390 | ~n13472;
  assign n11836 = ~PHYADDRPOINTER_REG_9__SCAN_IN | ~n13467;
  assign U2977 = ~n11844 | ~n11843;
  assign n11848 = ~n11846 | ~n11845;
  assign n11850 = ~n11848 | ~n11847;
  assign n11858 = ~n11850 | ~n11849;
  assign n11856 = ~n11852 & ~n11851;
  assign n11855 = ~n11854 & ~n11853;
  assign n11857 = ~n11856 & ~n11855;
  assign n11860 = ~n11858 | ~n11857;
  assign U3462 = ~n11863 | ~n11862;
  assign n11869 = ~n11872 & ~n12313;
  assign n11865 = ~n12312 & ~n11873;
  assign n11864 = ~n11874 & ~n12301;
  assign n11867 = ~n11865 & ~n11864;
  assign n11866 = ~n12317 | ~n11877;
  assign n11871 = ~n11869 & ~n11868;
  assign U3116 = ~n11871 | ~n11870;
  assign n11881 = ~n11872 & ~n12335;
  assign n11876 = ~n12334 & ~n11873;
  assign n11875 = ~n11874 & ~n12333;
  assign n11879 = ~n11876 & ~n11875;
  assign n11878 = ~n12338 | ~n11877;
  assign n11884 = ~n11881 & ~n11880;
  assign U3117 = ~n11884 | ~n11883;
  assign n13534 = n11887 ^ n11886;
  assign n11888 = ~n13534 | ~n13507;
  assign n11895 = ~n11894 & ~n11917;
  assign U3010 = ~n11899 | ~n11898;
  assign n11910 = ~n12946 & ~n12434;
  assign n11906 = ~n13329 & ~n12490;
  assign n11900 = ~n12617 | ~n11911;
  assign n11902 = ~n11901 & ~n12379;
  assign n11904 = ~n11902 & ~n12726;
  assign n11903 = ~n13334 | ~PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n11905 = ~n11904 | ~n11903;
  assign n11908 = ~n11906 & ~n11905;
  assign n11907 = ~n13335 | ~EBX_REG_10__SCAN_IN;
  assign n11913 = ~n12433 & ~n13333;
  assign U2817 = ~n11916 | ~n11915;
  assign n11927 = ~n12492 & ~n12502;
  assign n11923 = ~INSTADDRPOINTER_REG_9__SCAN_IN & ~n12499;
  assign n11922 = ~n11921;
  assign n11925 = ~n11923 & ~n11922;
  assign n11924 = ~n13507 | ~n12381;
  assign U3009 = ~n11930 | ~n11929;
  assign n11938 = ~n13329 & ~n12764;
  assign n11933 = ~n11966 | ~REIP_REG_13__SCAN_IN;
  assign n11932 = ~n13335 | ~EBX_REG_13__SCAN_IN;
  assign n11935 = ~n13334 | ~PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n11941 = ~n13330 | ~n11940;
  assign U2814 = ~n11946 | ~n11945;
  assign n11947 = ~n13333 | ~n13199;
  assign n11958 = n12298 & n11948;
  assign n11953 = EBX_REG_0__SCAN_IN & n13335;
  assign n11951 = ~n12926 | ~REIP_REG_0__SCAN_IN;
  assign n11950 = ~n11949 | ~n12587;
  assign n11952 = ~n11951 | ~n11950;
  assign n11956 = ~n11953 & ~n11952;
  assign n11955 = ~n12944 | ~n11954;
  assign U2827 = ~n11960 | ~n11959;
  assign n11962 = ~EBX_REG_31__SCAN_IN | ~n13560;
  assign n11961 = n13528 | n13440;
  assign U2828 = ~n11962 | ~n11961;
  assign n11974 = ~n13329 & ~n12769;
  assign n11964 = ~n12946 & ~n12742;
  assign n11963 = ~n12741 & ~n13333;
  assign n11972 = ~n11964 & ~n11963;
  assign n11965 = ~n13334 | ~PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n11970 = ~n12805 | ~n11965;
  assign n11968 = ~n11966 | ~REIP_REG_12__SCAN_IN;
  assign n11967 = ~n13335 | ~EBX_REG_12__SCAN_IN;
  assign n12398 = ~n11975;
  assign U2815 = ~n11978 | ~n11977;
  assign n11990 = ~n12126 & ~n12544;
  assign n11988 = ~n12538 | ~n12131;
  assign n11982 = n12324 | n12131;
  assign n11984 = ~n11983 | ~n11982;
  assign n12000 = ~n11990 & ~n11989;
  assign n11996 = ~n11991 & ~n12302;
  assign n11993 = ~n11992;
  assign n11998 = ~n12543 & ~n12127;
  assign n11997 = ~n12128 & ~n12536;
  assign n11999 = ~n11998 & ~n11997;
  assign U3025 = ~n12000 | ~n11999;
  assign n12004 = ~n12126 & ~n12347;
  assign n12002 = ~n12350 | ~n12131;
  assign n12008 = ~n12004 & ~n12003;
  assign n12006 = ~n12346 & ~n12127;
  assign n12005 = ~n12128 & ~n12345;
  assign n12007 = ~n12006 & ~n12005;
  assign U3023 = ~n12008 | ~n12007;
  assign n12012 = ~n12126 & ~n12359;
  assign n12010 = ~n7006 | ~n12131;
  assign n12016 = ~n12012 & ~n12011;
  assign n12014 = ~n12358 & ~n12127;
  assign n12013 = ~n12128 & ~n12357;
  assign n12015 = ~n12014 & ~n12013;
  assign U3024 = ~n12016 | ~n12015;
  assign n12020 = ~n12126 & ~n12368;
  assign n12018 = ~n7011 | ~n12131;
  assign n12024 = ~n12020 & ~n12019;
  assign n12022 = ~n12369 & ~n12127;
  assign n12021 = ~n12128 & ~n12370;
  assign n12023 = ~n12022 & ~n12021;
  assign U3027 = ~n12024 | ~n12023;
  assign n12027 = n12026 | n12025;
  assign n12034 = ~EBX_REG_15__SCAN_IN | ~n13335;
  assign n12032 = ~n12031 | ~n12607;
  assign n12036 = ~n13334 | ~PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n12042 = ~n13329 & ~n12045;
  assign n12041 = ~n12827 & ~n13333;
  assign U2812 = ~n12044 | ~n12043;
  assign n12048 = ~EBX_REG_15__SCAN_IN | ~n13560;
  assign U2844 = ~n12049 | ~n12048;
  assign n12062 = ~n12239 & ~n12335;
  assign n12060 = ~n12338 | ~n12243;
  assign n12054 = ~n12324 & ~n12243;
  assign n12071 = ~n12062 & ~n12061;
  assign n12066 = ~n12065 & ~n12156;
  assign n12069 = ~n12334 & ~n12240;
  assign n12068 = ~n12092 & ~n12333;
  assign n12070 = ~n12069 & ~n12068;
  assign U3133 = ~n12071 | ~n12070;
  assign n12075 = ~n12239 & ~n12536;
  assign n12073 = ~n12538 | ~n12243;
  assign n12079 = ~n12075 & ~n12074;
  assign n12077 = ~n12543 & ~n12240;
  assign n12076 = ~n12092 & ~n12544;
  assign n12078 = ~n12077 & ~n12076;
  assign U3137 = ~n12079 | ~n12078;
  assign n12083 = ~n12239 & ~n12370;
  assign n12081 = ~n7011 | ~n12243;
  assign n12080 = ~INSTQUEUE_REG_14__7__SCAN_IN | ~n12248;
  assign n12087 = ~n12083 & ~n12082;
  assign n12085 = ~n12369 & ~n12240;
  assign n12084 = ~n12092 & ~n12368;
  assign n12086 = ~n12085 & ~n12084;
  assign U3139 = ~n12087 | ~n12086;
  assign n12091 = ~n12239 & ~n12570;
  assign n12089 = ~n7004 | ~n12243;
  assign n12088 = ~INSTQUEUE_REG_14__6__SCAN_IN | ~n12248;
  assign n12096 = ~n12091 & ~n12090;
  assign n12094 = ~n12569 & ~n12240;
  assign n12093 = ~n12092 & ~n12560;
  assign n12095 = ~n12094 & ~n12093;
  assign U3138 = ~n12096 | ~n12095;
  assign n12100 = ~n12099 | ~DATAI_15_;
  assign U2876 = ~n12101 | ~n12100;
  assign n12107 = ~n12126 & ~n12333;
  assign n12103 = ~n12334 & ~n12127;
  assign n12102 = ~n12128 & ~n12335;
  assign n12105 = ~n12103 & ~n12102;
  assign n12104 = ~n12338 | ~n12131;
  assign U3021 = ~n12109 | ~n12108;
  assign n12115 = ~n12126 & ~n12301;
  assign n12111 = ~n12312 & ~n12127;
  assign n12110 = ~n12128 & ~n12313;
  assign n12113 = ~n12111 & ~n12110;
  assign n12112 = ~n12317 | ~n12131;
  assign U3020 = ~n12117 | ~n12116;
  assign n12123 = ~n12126 & ~n12555;
  assign n12119 = ~n12554 & ~n12127;
  assign n12118 = ~n12128 & ~n12549;
  assign n12121 = ~n12119 & ~n12118;
  assign n12120 = ~n7010 | ~n12131;
  assign U3022 = ~n12125 | ~n12124;
  assign n12135 = ~n12126 & ~n12560;
  assign n12130 = ~n12569 & ~n12127;
  assign n12129 = ~n12128 & ~n12570;
  assign n12133 = ~n12130 & ~n12129;
  assign n12132 = ~n7004 | ~n12131;
  assign U3026 = ~n12138 | ~n12137;
  assign n12153 = ~n12267 & ~n12536;
  assign n12151 = ~n12538 | ~n12271;
  assign n12143 = ~n12324 & ~n12271;
  assign n12303 = ~n12146 | ~n12145;
  assign n12328 = n12303 & STATE2_REG_2__SCAN_IN;
  assign n12162 = ~n12153 & ~n12152;
  assign n12157 = ~n12303 & ~n12156;
  assign n12160 = ~n12543 & ~n12268;
  assign n12159 = ~n12183 & ~n12544;
  assign n12161 = ~n12160 & ~n12159;
  assign U3073 = ~n12162 | ~n12161;
  assign n12166 = ~n12267 & ~n12345;
  assign n12164 = ~n12350 | ~n12271;
  assign n12170 = ~n12166 & ~n12165;
  assign n12168 = ~n12346 & ~n12268;
  assign n12167 = ~n12183 & ~n12347;
  assign n12169 = ~n12168 & ~n12167;
  assign U3071 = ~n12170 | ~n12169;
  assign n12174 = ~n12267 & ~n12357;
  assign n12172 = ~n7006 | ~n12271;
  assign n12178 = ~n12174 & ~n12173;
  assign n12176 = ~n12358 & ~n12268;
  assign n12175 = ~n12183 & ~n12359;
  assign n12177 = ~n12176 & ~n12175;
  assign U3072 = ~n12178 | ~n12177;
  assign n12182 = ~n12267 & ~n12549;
  assign n12180 = ~n7010 | ~n12271;
  assign n12187 = ~n12182 & ~n12181;
  assign n12185 = ~n12554 & ~n12268;
  assign n12184 = ~n12183 & ~n12555;
  assign n12186 = ~n12185 & ~n12184;
  assign U3070 = ~n12187 | ~n12186;
  assign n12191 = ~n12267 & ~n12570;
  assign n12189 = ~n7004 | ~n12271;
  assign n12188 = ~INSTQUEUE_REG_6__6__SCAN_IN | ~n12276;
  assign n12195 = ~n12191 & ~n12190;
  assign n12193 = ~n12569 & ~n12268;
  assign n12192 = ~n12183 & ~n12560;
  assign n12194 = ~n12193 & ~n12192;
  assign U3074 = ~n12195 | ~n12194;
  assign n12198 = ~n12196 & ~INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n12212 = ~n13504 & ~n12199;
  assign n12205 = ~n12204;
  assign n13546 = n12208 ^ n12207;
  assign n12209 = ~n13507 | ~n13546;
  assign U3012 = ~n12214 | ~n12213;
  assign n12220 = ~n12239 & ~n12313;
  assign n12216 = ~n12312 & ~n12240;
  assign n12215 = ~n12092 & ~n12301;
  assign n12218 = ~n12216 & ~n12215;
  assign n12217 = ~n12317 | ~n12243;
  assign U3132 = ~n12222 | ~n12221;
  assign n12228 = ~n12239 & ~n12345;
  assign n12224 = ~n12346 & ~n12240;
  assign n12223 = ~n12092 & ~n12347;
  assign n12226 = ~n12224 & ~n12223;
  assign n12225 = ~n12350 | ~n12243;
  assign U3135 = ~n12230 | ~n12229;
  assign n12236 = ~n12239 & ~n12357;
  assign n12232 = ~n12358 & ~n12240;
  assign n12231 = ~n12092 & ~n12359;
  assign n12234 = ~n12232 & ~n12231;
  assign n12233 = ~n7006 | ~n12243;
  assign U3136 = ~n12238 | ~n12237;
  assign n12247 = ~n12239 & ~n12549;
  assign n12242 = ~n12554 & ~n12240;
  assign n12241 = ~n12092 & ~n12555;
  assign n12245 = ~n12242 & ~n12241;
  assign n12244 = ~n7010 | ~n12243;
  assign U3134 = ~n12250 | ~n12249;
  assign n12256 = ~n12267 & ~n12313;
  assign n12252 = ~n12312 & ~n12268;
  assign n12251 = ~n12183 & ~n12301;
  assign n12254 = ~n12252 & ~n12251;
  assign n12253 = ~n12317 | ~n12271;
  assign U3068 = ~n12258 | ~n12257;
  assign n12264 = ~n12267 & ~n12335;
  assign n12260 = ~n12334 & ~n12268;
  assign n12259 = ~n12183 & ~n12333;
  assign n12262 = ~n12260 & ~n12259;
  assign n12261 = ~n12338 | ~n12271;
  assign U3069 = ~n12266 | ~n12265;
  assign n12275 = ~n12267 & ~n12370;
  assign n12270 = ~n12369 & ~n12268;
  assign n12269 = ~n12183 & ~n12368;
  assign n12273 = ~n12270 & ~n12269;
  assign n12272 = ~n7011 | ~n12271;
  assign U3075 = ~n12278 | ~n12277;
  assign n12281 = ~n12577 & ~REIP_REG_2__SCAN_IN;
  assign n12279 = ~PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n12280 = ~n13199 & ~n12279;
  assign n12283 = ~n12281 & ~n12280;
  assign n12282 = ~EBX_REG_2__SCAN_IN | ~n13335;
  assign n12291 = ~n12285 & ~n12284;
  assign n12289 = ~n12944 | ~n12286;
  assign n12288 = ~n12287 | ~n12587;
  assign n12290 = ~n12289 | ~n12288;
  assign n12294 = ~n12291 & ~n12290;
  assign n12293 = ~n13197 | ~n12292;
  assign U2825 = ~n12300 | ~n12299;
  assign n12321 = ~n12561 & ~n12301;
  assign n12311 = ~n12303 & ~n12302;
  assign n12315 = ~n12312 & ~n12568;
  assign n12314 = ~n12537 & ~n12313;
  assign n12319 = ~n12315 & ~n12314;
  assign n12318 = ~n12317 | ~n12562;
  assign n12332 = ~n12321 & ~n12320;
  assign n12325 = ~n12324 & ~n12562;
  assign n12327 = n12326 | n12325;
  assign U3036 = ~n12332 | ~n12331;
  assign n12342 = ~n12561 & ~n12333;
  assign n12337 = ~n12334 & ~n12568;
  assign n12336 = ~n12537 & ~n12335;
  assign n12340 = ~n12337 & ~n12336;
  assign n12339 = ~n12338 | ~n12562;
  assign n12344 = ~n12342 & ~n12341;
  assign U3037 = ~n12344 | ~n12343;
  assign n12354 = ~n12537 & ~n12345;
  assign n12349 = ~n12346 & ~n12568;
  assign n12348 = ~n12561 & ~n12347;
  assign n12352 = ~n12349 & ~n12348;
  assign n12351 = ~n12350 | ~n12562;
  assign n12356 = ~n12354 & ~n12353;
  assign U3039 = ~n12356 | ~n12355;
  assign n12365 = ~n12537 & ~n12357;
  assign n12361 = ~n12358 & ~n12568;
  assign n12360 = ~n12561 & ~n12359;
  assign n12363 = ~n12361 & ~n12360;
  assign n12362 = ~n7006 | ~n12562;
  assign n12367 = ~n12365 & ~n12364;
  assign U3040 = ~n12367 | ~n12366;
  assign n12376 = ~n12561 & ~n12368;
  assign n12372 = ~n12369 & ~n12568;
  assign n12371 = ~n12537 & ~n12370;
  assign n12374 = ~n12372 & ~n12371;
  assign n12373 = ~n7011 | ~n12562;
  assign n12378 = ~n12376 & ~n12375;
  assign U3043 = ~n12378 | ~n12377;
  assign n12388 = ~n12380 & ~n12379;
  assign n12383 = ~n12944 | ~n12381;
  assign n12382 = ~n13335 | ~EBX_REG_9__SCAN_IN;
  assign n12384 = ~n12383 | ~n12382;
  assign n12386 = ~n12726 & ~n12384;
  assign n12385 = ~n13334 | ~PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n12393 = ~n12390 | ~n13197;
  assign n12392 = ~n13330 | ~n12391;
  assign U2818 = ~n12397 | ~n12396;
  assign n12399 = ~n12617 | ~n12398;
  assign n12400 = ~REIP_REG_11__SCAN_IN | ~n12399;
  assign n12407 = ~n12400 & ~n12721;
  assign n12402 = ~n12944 | ~n12509;
  assign n12401 = ~n13335 | ~EBX_REG_11__SCAN_IN;
  assign n12403 = ~n12402 | ~n12401;
  assign n12405 = ~n12726 & ~n12403;
  assign n12404 = ~n13334 | ~PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n12409 = ~n13197 | ~n12463;
  assign U2816 = ~n12414 | ~n12413;
  assign n12426 = ~n12946 & ~n13539;
  assign n12416 = ~n13199 & ~n12415;
  assign n12424 = ~n12416 & ~n12726;
  assign n12422 = ~n12418 & ~n12448;
  assign n12420 = ~n12944 | ~n13540;
  assign n12419 = ~n13335 | ~EBX_REG_7__SCAN_IN;
  assign n12421 = ~n12420 | ~n12419;
  assign n12423 = ~n12422 & ~n12421;
  assign n12430 = ~n12427 & ~REIP_REG_7__SCAN_IN;
  assign n12429 = ~n12428 & ~n13333;
  assign U2820 = ~n12432 | ~n12431;
  assign U2976 = ~n12445 | ~n12495;
  assign n12446 = ~n12650 & ~REIP_REG_6__SCAN_IN;
  assign n12460 = ~n12448 & ~n12447;
  assign n12451 = ~n12946 & ~n13545;
  assign n12450 = ~n12449 & ~n13333;
  assign n12458 = ~n12451 & ~n12450;
  assign n12452 = ~n13334 | ~PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n12456 = ~n12805 | ~n12452;
  assign n12454 = ~n12944 | ~n13546;
  assign n12453 = ~n13335 | ~EBX_REG_6__SCAN_IN;
  assign n12455 = ~n12454 | ~n12453;
  assign n12457 = ~n12456 & ~n12455;
  assign U2821 = ~n12462 | ~n12461;
  assign n12464 = ~PHYADDRPOINTER_REG_11__SCAN_IN | ~n13467;
  assign U2975 = ~n12475 | ~n12474;
  assign n12479 = ~n12528;
  assign n12482 = ~EBX_REG_16__SCAN_IN | ~n13560;
  assign U2843 = ~n12483 | ~n12482;
  assign n12485 = ~n13177 | ~DATAI_0_;
  assign n12484 = ~n7008 | ~DATAI_16_;
  assign n12488 = ~EAX_REG_16__SCAN_IN | ~n13178;
  assign U2875 = ~n12489 | ~n12488;
  assign n12503 = ~n12502 | ~n12501;
  assign U3008 = ~n12506 | ~n12505;
  assign U3453 = ~n12508 | ~n12507;
  assign n12522 = ~n13049 & ~n12519;
  assign n12521 = ~n13045 & ~n12520;
  assign U3007 = ~n12526 | ~n12525;
  assign n12529 = n12528 | n12527;
  assign n12531 = ~n13177 | ~DATAI_1_;
  assign n12530 = ~n7008 | ~DATAI_17_;
  assign n12534 = ~EAX_REG_17__SCAN_IN | ~n13178;
  assign U2874 = ~n12535 | ~n12534;
  assign n12542 = ~n12537 & ~n12536;
  assign n12540 = ~n12538 | ~n12562;
  assign n12546 = ~n12543 & ~n12568;
  assign n12545 = ~n12561 & ~n12544;
  assign n12547 = ~n12546 & ~n12545;
  assign U3041 = ~n12548 | ~n12547;
  assign n12553 = ~n12537 & ~n12549;
  assign n12551 = ~n7010 | ~n12562;
  assign n12557 = ~n12554 & ~n12568;
  assign n12556 = ~n12561 & ~n12555;
  assign n12558 = ~n12557 & ~n12556;
  assign U3038 = ~n12559 | ~n12558;
  assign n12567 = ~n12561 & ~n12560;
  assign n12565 = ~n7004 | ~n12562;
  assign n12572 = ~n12569 & ~n12568;
  assign n12571 = ~n12537 & ~n12570;
  assign n12573 = ~n12572 & ~n12571;
  assign U3042 = ~n12574 | ~n12573;
  assign n12586 = ~n12575 & ~n13333;
  assign n12582 = ~n13199 & ~n12576;
  assign n12578 = ~REIP_REG_3__SCAN_IN & ~n12577;
  assign n12580 = ~n12578 | ~REIP_REG_2__SCAN_IN;
  assign n12579 = ~n12944 | ~n13558;
  assign n12581 = ~n12580 | ~n12579;
  assign n12584 = ~n12582 & ~n12581;
  assign n12583 = ~n13335 | ~EBX_REG_3__SCAN_IN;
  assign n12589 = ~n12588 | ~n12587;
  assign U2824 = ~n12595 | ~n12594;
  assign n12599 = ~n13329 & ~n12841;
  assign n12597 = ~n13335 | ~EBX_REG_14__SCAN_IN;
  assign n12596 = ~n13334 | ~PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n12614 = ~n12613 | ~n13197;
  assign U2813 = ~n12615 | ~n12614;
  assign n12629 = ~n12616 & ~n13333;
  assign n12625 = ~n12946 & ~n13533;
  assign n12618 = ~n12617 & ~n12721;
  assign n12620 = ~n12618 | ~REIP_REG_8__SCAN_IN;
  assign n12619 = ~n12944 | ~n13534;
  assign n12621 = ~n12620 | ~n12619;
  assign n12623 = ~n12726 & ~n12621;
  assign n12622 = ~n13334 | ~PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n12626 = ~n13335 | ~EBX_REG_8__SCAN_IN;
  assign U2819 = ~n12633 | ~n12632;
  assign n12649 = ~n12634 & ~n13333;
  assign n12645 = ~n12635 & ~n13551;
  assign n12637 = ~n12636 & ~n12721;
  assign n12643 = ~n12637 | ~REIP_REG_5__SCAN_IN;
  assign n12641 = ~n13199 & ~n12638;
  assign n12639 = ~n12944 | ~n13552;
  assign n12640 = ~n12639 | ~n12805;
  assign n12642 = ~n12641 & ~n12640;
  assign U2822 = ~n12653 | ~n12652;
  assign n12657 = ~EAX_REG_18__SCAN_IN | ~n13178;
  assign n12661 = ~n13177 | ~DATAI_2_;
  assign U2873 = ~n12662 | ~n12661;
  assign n12666 = ~n13334 | ~PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n12671 = ~n12805 | ~n12666;
  assign n12668 = ~n13335 | ~EBX_REG_16__SCAN_IN;
  assign U2811 = ~n12679 | ~n12678;
  assign n12682 = ~n12681 | ~n12680;
  assign n12688 = n12683 | n12682;
  assign U3149 = ~n12694 | ~n12693;
  assign n12698 = n13528 | n13059;
  assign n12697 = ~EBX_REG_19__SCAN_IN | ~n13560;
  assign U2840 = ~n12702 | ~n12701;
  assign n12706 = ~REIP_REG_17__SCAN_IN | ~n12705;
  assign n12708 = ~n13199 & ~n12707;
  assign n12710 = ~n12708 & ~n12726;
  assign n12709 = ~n13335 | ~EBX_REG_17__SCAN_IN;
  assign n12719 = n13329 | n13527;
  assign U2810 = ~n12720 | ~n12719;
  assign n12730 = ~n12993 & ~n13333;
  assign n12724 = ~n12810 | ~REIP_REG_18__SCAN_IN;
  assign n12723 = ~n13335 | ~EBX_REG_18__SCAN_IN;
  assign n12727 = ~n13334 | ~PHYADDRPOINTER_REG_18__SCAN_IN;
  assign U2809 = ~n12740 | ~n12739;
  assign U2974 = ~n12753 | ~n12779;
  assign n12757 = ~n12754 | ~n13371;
  assign n12756 = ~n13374 | ~n12755;
  assign U3005 = ~n12768 | ~n12767;
  assign n12772 = ~n12771 | ~n12770;
  assign U3006 = ~n12785 | ~n12784;
  assign n12788 = ~EBX_REG_20__SCAN_IN | ~n13560;
  assign U2839 = ~n12789 | ~n12788;
  assign n12795 = ~n13177 | ~DATAI_3_;
  assign U2872 = ~n12796 | ~n12795;
  assign n12797 = ~EAX_REG_20__SCAN_IN | ~n13178;
  assign n12802 = ~n13177 | ~DATAI_4_;
  assign U2871 = ~n12803 | ~n12802;
  assign n12804 = ~n13334 | ~PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n12809 = ~n12805 | ~n12804;
  assign n12807 = ~n13335 | ~EBX_REG_19__SCAN_IN;
  assign n12806 = ~n13197 | ~n12917;
  assign n12808 = ~n12807 | ~n12806;
  assign n12812 = ~n12809 & ~n12808;
  assign n12814 = n13329 | n13059;
  assign U2808 = ~n12820 | ~n12819;
  assign n12824 = ~n13164 & ~n12821;
  assign n12831 = n12830 | n13465;
  assign U2971 = ~n12832 | ~n12831;
  assign n12843 = ~n12840;
  assign n12846 = n12843 | n12842;
  assign U3004 = ~n12850 | ~n12849;
  assign n12851 = n13560 & EBX_REG_22__SCAN_IN;
  assign U2837 = ~n12855 | ~n12854;
  assign n12857 = n13560 & EBX_REG_23__SCAN_IN;
  assign U2836 = ~n12861 | ~n12860;
  assign n12865 = n13467 & PHYADDRPOINTER_REG_16__SCAN_IN;
  assign U2970 = ~n12872 | ~n12871;
  assign n12876 = n12875 | n12874;
  assign n12877 = n13560 & EBX_REG_24__SCAN_IN;
  assign U2835 = ~n12880 | ~n12879;
  assign n12884 = ~n13560 | ~EBX_REG_25__SCAN_IN;
  assign U2834 = ~n12887 | ~n12886;
  assign n12980 = ~n12889 | ~n12888;
  assign n12892 = n13467 & PHYADDRPOINTER_REG_17__SCAN_IN;
  assign U2969 = ~n12898 | ~n12897;
  assign n12902 = ~n12961;
  assign n12906 = n13177 & DATAI_10_;
  assign n12904 = ~n7008 | ~DATAI_26_;
  assign n12903 = ~n13178 | ~EAX_REG_26__SCAN_IN;
  assign U2865 = ~n12908 | ~n12907;
  assign n12915 = ~n13467 | ~PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n12918 = n13472 & n12917;
  assign U2967 = ~n12921 | ~n12920;
  assign n12922 = n13560 & EBX_REG_26__SCAN_IN;
  assign U2833 = ~n12925 | ~n12924;
  assign n12927 = ~n12926 | ~REIP_REG_24__SCAN_IN;
  assign n12930 = n12929 | REIP_REG_24__SCAN_IN;
  assign U2803 = ~n12943 | ~n12942;
  assign n12952 = n13333 | n12951;
  assign U2802 = ~n12959 | ~n12958;
  assign n13232 = ~n12963 & ~n12962;
  assign n12967 = n13177 & DATAI_11_;
  assign n12965 = ~n7008 | ~DATAI_27_;
  assign n12964 = ~n13178 | ~EAX_REG_27__SCAN_IN;
  assign U2864 = ~n12969 | ~n12968;
  assign n12974 = n13560 & EBX_REG_27__SCAN_IN;
  assign U2832 = ~n12977 | ~n12976;
  assign n12997 = n13115 | n13465;
  assign U2968 = ~n12997 | ~n12996;
  assign U3001 = ~n13011 | ~n13010;
  assign n13015 = n13177 & DATAI_12_;
  assign n13013 = ~n7008 | ~DATAI_28_;
  assign n13012 = ~n13178 | ~EAX_REG_28__SCAN_IN;
  assign U2863 = ~n13017 | ~n13016;
  assign n13018 = n13560 & EBX_REG_28__SCAN_IN;
  assign U2831 = ~n13021 | ~n13020;
  assign n13042 = n13329 | n13022;
  assign n13032 = ~n13199 & ~n13163;
  assign n13025 = ~n13024 | ~n13035;
  assign n13027 = ~n13026 | ~n13025;
  assign n13030 = n13028 | n13027;
  assign n13038 = n13036 | n13035;
  assign U2801 = ~n13042 | ~n13041;
  assign n13047 = ~n13043 & ~INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n13046 = ~n13045 & ~n13044;
  assign n13052 = ~n13047 & ~n13046;
  assign n13050 = ~n13049 & ~n13048;
  assign n13051 = ~n13050 & ~n13377;
  assign n13063 = n13055 | n13054;
  assign U2999 = ~n13063 | ~n13062;
  assign U2800 = n13075 | n13074;
  assign n13084 = n13467 & PHYADDRPOINTER_REG_20__SCAN_IN;
  assign U2966 = ~n13090 | ~n13089;
  assign n13331 = ~n13094 & ~n13093;
  assign n13098 = n13177 & DATAI_13_;
  assign n13096 = ~n7008 | ~DATAI_29_;
  assign n13095 = ~n13178 | ~EAX_REG_29__SCAN_IN;
  assign U2862 = ~n13100 | ~n13099;
  assign n13104 = n13102 | n13101;
  assign n13105 = n13560 & EBX_REG_29__SCAN_IN;
  assign U2830 = ~n13108 | ~n13107;
  assign n13123 = n13110 | n13109;
  assign n13113 = ~n13112 | ~n13111;
  assign n13116 = n13491 & REIP_REG_18__SCAN_IN;
  assign U3000 = ~n13123 | ~n13122;
  assign n13143 = n13130 | n13129;
  assign n13137 = ~n13333 & ~n13133;
  assign n13135 = ~n13334 | ~PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n13134 = ~n13335 | ~EBX_REG_28__SCAN_IN;
  assign U2799 = ~n13143 | ~n13142;
  assign U2965 = ~n13158 | ~n13157;
  assign n13166 = ~n13162;
  assign n13165 = ~n13164 & ~n13163;
  assign n13167 = ~n13166 & ~n13165;
  assign U2960 = ~n13173 | ~n13172;
  assign n13182 = n13177 & DATAI_14_;
  assign n13180 = ~n7008 | ~DATAI_30_;
  assign n13179 = ~n13178 | ~EAX_REG_30__SCAN_IN;
  assign U2861 = ~n13184 | ~n13183;
  assign n13192 = n13560 & EBX_REG_30__SCAN_IN;
  assign U2829 = ~n13195 | ~n13194;
  assign n13198 = ~PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n13208 = ~n13199 & ~n13198;
  assign n13201 = ~n13200 & ~REIP_REG_30__SCAN_IN;
  assign n13203 = ~n13335 | ~EBX_REG_30__SCAN_IN;
  assign U2797 = ~n13214 | ~n13213;
  assign n13231 = n13416 | n13465;
  assign n13223 = n13467 & PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n13226 = ~n13223 & ~n13417;
  assign U2964 = ~n13231 | ~n13230;
  assign n13233 = ~n13467 | ~PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n13236 = ~n13363 | ~n13233;
  assign n13235 = ~n13316 & ~n13234;
  assign n13237 = ~n13236 & ~n13235;
  assign n13242 = ~n13240;
  assign U2959 = ~n13248 | ~n13247;
  assign n13255 = ~n13249;
  assign n13252 = ~n13251 & ~n13250;
  assign n13253 = ~INSTADDRPOINTER_REG_19__SCAN_IN & ~n13252;
  assign n13254 = ~n13253 & ~n13257;
  assign U2998 = ~n13268 | ~n13267;
  assign n13276 = ~n13272 | ~n13481;
  assign n13275 = ~n13274 | ~n13273;
  assign n13277 = ~n13276 & ~n13275;
  assign n13282 = ~INSTADDRPOINTER_REG_26__SCAN_IN | ~INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n13284 = ~n13297 & ~n13282;
  assign n13285 = ~n13284 | ~n13283;
  assign n13436 = ~n13287 | ~n13286;
  assign n13432 = ~INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n13290 = ~n13467 | ~PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n13292 = ~n13306 | ~n13290;
  assign n13291 = ~n13316 & ~n13332;
  assign U2957 = n13296 | n13295;
  assign n13397 = ~n13432 & ~n13297;
  assign n13426 = n13299 | n13298;
  assign n13304 = ~n13396;
  assign U2989 = ~n13311 | ~n13310;
  assign n13313 = ~n13467 | ~PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n13318 = ~n13314 | ~n13313;
  assign n13317 = ~n13316 & ~n13315;
  assign n13321 = n13318 | n13317;
  assign U2963 = ~n13323 | ~n13322;
  assign n13326 = n13325 | REIP_REG_29__SCAN_IN;
  assign n13339 = ~n13333 & ~n13332;
  assign n13337 = ~n13334 | ~PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n13336 = ~n13335 | ~EBX_REG_29__SCAN_IN;
  assign U2798 = ~n13345 | ~n13344;
  assign n13351 = ~n13491 | ~REIP_REG_24__SCAN_IN;
  assign n13350 = ~n13467 | ~PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n13354 = n13351 & n13350;
  assign U2962 = ~n13358 | ~n13357;
  assign n13361 = n13398 | INSTADDRPOINTER_REG_27__SCAN_IN;
  assign U2991 = ~n13369 | ~n13368;
  assign U2997 = ~n13388 | ~n13387;
  assign n13390 = ~n13464 | ~n13389;
  assign n13392 = n13391 | EAX_REG_31__SCAN_IN;
  assign U2860 = ~n13395 | ~n13394;
  assign n13431 = ~INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n13430 = ~n13404 | ~n13403;
  assign U2988 = ~n13409 | ~n13408;
  assign n13482 = ~n13410;
  assign n13411 = ~INSTADDRPOINTER_REG_21__SCAN_IN & ~INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n13412 = ~n13482 & ~n13411;
  assign n13420 = n13490 | n13419;
  assign U2996 = ~n13425 | ~n13424;
  assign n13427 = n13426 & INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n13433 = ~n13432 | ~n13431;
  assign n13435 = ~n13434 & ~n13433;
  assign n13439 = ~n13438 & ~n13437;
  assign n13446 = n13445 | n13444;
  assign U2987 = ~n13449 | ~n13448;
  assign U2956 = n13462 | n13461;
  assign n13470 = n13467 & PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n13469 = ~n13468;
  assign n13474 = ~n13470 & ~n13469;
  assign U2955 = ~n13478 | ~n13477;
  assign n13483 = ~n13481 | ~n13480;
  assign n13485 = ~n13483 | ~n13482;
  assign n13486 = n13485 | n13484;
  assign n13492 = n13491 & REIP_REG_24__SCAN_IN;
  assign U2994 = ~n13499 | ~n13498;
  assign n13502 = n13501 | INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n13511 = ~n13505 & ~n13504;
  assign n13512 = ~n13511 & ~n13510;
  assign U2993 = ~n13513 | ~n13512;
  assign n13516 = ~n13514 & ~D_C_N_REG_SCAN_IN;
  assign n13519 = ~n13516 & ~n13515;
  assign n13518 = ~CODEFETCH_REG_SCAN_IN & ~n13517;
  assign U2791 = n13519 | n13518;
  assign U2841 = n13525 | n13524;
  assign n13530 = n13528 | n13527;
  assign n13529 = ~EBX_REG_17__SCAN_IN | ~n13560;
  assign U2842 = n13532 | n13531;
  assign n13535 = ~EBX_REG_8__SCAN_IN | ~n13560;
  assign U2851 = n13538 | n13537;
  assign n13544 = ~n8806 & ~n13539;
  assign n13541 = ~EBX_REG_7__SCAN_IN | ~n13560;
  assign U2852 = n13544 | n13543;
  assign n13550 = ~n8806 & ~n13545;
  assign n13547 = ~EBX_REG_6__SCAN_IN | ~n13560;
  assign U2853 = n13550 | n13549;
  assign n13556 = ~n8806 & ~n13551;
  assign n13553 = ~EBX_REG_5__SCAN_IN | ~n13560;
  assign U2854 = n13556 | n13555;
  assign n13564 = ~n8806 & ~n13557;
  assign n13561 = ~EBX_REG_3__SCAN_IN | ~n13560;
  assign U2856 = n13564 | n13563;
  assign n13569 = ~n13566 | ~DATAI_15_;
  assign n13568 = ~LWORD_REG_15__SCAN_IN | ~n13567;
  assign U2954 = n13571 | n13570;
endmodule


