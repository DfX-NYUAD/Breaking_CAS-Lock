// Benchmark "b21_C" written by ABC on Thu Mar  5 01:05:11 2020

module b21_C ( 
    P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
    SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_,
    SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_,
    SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
    P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
    P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
    P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
    P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
    P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
    P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
    P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
    P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
    P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
    P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
    P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
    P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
    P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
    P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
    P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
    P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
    P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
    P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
    P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
    P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
    P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
    P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
    P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
    P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN,
    ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
    ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
    ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
    ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
    U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348,
    P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341,
    P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334,
    P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327,
    P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441,
    P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315,
    P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308,
    P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301,
    P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294,
    P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466,
    P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487,
    P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508,
    P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516,
    P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523,
    P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530,
    P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537,
    P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544,
    P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551,
    P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288,
    P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281,
    P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274,
    P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267,
    P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261,
    P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254,
    P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247,
    P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555,
    P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562,
    P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569,
    P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576,
    P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583,
    P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237,
    P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230,
    P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223,
    P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216,
    P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083,
    P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353,
    P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346,
    P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339,
    P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332,
    P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438,
    P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320,
    P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313,
    P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306,
    P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299,
    P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534,
    P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541,
    P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548,
    P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293,
    P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286,
    P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279,
    P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272,
    P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265,
    P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
    P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
    P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566,
    P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573,
    P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580,
    P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151,
    P2_U3966  );
  input  P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_,
    SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
    SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
    SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
    P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
    P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
    P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
    P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
    P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
    P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
    P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
    P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
    P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
    P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
    P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
    P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
    P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
    P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
    P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
    P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
    P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
    P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
    P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
    P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
    P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
    P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
    P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
    P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
    ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
    ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
    ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
    U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348,
    P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341,
    P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334,
    P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327,
    P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441,
    P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315,
    P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308,
    P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301,
    P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294,
    P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466,
    P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487,
    P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508,
    P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516,
    P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523,
    P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530,
    P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537,
    P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544,
    P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551,
    P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288,
    P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281,
    P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274,
    P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267,
    P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261,
    P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254,
    P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247,
    P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555,
    P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562,
    P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569,
    P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576,
    P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583,
    P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237,
    P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230,
    P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223,
    P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216,
    P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083,
    P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353,
    P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346,
    P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339,
    P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332,
    P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438,
    P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320,
    P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313,
    P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306,
    P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299,
    P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534,
    P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541,
    P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548,
    P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293,
    P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286,
    P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279,
    P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272,
    P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265,
    P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
    P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
    P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566,
    P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573,
    P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580,
    P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151,
    P2_U3966;
  wire n15720, n15434, n15465, n17063, n15298, n16449, n11236, n15154,
    n11075, n14968, n16854, n16503, n14908, n14669, n11217, n14590, n14470,
    n14225, n14997, n14048, n16302, n13952, n15914, n14510, n14447, n13350,
    n13117, n10922, n13206, n13024, n12651, n12618, n11296, n9179, n9035,
    n15212, n16491, n10630, n10586, n10639, n10239, n10632, n9106, n10237,
    n10209, n9304, n9092, n9044, n9093, n10261, n11222, n13555, n10973,
    n11232, n11251, n11212, n11012, n11227, n11238, n10891, n10278, n10940,
    n15395, n15634, n10224, n15739, n12522, n14731, n14266, n9169, n16976,
    n13581, n10768, n10771, n10769, n10772, n15960, n9666, n16048, n10578,
    n15160, n16778, n12043, n15201, n17018, n10796, n9112, n9915, n11207,
    n11315, n11191, n11121, n16502, n14216, n16124, n15961, n15850, n15845,
    n11089, n16957, n15763, n15867, n15488, n15369, n13390, n11613, n12117,
    n10309, n9209, n9205, n9138, n12534, n11807, n10256, n9033, n9180,
    n12537, n12806, n15733, n15722, n15782, n16481, n15732, n16477, n15781,
    n17081, n15490, n16037, n15573, n17080, n15703, n16046, n15663, n17077,
    n15572, n16467, n17076, n17034, n16840, n16045, n16044, n15496, n16036,
    n15543, n15368, n15449, n15522, n15349, n15485, n16835, n15346, n15295,
    n16846, n15591, n15365, n16043, n15136, n17032, n15677, n15253, n15618,
    n16834, n15655, n15123, n16965, n15133, n15774, n16845, n15293, n15250,
    n17071, n16459, n16466, n15251, n16849, n15134, n15223, n16964, n15344,
    n15654, n17069, n15292, n11204, n15747, n16464, n15966, n15358, n16961,
    n15222, n15574, n15355, n11184, n15059, n16457, n15248, n15433, n17070,
    n15131, n15840, n15122, n15420, n15049, n15390, n15062, n15656, n15387,
    n15241, n15430, n15617, n16029, n17030, n15129, n15111, n15965, n16960,
    n15416, n16465, n15642, n16458, n16839, n16455, n15556, n16842, n15380,
    n17145, n15048, n16806, n16454, n16958, n16423, n9968, n15334, n15056,
    n15453, n16447, n15968, n15057, n15379, n15210, n15419, n15321, n15266,
    n15959, n16824, n15331, n15037, n16832, n15640, n15055, n15217, n15183,
    n15418, n15771, n15830, n15008, n15958, n15209, n15405, n15265, n15351,
    n11140, n15796, n15005, n16027, n15711, n14966, n15197, n17144, n16451,
    n15554, n15194, n15152, n16805, n16830, n16956, n16446, n16953, n15320,
    n15855, n15955, n11083, n17121, n17067, n15195, n17149, n15213, n16799,
    n17025, n15795, n15375, n16443, n16506, n15769, n15730, n15653, n15002,
    n11342, n15792, n15098, n11065, n16417, n15291, n16529, n15308, n15319,
    n16798, n15483, n17060, n11058, n16444, n15853, n17061, n11139, n15675,
    n15182, n15728, n15780, n15949, n15374, n17124, n16528, n15256, n11322,
    n16505, n11129, n17143, n15481, n15400, n16801, n15023, n17058, n16823,
    n15001, n15651, n11203, n15674, n15181, n11340, n11338, n15672, n15282,
    n14817, n14789, n16504, n15165, n15396, n14820, n15184, n11344, n15948,
    n17142, n15075, n17120, n14958, n17115, n16794, n15953, n16425, n17123,
    n15072, n17108, n15083, n15779, n15414, n14711, n15615, n15394, n14714,
    n17057, n17122, n11066, n15648, n14991, n15759, n14807, n15613, n15879,
    n15304, n14940, n15859, n15069, n14814, n11068, n14943, n15821, n11200,
    n14863, n10741, n15624, n10172, n14788, n15643, n14813, n15662, n15167,
    n17020, n16776, n14777, n14709, n10736, n17117, n15946, n10059, n15110,
    n10170, n15820, n15623, n14992, n16403, n15877, n15569, n15257, n16775,
    n15661, n14937, n15070, n16401, n15157, n15686, n14765, n15702, n15705,
    n14575, n15645, n15876, n11301, n15817, n14929, n14706, n14762, n11268,
    n15109, n15424, n16020, n14922, n15410, n14469, n11288, n15471, n14466,
    n15943, n11292, n17050, n16808, n15685, n15180, n15036, n10685, n17024,
    n16436, n15495, n15700, n11305, n16814, n9998, n14752, n15542, n15341,
    n16400, n14390, n14915, n11044, n15299, n15179, n14759, n14938, n11286,
    n14973, n15494, n11183, n15035, n15699, n15326, n14697, n15590, n15316,
    n14700, n15559, n15189, n15565, n11006, n15245, n15561, n15695, n14554,
    n15066, n14464, n14197, n14989, n15325, n11182, n15588, n15558, n11128,
    n14745, n15464, n15288, n15408, n15540, n15289, n11304, n15448, n15338,
    n11037, n14694, n14101, n14687, n15938, n14615, n11127, n15587, n15186,
    n14760, n14913, n14538, n15521, n14612, n16386, n14665, n15065, n10860,
    n14535, n15063, n14212, n14776, n15584, n15519, n16382, n16763, n14456,
    n16771, n16373, n15274, n15531, n15446, n14682, n14661, n15936, n14037,
    n11034, n16378, n11031, n14609, n14126, n15151, n14488, n14491, n15517,
    n15312, n14209, n15175, n13949, n17051, n15934, n10987, n14987, n15283,
    n16760, n14775, n13942, n14736, n15240, n14695, n16359, n11160, n15239,
    n16865, n15128, n14692, n14658, n14504, n14123, n16362, n14921, n14525,
    n16342, n10062, n14610, n11005, n14113, n15149, n16768, n10023, n15268,
    n10684, n14062, n15932, n15120, n9940, n11161, n14110, n10683, n13810,
    n15022, n15161, n14443, n14485, n15227, n14109, n15118, n10875, n16358,
    n14933, n14195, n14654, n15511, n14121, n14463, n14049, n14320, n15236,
    n14092, n14501, n16762, n14674, n9909, n15930, n15097, n15127, n10980,
    n11115, n14194, n11113, n13937, n11164, n15020, n9937, n10859, n15046,
    n11147, n16351, n9908, n14021, n14108, n15095, n14462, n14597, n16754,
    n15054, n16348, n14074, n15235, n16747, n14317, n10874, n14486, n9911,
    n14435, n14756, n11137, n14263, n14287, n14181, n11002, n15053, n14001,
    n15076, n14008, n11146, n13707, n13712, n14103, n11234, n14982, n14492,
    n15094, n14208, n14904, n15115, n16869, n14288, n14381, n16737, n14017,
    n13921, n16010, n10969, n13805, n14980, n14981, n16741, n14945, n14377,
    n14239, n14957, n14401, n14308, n15000, n9951, n14207, n14369, n14475,
    n16552, n14902, n14378, n14728, n16328, n9903, n10011, n14010, n14178,
    n14016, n14259, n13918, n14592, n15087, n14305, n14161, n13927, n13708,
    n14955, n16317, n16546, n14357, n14398, n14726, n13995, n14944, n13827,
    n10856, n14847, n14786, n14812, n14274, n13899, n14122, n15078, n14358,
    n16316, n14691, n14767, n11094, n14058, n16732, n13981, n13895, n14301,
    n13826, n9920, n13996, n13680, n16321, n14270, n14034, n14175, n14953,
    n13917, n14715, n13910, n11226, n14302, n14163, n14603, n11145, n14234,
    n16738, n11141, n14746, n14255, n9947, n14030, n14157, n14845, n14233,
    n14353, n14651, n13894, n13677, n16292, n13978, n16879, n13992, n9906,
    n9880, n13817, n11174, n14156, n16298, n16290, n13676, n14948, n13896,
    n13972, n14539, n10849, n14916, n14053, n14705, n13334, n14155, n11098,
    n11221, n14479, n14071, n14608, n14889, n14069, n13909, n9853, n14739,
    n9858, n11220, n14026, n16887, n14461, n16878, n11085, n14206, n14748,
    n10995, n14397, n16537, n10602, n14348, n14540, n14149, n14484, n13667,
    n13844, n14515, n11091, n14844, n11087, n14667, n13958, n14783, n14885,
    n14228, n13670, n14235, n14600, n13749, n14883, n14840, n14480, n13500,
    n14516, n14031, n13745, n16540, n14792, n14227, n14267, n9788, n13664,
    n14524, n14598, n14573, n13719, n9792, n9822, n10627, n13497, n14024,
    n14523, n13737, n13802, n10662, n14570, n16885, n16880, n13616, n13955,
    n9893, n14839, n14666, n13404, n16881, n15881, n10731, n14522, n13401,
    n14841, n9759, n13663, n16056, n14343, n14879, n14355, n13701, n14568,
    n14835, n14884, n13417, n11022, n14354, n14878, n13832, n10661, n11021,
    n13396, n13830, n11011, n16699, n14283, n13414, n10590, n9753, n9834,
    n14831, n16940, n14871, n9757, n14279, n14440, n14476, n14870, n14822,
    n14439, n13960, n9831, n9720, n14830, n16279, n16884, n14565, n17002,
    n11016, n16272, n13244, n15905, n15882, n9629, n14106, n14620, n11020,
    n10844, n10577, n14632, n14560, n10665, n14362, n14129, n14617, n14628,
    n13847, n9738, n9715, n16922, n10862, n10562, n9668, n16931, n9731,
    n10978, n16270, n14323, n13597, n9626, n14331, n14082, n14264, n14344,
    n10570, n16700, n16998, n10666, n9663, n13593, n9630, n14132, n14226,
    n10977, n14321, n14329, n13866, n14080, n14184, n16680, n13548, n13763,
    n10664, n13776, n15994, n13867, n14275, n10948, n9700, n13772, n16919,
    n9619, n13876, n13225, n14251, n14252, n13845, n9623, n10835, n13846,
    n10529, n13760, n14130, n13877, n9724, n15992, n10537, n14002, n16252,
    n13982, n13388, n13538, n14159, n9650, n9591, n13759, n10834, n9627,
    n13963, n16643, n13537, n14171, n10511, n13106, n14247, n13566, n13532,
    n12922, n14144, n15839, n16225, n13720, n13565, n16661, n14158, n13459,
    n9606, n13717, n13453, n15902, n12988, n10653, n10833, n15598, n13518,
    n13645, n15716, n15988, n13451, n15989, n9469, n10468, n12976, n9556,
    n13614, n9503, n15986, n12584, n15834, n12915, n9579, n13517, n9551,
    n13688, n13554, n9633, n10938, n13974, n12984, n13646, n13485, n16637,
    n16934, n16987, n13595, n15895, n16914, n12583, n15752, n10934, n13309,
    n10832, n12483, n10392, n12474, n16220, n16203, n16175, n10932, n9466,
    n12472, n9461, n15563, n15890, n13022, n13203, n12309, n10933, n10445,
    n12578, n11316, n12480, n13185, n13173, n15281, n10831, n9486, n13266,
    n15566, n9539, n14047, n15984, n12469, n15486, n12577, n12308, n12479,
    n15888, n15865, n13295, n12372, n10456, n10475, n10163, n12101, n12108,
    n9561, n15848, n15847, n10965, n10159, n10078, n13294, n11329, n12084,
    n13003, n15724, n16606, n16405, n12303, n11225, n16393, n16367, n16265,
    n16853, n9476, n16135, n10376, n9450, n12646, n15030, n15031, n16248,
    n16609, n10830, n12106, n11977, n10882, n13988, n16338, n15869, n16054,
    n12083, n12302, n16379, n15913, n10657, n14642, n16164, n15557, n11971,
    n11975, n16160, n11788, n11278, n10963, n12091, n11965, n16209, n16816,
    n10156, n12334, n10956, n16347, n15452, n16511, n11313, n16516, n11262,
    n9473, n17126, n10623, n10829, n11170, n11104, n10678, n16787, n11260,
    n10728, n10598, n11122, n11196, n11312, n12090, n11964, n11157, n10252,
    n15689, n13443, n10345, n15762, n10483, n11751, n10073, n11762, n10466,
    n16087, n10544, n11748, n11758, n16781, n15509, n9379, n15758, n12002,
    n13020, n10250, n10676, n11103, n11156, n11169, n11277, n11311, n16452,
    n15967, n10727, n17147, n9990, n15578, n10253, n11745, n10828, n9350,
    n11755, n11195, n10525, n10508, n13317, n11270, n12009, n12005, n15745,
    n15725, n11954, n10751, n9208, n12539, n12120, n11259, n16544, n10287,
    n11719, n11714, n9309, n10474, n10553, n10569, n10536, n10070, n9040,
    n10589, n11814, n14906, n9274, n10147, n10315, n15512, n10497, n13366,
    n11686, n10034, n10616, n10720, n10235, n16534, n10455, n10430, n15806,
    n10409, n15801, n16713, n10826, n15360, n11190, n13818, n16739, n15088,
    n10764, n10644, n15789, n15258, n12181, n16837, n11294, n10008, n10040,
    n9849, n15335, n10002, n9978, n11255, n9818, n9588, n13474, n9960,
    n15372, n11248, n9876, n11097, n13228, n9339, n15451, n9929, n11733,
    n11150, n11144, n17062, n11318, n9890, n11163, n11167, n11154, n15832,
    n9972, n9202, n10824, n14825, n11373, n10765, n15404, n10120, n16474,
    n15713, n11119, n9954, n12855, n10887, n9290, n10642, n9616, n9749,
    n9660, n11544, n9712, n10721, n11101, n10774, n11364, n9449, n15766,
    n9217, n9342, n9538, n9699, n9842, n12934, n9737, n9776, n9649, n11967,
    n9578, n10550, n9485, n10822, n9923, n10225, n9285, n12088, n10761,
    n10050, n9037, n9899, n15594, n11417, n10217, n10549, n9884, n10675,
    n9952, n11436, n17091, n14876, n9870, n15595, n10760, n9038, n11369,
    n10715, n10620, n9521, n10470, n11365, n13968, n14099, n15793, n15791,
    n11671, n10175, n9844, n10114, n10638, n10450, n10220, n11944, n9520,
    n14038, n16967, n11378, n16847, n10593, n9266, n13461, n9128, n10533,
    n17092, n10557, n10042, n10113, n9597, n9671, n9594, n11046, n12135,
    n10449, n9438, n9805, n9812, n9726, n10227, n9632, n10538, n10634,
    n9232, n10491, n9407, n9596, n9562, n11532, n9517, n11363, n11846,
    n10045, n9569, n9861, n9980, n11935, n9570, n9400, n9440, n9524, n9532,
    n9892, n9368, n9864, n11033, n9482, n10061, n9762, n9680, n9704, n9772,
    n10131, n11042, n11043, n9830, n9635, n9796, n9863, n9284, n9945,
    n9634, n9289, n9640, n9530, n9399, n9367, n9568, n9894, n9231, n9405,
    n9764, n11067, n9798, n9265, n9652, n14388, n10129, n9186, n9832,
    n9694, n9080, n10066, n9566, n9283, n14582, n11038, n10564, n9835,
    n10718, n11059, n9801, n10126, n10018, n10499, n9077, n9479, n9866,
    n9600, n10404, n9602, n9288, n9230, n14577, n9638, n9494, n9684, n9099,
    n9188, n9491, n10436, n10432, n9097, n9421, n9034, n10189, n9096,
    n10385, n9113, n9418, n10398, n10179, n10188, n9318, n10203, n10193,
    n10128, n9079, n9089, n9124, n10365, n9056, n10207, n10226, n9683,
    n9111, n9109, n9703, n9123, n9733, n10606, n10608, n9063, n9643, n9060,
    n10182, n10181, n9061, n9639, n10210, n10247, n10201, n10202, n10192,
    n10127, n10197, n10810, n9119, n10015, n10249, n9651, n10403, n9101,
    n10019, n10629, n10485, n9300, n10198, n10635, n15858, n15857, n15785,
    n15788, n15667, n15670, n16479, n15503, n15731, n15719, n15822, n15500,
    n16851, n15665, n15826, n15773, n15497, n15680, n10033, n15487, n17075,
    n15472, n15683, n15491, n17033, n15790, n17078, n15562, n11250, n15629,
    n15632, n15607, n16963, n16844, n15460, n15457, n16434, n16032, n15676,
    n15113, n15362, n15224, n15626, n15130, n15718, n16825, n15363, n15361,
    n15381, n15455, n15717, n15060, n15454, n15616, n16959, n15625, n15604,
    n15121, n15748, n15039, n16807, n15505, n15269, n17028, n16955, n15352,
    n16426, n15384, n15427, n15267, n15353, n17066, n15047, n16786, n15211,
    n16422, n15426, n15385, n15383, n15311, n17027, n15605, n11131, n15169,
    n15484, n15770, n16025, n15328, n16804, n16432, n16827, n17035, n17125,
    n15343, n15406, n15191, n15599, n16023, n15327, n17148, n15003, n9938,
    n15190, n15342, n11138, n15166, n15854, n17059, n15652, n15768, n15761,
    n11341, n17116, n15852, n9910, n17022, n11321, n15650, n15247, n16862,
    n16413, n15825, n16024, n11202, n15727, n15794, n15729, n16950, n17102,
    n15673, n14779, n15778, n15246, n15309, n15846, n17106, n14818, n16860,
    n9883, n17021, n17114, n17119, n14589, n14712, n14581, n14990, n14815,
    n14905, n15412, n17118, n16527, n14408, n15411, n16946, n15647, n14787,
    n11308, n11324, n14941, n14413, n16021, n10080, n10737, n10082, n15622,
    n17054, n17056, n15568, n15660, n10169, n16945, n16439, n14729, n14928,
    n14707, n10079, n14976, n10735, n15417, n14763, n15575, n15707, n15816,
    n14979, n10057, n15723, n10054, n15067, n16856, n15684, n15423, n15945,
    n15828, n16019, n15600, n16810, n14202, n10052, n15409, n14467, n15602,
    n10055, n15609, n14751, n15493, n14650, n11290, n16398, n15296, n16863,
    n16788, n15940, n14698, n14934, n15177, n16376, n11285, n9999, n14387,
    n16383, n10028, n10996, n10031, n14738, n15314, n14214, n16764, n16868,
    n14686, n16874, n10029, n10026, n15402, n15539, n14520, n14211, n14042,
    n15287, n16385, n16370, n14098, n11181, n9991, n14757, n9996, n16782,
    n14128, n15935, n15337, n14125, n15173, n16929, n15100, n14613, n15468,
    n14115, n16870, n15172, n9992, n15306, n9989, n15445, n14112, n15581,
    n15276, n14657, n11176, n14676, n16355, n14445, n14093, n15506, n13946,
    n14986, n10986, n15516, n9964, n15171, n14983, n15579, n14077, n14489,
    n13940, n11030, n16341, n16366, n14023, n14290, n14020, n14293, n14503,
    n9970, n11004, n15929, n15119, n9939, n9963, n14494, n13920, n9933,
    n14370, n13923, n14380, n15928, n14744, n14291, n11177, n13808, n13752,
    n16353, n14383, n10858, n15052, n14310, n14399, n14067, n15081, n16866,
    n16736, n14402, n16745, n15044, n9932, n14978, n15018, n15114, n14061,
    n16350, n14717, n15924, n13897, n14060, n14306, n11148, n10953, n13900,
    n14162, n16735, n15092, n14303, n13705, n15080, n13710, n16333, n14368,
    n14035, n11135, n14176, n14376, n16008, n16744, n9901, n14257, n9904,
    n15922, n16867, n16547, n14716, n15043, n14032, n16734, n14073, n17010,
    n14810, n14846, n14811, n15919, n9907, n15920, n14998, n15917, n11223,
    n13916, n14766, n14300, n16535, n13906, n14690, n14952, n14142, n9879,
    n13732, n13986, n9882, n16875, n10734, n14749, n16549, n14601, n14230,
    n13728, n11111, n16720, n14248, n14704, n11092, n13812, n14599, n16723,
    n16543, n16530, n14684, n9855, n9852, n16721, n14396, n9791, n11134,
    n16711, n13957, n13746, n13731, n15909, n9790, n14482, n10236, n15906,
    n10992, n9824, n9787, n9821, n14606, n16706, n15904, n15883, n11208,
    n10600, n13627, n9756, n13600, n13700, n13787, n13448, n15907, n14347,
    n13690, n14875, n16001, n14284, n9751, n9755, n14051, n15997, n16280,
    n11015, n14562, n10863, n13442, n11013, n17000, n16257, n14070, n15891,
    n14868, n16677, n11010, n14426, n16659, n9797, n15996, n9667, n11014,
    n9714, n14557, n13869, n13994, n9718, n16260, n14416, n10394, n10972,
    n14068, n10545, n10974, n9622, n16645, n13878, n10554, n14148, n16672,
    n9662, n16996, n10663, n13864, n9727, n9618, n16994, n13770, n13873,
    n13911, n10517, n9508, n13197, n13637, n16198, n16989, n12921, n13531,
    n15553, n9555, n13102, n16624, n9507, n9468, n10498, n12869, n12836,
    n13599, n16935, n12914, n13738, n16915, n9550, n15894, n9467, n12573,
    n14448, n12694, n16427, n13837, n16985, n9363, n16983, n15736, n16151,
    n14078, n15977, n11330, n14079, n15861, n17131, n11201, n15971, n15482,
    n9362, n12321, n9354, n15976, n16148, n11130, n16146, n10431, n12873,
    n9393, n9389, n9360, n17128, n16514, n13184, n16510, n15532, n16132,
    n16110, n12994, n16226, n14796, n16244, n14506, n16277, n16192, n14167,
    n10077, n15849, n16051, n13642, n13424, n10894, n13288, n12140, n15765,
    n12779, n10526, n10153, n15313, n9327, n10509, n12502, n12501, n10444,
    n10410, n12876, n10877, n12007, n9511, n16979, n10155, n15696, n10679,
    n12819, n17041, n16115, n10152, n10726, n11464, n11664, n15800, n15804,
    n11646, n10766, n10465, n12687, n10484, n9240, n11105, n11102, n10516,
    n11123, n10673, n10288, n11168, n11155, n11120, n10588, n10568, n13783,
    n13855, n14605, n10723, n11635, n11307, n13121, n16568, n10749, n10300,
    n10234, n16666, n16678, n14527, n16717, n9369, n10123, n11611, n13104,
    n10615, n16693, n10717, n10880, n10722, n12157, n10233, n10552, n9132,
    n10614, n12794, n9036, n10724, n10122, n15407, n12668, n11372, n10714,
    n9172, n11007, n15549, n12153, n16492, n14833, n10719, n9147, n9921,
    n9194, n10137, n10471, n9868, n15203, n12311, n9987, n16471, n14655,
    n10024, n11368, n14424, n16478, n10223, n10548, n10115, n10215, n10141,
    n15619, n11303, n9672, n10513, n9682, n10212, n17084, n9518, n9560,
    n10532, n16843, n14836, n10637, n10111, n9950, n9646, n9642, n10208,
    n9837, n9803, n9730, n10022, n9741, n9083, n10010, n10486, n9943,
    n9086, n9631, n11036, n10211, n9681, n9512, n9519, n11423, n9913,
    n9127, n10064, n9120, n9228, n9125, n9514, n9523, n9185, n10519, n9103,
    n9262, n10426, n11049, n9644, n14094, n9090, n9371, n9918, n9948,
    n9442, n10017, n9153, n9676, n9677, n9985, n9292, n9122, n9528, n9897,
    n9475, n9584, n9728, n10047, n9264, n9403, n9767, n9637, n9100, n9267,
    n9867, n9527, n9402, n9729, n10048, n11090, n9534, n9565, n9898,
    n14962, n9768, n9291, n9986, n9286, n10480, n9599, n9802, n9836, n9919,
    n9233, n10067, n9370, n9474, n9949, n9441, n9234, n9152, n10124, n9287,
    n9268, n10190, n10204, n10200, n10289, n9046, n9062, n9053, n10180,
    n9057, n10183, n9164, n9163, n10214, n10312, n9085, n9050, n10565,
    n10270, n12666, n14583, n10310, n16969, n9039, n17104, n11061, n17110,
    n9934, n9072, n12014, n16080, n12388, n12346, n16070, n10016, n13250,
    n9857, n9851, n9995, n15214, n9183, n16006, n14147, n10918, n10950,
    n10941, n15829, n9531, n13204, n11267, n10245, n15461, n10587, n10393,
    n9750, n9994, n9826, n9820, n9752, n9601, n9774, n11245, n10476,
    n10567, n10551, n10535, n10375, n12006, n9965, n9859, n12046, n16079,
    n16273, n16061, n16729, n16450, n15709, n11159, n15104, n10628, n16143,
    n10276, n9174, n9770, n9121, n9689, n9515, n9526, n9513, n11298,
    n10904, n11239, n11244, n10901, n13556, n11213, n10555, n10539, n10540,
    n11804, n13865, n10299, n10886, n15371, n15492, n15278, n11116, n10672,
    n10998, n12993, n10490, n9661, n9967, n9962, n10081, n9878, n9881,
    n10032, n10027, n10030, n9786, n9993, n9931, n9553, n10058, n10053,
    n10056, n9314, n9137, n11759, n14591, n12451, n15635, n16531, n14215,
    n13587, n13583, n9237, n10014, n9896, n9763, n9678, n9563, n9471,
    n10383, n11323, n11320, n10439, n10440, n11228, n15010, n11254, n11252,
    n11264, n11265, n14433, n16285, n11193, n11166, n11153, n11118, n11100,
    n10677, n10251, n10242, n10622, n10621, n10619, n10597, n10596, n10592,
    n10573, n12307, n13875, n14567, n14881, n15051, n14701, n14102, n10473,
    n13696, n13740, n10362, n16038, n10281, n14703, n14116, n14119, n14083,
    n14014, n13399, n10531, n10547, n9902, n9905, n14146, n10000, n9758,
    n9810, n9808, n9848, n12041, n11675, n9614, n9071, n9612, n9215, n9214,
    n9144, n9143, n9074, n9075, n9069, n11691, n14834, n15198, n9605,
    n9603, n15743, n14277, n14371, n14294, n14391, n13657, n13407, n13342,
    n13166, n13425, n17073, n9773, n14627, n9481, n9446, n10477, n14895,
    n11025, n11024, n15439, n10515, n13653, n13650, n13017, n14425, n13886,
    n13734, n13715, n13496, n14850, n14849, n14860, n14859, n13861, n14826,
    n14823, n14693, n14680, n14852, n14502, n14318, n9082, n16091, n16106,
    n16102, n16145, n16194, n16206, n16219, n16217, n16238, n16627, n16259,
    n16275, n16656, n16648, n16673, n16684, n16698, n16312, n16709, n16708,
    n16705, n16707, n16696, n16697, n16329, n16731, n16726, n16727, n16545,
    n15901, n15897, n15893, n16356, n16354, n16372, n16749, n16748, n16746,
    n16759, n16752, n16758, n16757, n16756, n15915, n15912, n15910, n16387,
    n16374, n16399, n16770, n16767, n16765, n16796, n16523, n15931, n15925,
    n16415, n17046, n16813, n16429, n16442, n16873, n16872, n16859, n16819,
    n16817, n16818, n16815, n16820, n16811, n16812, n16785, n16803, n17013,
    n15941, n15918, n15899, n17055, n17053, n17052, n17049, n16829, n16949,
    n17005, n9055, n9516, n10935, n10395, n10923, n10947, n10928, n16026,
    n16028, n16453, n16251, n10297, n16410, n11188, n11084, n10667, n16062,
    n16063, n16243, n13689, n16165, n16166, n16150, n10186, n10187, n17065,
    n16841, n17029, n9571, n9533, n16628, n9408, n9775, n14133, n16892,
    n10787, n12373, n9094, n9098, n9725, n9404, n10382, n10494, n11019,
    n11218, n11229, n10944, n10897, n13021, n10521, n10522, n10523, n10504,
    n10505, n10506, n10461, n10462, n10464, n12064, n11934, n12582, n12586,
    n12920, n13536, n10957, n11327, n15466, n15467, n14566, n10534, n10472,
    n10656, n10364, n10355, n15833, n15708, n15777, n15712, n15710, n15544,
    n15550, n15548, n15552, n15270, n15271, n11189, n15105, n15029, n11106,
    n11107, n14771, n14702, n10729, n10626, n10625, n10852, n14054, n14005,
    n13983, n13908, n13730, n10419, n10652, n10649, n12900, n10218, n10447,
    n10396, n17135, n9430, n15690, n9465, n9628, n12774, n9356, n11683,
    n11696, n11724, n13462, n13761, n14336, n14827, n14236, n11981, n9604,
    n11524, n9372, n9315, n15163, n15593, n15393, n15300, n15170, n15155,
    n14969, n14909, n14732, n14670, n14593, n14471, n14349, n14150, n14229,
    n13965, n13782, n13596, n13592, n13792, n9293, n9332, n10021, n9984,
    n9641, n9673, n9636, n9567, n9559, n9525, n9529, n9445, n9439, n9397,
    n9365, n9330, n9154, n9110, n15138, n10481, n10482, n10478, n12406,
    n14638, n11300, n11299, n13297, n12325, n16076, n14891, n15524, n10514,
    n14256, n10479, n12415, n11209, n11215, n11216, n16392, n11314, n11274,
    n11276, n15564, n11261, n11192, n10561, n10560, n10543, n10324, n10254,
    n11803, n12129, n12123, n12913, n13530, n11662, n16501, n15776, n15824,
    n15659, n15473, n15478, n15125, n16337, n14996, n14809, n10732, n14458,
    n10841, n14117, n14012, n14011, n13932, n13890, n13438, n10641, n15547,
    n12008, n16500, n15775, n15658, n15336, n15027, n14808, n14459, n14457,
    n14204, n10846, n10845, n14203, n15657, n14072, n13893, n13892, n13619,
    n13620, n13628, n13626, n13743, n13495, n13397, n14993, n10883, n12021,
    n14961, n10238, n16487, n10191, n10636, n10493, n10271, n11487, n9361,
    n12749, n12748, n16524, n9243, n9856, n17111, n12822, n16689, n9793,
    n9794, n9997, n12663, n13274, n9624, n9625, n13594, n13961, n9554,
    n9557, n10861, n10136, n12780, n12781, n15809, n17079, n10039, n10007,
    n9977, n9959, n9928, n9889, n9875, n9817, n9252, n9198, n11516, n11512,
    n14333, n13452, n13455, n13773, n14325, n15764, n17127, n15621, n15610,
    n15812, n15323, n15691, n15585, n15510, n14977, n14925, n14930, n15231,
    n15230, n14753, n14688, n14495, n16728, n14311, n16712, n16687, n14217,
    n15671, n15639, n15620, n15421, n15322, n15068, n14931, n14754, n14689,
    n14656, n14478, n15185, n13601, n13358, n13160, n9116, n12180, n12182,
    n15254, n14574, n11306, n11845, n10065, n10119, n14095, n10049, n9084,
    n13943, n9078, n9081, n13508, n17037, n9104, n11096, n9865, n17072,
    n13065, n12842, n12680, n14328, n12427, n12295, n12146, n12077, n9572,
    n11995, n11822, n11831, n11721, n11778, n11693, n9410, n11739, n11626,
    n11537, n11474, n9281, n10417, n10418, n10952, n15142, n15141, n15139,
    n13524, n14639, n14647, n10443, n14894, n14892, n14900, n15529, n15528,
    n15525, n14444, n14442, n15438, n13561, n14780, n14719, n14724, n10964,
    n15040, n15013, n15011, n10268, n14505, n14519, n14517, n15527, n10884,
    n11269, n15530, n10881, n10981, n11263, n11257, n11194, n11171, n11165,
    n11158, n11152, n11117, n11099, n10674, n10243, n10624, n10618, n10599,
    n10591, n10575, n10576, n16230, n16189, n16195, n16177, n10390, n10391,
    n10373, n10374, n10344, n16116, n10308, n10306, n12273, n12070, n13543,
    n14422, n14421, n14569, n14561, n14873, n15450, n15382, n11180, n11136,
    n14784, n14640, n10850, n14091, n14086, n13931, n13702, n13176, n13147,
    n14708, n14120, n14018, n14015, n13915, n13011, n12020, n11612, n13947,
    n13806, n12681, n13874, n13535, n12919, n12581, n12306, n11962, n10133,
    n14186, n15508, n13486, n12731, n17146, n17150, n16629, n15085, n15084,
    n15082, n15688, n14526, n14543, n14541, n15577, n14947, n14946, n15582,
    n15229, n14795, n14794, n14804, n16777, n15811, n14136, n10866, n10864,
    n9850, n9615, n9323, n9346, n9347, n12495, n9218, n9142, n9076, n14340,
    n14625, n14623, n15359, n15350, n14975, n14936, n14920, n14758, n14743,
    n14927, n13971, n13834, n15218, n10763, n15805, n14278, n14375, n14299,
    n14395, n13247, n13169, n13383, n12745, n11074, n11060, n14409, n14385,
    n13938, n13155, n14828, n9807, n13774, n13458, n12983, n12477, n9574,
    n12105, n11974, n9480, n11614, n11469, n11480, n11486, n9161, n11361,
    n10820, n11345, n11032, n13656, n13889, n14050, n14007, n13735, n13635,
    n13269, n13681, n13750, n13498, n13678, n13747, n13501, n14862, n13862,
    n14681, n14664, n14500, n14319, n14316, n14241, n13608, n13668, n13800,
    n13665, n13803, n13757, n9170, n10888, n9041, n16391, n16461, n9042,
    n16071, n9043, n16082, n16147, n16212, n15889, n16306, n16375, n16390,
    n16822, n15954, n10931, n11926, n10892, n10397, n11093, n11692, n9443,
    n16660, n16616, n10503, n11175, n14104, n9394, n9912, n15751, n14151,
    n9406, n9254, n11243, n10248, n16199, n16701, n13371, n9827, n9701,
    n9779, n9488, n11494, n15646, n14984, n14924, n9800, n9564, n11632,
    n12418, n10367, n15103, n10240, n11562, n12986, n15205, n9065, n9761,
    n9595, n10221, n14096, n11475, n13598, n16161, n12671, n9189, n9045,
    n9224, n9302, n9047, n9409, n9049, n9048, n9051, n9052, n9054, n9095,
    n9058, n9059, n9107, n9105, n11079, n9064, n9066, n9067, n9070, n9068,
    n9544, n11054, n9073, n9656, n10130, n13753, n9088, n9087, n11416,
    n9573, n9126, n9091, n9102, n9118, n9133, n9108, n9114, n9115, n11357,
    n9117, n12282, n13503, n16962, n10791, n9271, n9131, n9129, n9130,
    n11844, n9134, n17107, n9140, n12281, n14237, n9136, n9135, n11843,
    n9139, n9178, n9141, n9145, n9146, n12629, n9148, n9149, n9150, n9151,
    n9155, n9156, n9160, n9157, n9158, n9159, n9184, n9162, n9166, n9165,
    n9167, n11424, n9168, n9171, n12542, n17109, n9173, n9175, n12550,
    n9935, n9177, n9176, n9182, n9181, n12538, n10746, n9229, n9187,
    n11545, n9192, n9190, n11859, n9191, n9195, n9839, n9193, n12559,
    n16561, n9204, n9196, n9197, n9200, n9199, n9201, n12721, n9203,
    n16562, n9207, n9206, n10745, n9211, n9210, n12730, n9212, n9213,
    n9216, n9239, n9219, n9227, n9220, n9221, n9223, n9222, n9225, n9257,
    n11428, n9226, n9263, n11386, n9235, n9236, n12720, n9238, n9244,
    n9242, n16567, n9241, n9246, n9245, n12664, n9248, n9957, n9247,
    n12791, n9250, n9249, n9251, n12825, n9273, n11395, n9261, n9253,
    n9256, n9255, n9259, n9334, n9258, n11452, n9260, n9270, n9282, n9269,
    n9272, n9277, n9276, n9275, n9278, n9279, n9280, n12776, n9331, n9366,
    n9294, n9307, n9295, n9296, n9298, n9299, n9297, n9305, n9301, n9303,
    n9374, n9306, n9308, n13114, n9326, n9310, n9313, n9311, n9312, n9324,
    n9322, n9317, n9316, n9319, n12767, n9320, n9321, n16595, n9325, n9357,
    n9329, n9328, n9333, n9337, n9335, n9336, n9338, n12435, n9349, n9340,
    n9341, n9343, n12818, n9345, n9344, n12763, n9348, n12775, n9352,
    n9351, n9353, n9364, n9355, n9359, n9358, n12751, n9398, n9373, n9377,
    n9375, n9376, n9378, n13364, n9388, n9382, n9380, n9381, n9386, n13420,
    n9384, n9383, n9385, n9387, n9392, n9391, n9390, n9396, n9395, n9433,
    n9401, n9414, n9412, n9411, n9413, n13223, n9429, n9417, n9415, n9416,
    n9427, n9425, n9420, n9419, n9422, n13130, n9423, n9424, n9426, n9428,
    n9434, n12955, n9432, n9431, n12957, n9437, n9436, n9435, n12956,
    n13273, n9464, n9472, n9448, n9444, n9447, n13280, n9460, n13285,
    n9451, n9454, n9452, n9453, n9458, n9456, n9455, n9457, n9459, n9463,
    n9462, n9470, n9506, n9477, n9484, n9478, n9483, n13611, n9502, n9487,
    n9490, n9489, n9500, n9498, n9493, n9492, n9495, n13473, n9496, n9497,
    n9499, n9501, n13484, n9505, n9504, n9510, n9509, n13483, n13568,
    n9522, n9537, n9535, n9536, n9540, n9543, n9541, n9542, n9548, n9546,
    n13842, n9545, n9547, n9549, n9552, n9558, n9577, n9686, n9575, n9576,
    n13973, n9590, n9580, n9583, n9581, n9582, n9586, n13811, n9585, n9587,
    n9589, n9593, n9592, n9598, n16668, n9607, n13979, n9608, n9611, n9609,
    n9610, n9613, n9617, n9621, n9620, n13852, n9674, n9648, n9645, n9647,
    n16657, n14218, n9655, n9653, n9654, n9658, n9657, n9659, n14182,
    n9665, n9664, n9670, n9669, n14183, n10865, n9716, n9675, n9679, n9723,
    n9698, n9685, n9687, n9688, n9690, n9693, n9691, n9692, n9696, n9695,
    n9697, n14296, n9702, n10867, n9705, n9740, n9708, n9706, n9707, n9710,
    n9709, n9711, n9713, n9719, n9717, n9722, n9721, n9732, n9736, n9734,
    n9735, n16692, n9739, n9742, n14536, n9745, n9743, n9744, n9747, n9746,
    n9748, n9754, n9760, n14542, n9766, n9765, n9769, n9777, n9771, n9804,
    n16716, n9778, n9781, n9780, n9785, n14544, n9783, n9782, n9784, n9789,
    n9795, n9825, n9799, n9811, n9806, n9809, n14797, n9819, n9814, n9813,
    n9815, n9816, n14790, n9823, n9829, n9828, n14791, n14848, n9833,
    n9862, n9843, n9838, n9841, n9840, n16548, n9846, n9845, n14659, n9847,
    n9854, n9860, n15077, n9869, n9877, n9872, n9871, n9873, n9874, n9891,
    n9886, n9885, n9887, n9888, n9895, n9914, n9900, n9917, n9916, n9944,
    n9922, n9930, n9925, n9924, n9926, n9927, n15225, n9936, n9942, n9941,
    n15226, n9966, n9946, n9981, n9982, n9953, n9961, n9956, n9955, n14974,
    n9958, n15159, n15504, n9969, n9971, n15576, n9979, n9974, n9973,
    n9975, n9976, n15697, n9983, n10012, n9988, n10001, n15687, n10009,
    n10004, n10003, n10005, n10006, n10013, n10043, n10020, n10044, n10025,
    n15810, n10041, n10036, n10035, n10037, n10038, n10046, n10063, n10051,
    n10060, n17103, n11035, n10069, n10068, n10071, n10072, n10075, n10074,
    n10076, n10084, n10083, n10088, n10086, n10085, n10087, n10110, n10090,
    n10089, n10091, n10108, n10093, n10092, n10097, n10095, n10094, n10096,
    n10105, n10099, n10098, n10103, n10101, n10100, n10102, n10104, n10106,
    n10107, n10109, n10116, n10112, n10117, n12154, n10118, n12158, n10121,
    n10125, n17086, n10174, n17089, n15422, n10222, n10132, n10173, n10134,
    n17136, n10171, n10135, n12156, n10140, n10138, n10139, n10146, n10144,
    n10142, n13152, n10143, n10145, n17130, n15086, n10167, n10150, n15636,
    n10148, n10149, n17132, n10154, n10151, n10157, n10158, n10161, n10160,
    n10162, n17112, n10165, n10164, n10166, n10168, n10177, n10176, n10178,
    n10349, n10184, n10185, n10311, n10326, n10350, n10196, n10199, n10194,
    n10195, n10232, n10205, n10206, n10229, n10716, n10213, n10219, n10216,
    n10725, n13709, n10228, n14404, n10230, n10231, n10579, n10605, n10611,
    n16472, n10241, n10244, n14576, n10412, n10246, n10255, n10259, n10257,
    n10258, n12383, n16081, n10260, n10742, n10263, n10262, n10645, n12345,
    n10280, n10265, n10264, n10269, n10267, n10266, n10273, n10272, n10274,
    n11653, n10275, n10277, n12351, n10279, n10282, n16090, n12596, n10284,
    n10283, n10286, n10285, n16073, n10290, n10293, n10291, n10292, n10295,
    n10294, n11655, n12236, n10296, n10298, n13050, n16093, n10301, n10302,
    n16104, n12888, n10305, n10303, n10304, n10307, n10313, n11657, n10314,
    n10317, n10316, n13144, n12889, n10319, n16125, n10318, n12691, n10321,
    n10320, n10325, n10323, n12848, n10322, n12890, n11481, n10334, n10327,
    n10330, n10328, n10329, n10332, n10331, n11659, n10333, n10336, n10335,
    n12695, n10338, n10337, n12865, n10341, n10339, n13075, n10340, n10343,
    n10342, n13014, n10356, n10354, n10346, n10348, n10347, n10352, n10399,
    n10351, n10353, n13078, n16111, n16136, n15969, n12866, n10358, n10357,
    n10363, n10361, n10359, n10360, n13032, n10370, n10366, n13033, n10368,
    n10369, n10372, n10371, n13251, n10378, n10377, n10384, n10379, n10380,
    n10381, n13265, n10387, n13260, n10386, n10389, n10388, n15981, n13172,
    n10408, n10400, n10402, n10401, n10406, n10405, n10407, n10414, n13293,
    n10411, n10413, n10416, n10415, n16181, n10420, n13312, n10421, n10429,
    n10422, n10425, n10423, n10424, n10427, n10428, n16176, n10433, n10435,
    n10434, n10437, n10458, n13549, n10438, n10442, n10441, n16180, n10446,
    n10448, n10451, n10454, n10452, n10453, n16205, n10457, n10459, n13683,
    n10460, n10463, n10467, n10469, n13618, n16188, n13654, n10487, n10488,
    n10489, n10492, n10496, n10495, n16229, n10501, n10500, n10502, n14164,
    n10507, n10510, n10512, n13902, n14261, n10518, n10520, n14242, n13924,
    n10524, n10527, n10530, n10528, n13993, n16247, n13997, n10542, n10541,
    n10546, n14063, n16266, n10556, n10559, n14087, n10558, n10563, n10566,
    n10572, n14432, n10571, n10574, n10840, n10601, n10580, n10583, n10581,
    n10582, n10585, n10584, n16053, n13882, n10594, n10595, n10603, n15884,
    n16003, n10989, n10617, n10604, n10607, n10610, n10609, n10613, n10612,
    n16293, n16067, n11086, n10631, n10633, n16031, n10885, n10640, n10643,
    n14769, n16084, n12338, n10646, n12594, n10647, n10648, n12895, n10651,
    n10650, n12999, n10654, n13256, n10655, n13180, n10658, n15887, n10659,
    n13695, n15892, n10660, n13625, n13729, n13907, n13985, n14052, n10668,
    n10851, n10669, n10997, n10670, n11112, n16469, n10671, n16299, n11631,
    n10681, n16488, n10680, n10682, n10687, n10686, n10691, n10689, n10688,
    n10690, n10713, n10693, n10692, n10694, n10711, n10696, n10695, n10700,
    n10698, n10697, n10699, n10708, n10702, n10701, n10706, n10704, n10703,
    n10705, n10707, n10709, n10710, n10712, n10878, n16486, n16468, n14995,
    n12004, n15272, n15285, n10733, n13071, n10730, n12899, n10739, n10738,
    n10740, n10744, n10743, n10747, n10753, n12521, n10748, n10750, n12628,
    n10752, n10759, n10755, n10754, n10757, n10756, n10758, n10800, n10762,
    n16981, n16554, n16553, n16563, n16974, n12553, n10767, n10781, n16574,
    n16896, n16581, n17043, n16579, n16971, n10770, n12449, n16888, n16901,
    n12362, n16890, n16598, n13113, n10775, n10773, n13329, n15738, n10777,
    n10776, n10795, n12167, n10778, n10780, n10779, n12549, n10783, n10782,
    n12500, n16569, n10784, n12456, n16972, n10786, n10785, n16590, n10788,
    n16589, n13100, n12738, n10789, n10790, n10793, n10792, n10794, n12739,
    n12789, n13107, n10797, n10798, n10799, n10802, n10801, n10809, n15174,
    n12560, n12506, n12505, n10803, n10804, n13365, n12370, n16596, n10805,
    n12735, n10807, n10806, n10808, n10839, n10837, n13386, n13195, n12834,
    n12571, n12319, n12138, n12000, n11812, n10827, n10825, n10823, n10821,
    n11379, n10819, n10817, n10815, n11356, n10813, n11348, n11351, n11350,
    n10811, n11354, n11353, n10812, n11355, n10814, n11360, n10816, n11362,
    n10818, n11435, n11543, n11732, n11813, n12001, n12139, n12320, n12572,
    n12835, n13196, n13387, n13547, n10836, n10838, n10843, n10842, n10848,
    n14205, n10847, n10854, n10853, n10855, n10857, n14853, n10876, n10872,
    n10868, n13465, n10870, n10869, n10871, n10873, n10960, n10879, n10954,
    n16039, n10975, n10890, n12386, n10889, n12326, n12327, n10893, n12416,
    n10895, n12414, n10896, n10898, n12405, n10899, n10900, n10903, n10902,
    n10905, n12617, n12619, n10907, n10906, n10908, n10909, n10910, n12650,
    n12649, n10911, n10912, n10913, n10914, n10917, n10916, n10915, n10919,
    n10921, n10920, n10924, n10927, n10926, n10925, n10929, n10930, n13520,
    n10936, n10939, n10937, n13648, n10942, n10945, n10943, n10946, n14170,
    n10949, n10951, n10955, n15535, n10958, n12926, n10962, n10959, n15872,
    n10961, n10967, n10966, n10968, n10971, n10970, n10988, n10979, n10976,
    n14436, n14434, n11017, n10982, n13529, n10984, n10983, n10985, n10991,
    n10990, n10994, n10993, n11000, n10999, n11001, n11003, n11009, n11008,
    n14437, n11023, n11018, n11205, n11026, n14415, n11028, n11027, n11029,
    n11039, n11041, n11040, n11045, n11302, n11048, n11047, n11051, n11050,
    n11053, n11052, n14384, n11056, n14585, n11055, n11057, n11063, n11062,
    n11064, n11070, n11069, n11072, n11071, n11073, n11076, n11077, n11078,
    n11081, n11080, n11082, n11088, n14768, n11095, n11109, n11108, n13335,
    n16322, n11142, n11110, n14994, n16294, n14770, n15916, n11114, n11185,
    n11125, n16334, n11124, n11126, n11133, n11132, n15025, n11143, n15926,
    n16012, n15024, n15101, n11151, n11149, n16014, n15099, n11172, n11162,
    n16363, n16016, n11173, n15242, n11178, n15244, n11179, n11186, n15028,
    n11187, n15275, n11198, n15463, n11197, n11199, n11206, n11210, n11211,
    n14518, n11214, n14637, n11219, n14718, n11224, n14893, n14890, n11230,
    n11231, n15012, n11233, n15009, n11237, n11235, n15140, n15137, n11242,
    n11240, n11241, n15436, n11247, n11246, n15435, n15526, n11249, n13944,
    n15523, n11253, n11291, n11256, n11258, n11266, n11289, n11279, n11272,
    n11271, n11273, n11275, n15704, n11287, n11283, n11281, n11280, n11282,
    n11284, n11293, n15860, n11297, n11295, n14198, n15863, n15202, n11310,
    n11309, n11317, n15868, n11319, n11343, n11339, n11337, n11335, n11326,
    n11325, n11331, n11328, n11333, n11332, n11334, n11336, n11347, n11346,
    n11349, n11352, n11359, n11358, n11367, n11366, n11371, n11370, n11375,
    n11374, n11377, n11376, n11381, n11380, n11383, n11382, n11385, n11384,
    n11388, n11387, n11390, n11389, n11392, n11391, n11394, n11393, n11399,
    n11397, n11396, n11398, n11403, n11401, n11584, n11400, n11402, n11405,
    n11404, n11407, n11406, n12726, n11570, n11569, n11572, n11408, n11852,
    n11851, n11853, n11409, n11413, n11412, n11411, n14411, n11410, n11414,
    n11444, n11415, n11421, n17096, n14842, n11419, n14386, n11422, n14837,
    n11449, n11418, n11420, n11434, n11492, n11836, n11838, n11576, n11578,
    n11425, n11857, n11856, n11427, n11426, n11431, n11430, n11429, n11432,
    n11451, n11433, n11463, n11438, n11437, n11440, n11439, n11442, n11441,
    n12766, n11443, n11911, n11910, n11912, n11907, n11445, n11556, n11555,
    n11557, n11446, n11515, n11447, n11448, n11460, n11450, n11905, n11904,
    n11454, n11453, n11551, n11550, n11552, n11455, n11508, n11507, n11456,
    n11458, n11517, n11457, n11459, n11462, n11461, n11466, n11465, n11468,
    n11467, n11471, n11470, n11473, n11472, n11477, n11476, n11479, n11478,
    n11485, n11483, n11482, n11484, n11491, n11489, n11488, n11490, n11496,
    n11493, n11495, n11497, n11501, n11499, n11498, n11500, n11506, n11503,
    n11502, n11504, n11505, n11510, n11509, n11511, n11514, n11513, n11529,
    n11519, n11518, n11521, n11520, n11523, n11522, n11525, n12755, n11527,
    n11689, n11526, n11528, n11531, n11530, n11534, n11533, n11536, n11535,
    n11540, n11538, n11539, n11542, n11541, n11547, n11546, n11549, n11548,
    n11554, n11553, n11566, n11559, n11558, n11561, n11560, n12826, n11564,
    n11563, n11565, n11568, n11567, n11571, n11573, n11575, n11574, n11583,
    n11581, n11577, n11579, n11580, n11582, n11586, n11585, n11588, n11587,
    n11590, n11589, n11592, n11591, n11594, n11593, n11596, n11595, n11598,
    n11597, n11600, n11599, n11602, n11601, n11604, n11603, n11606, n11605,
    n11608, n11607, n11610, n11609, n11616, n11615, n11618, n11617, n11625,
    n11620, n11619, n11623, n11621, n11622, n11624, n11628, n11927, n11627,
    n11630, n11629, n12644, n11633, n11634, n14864, n11636, n11652, n12187,
    n12247, n12246, n12249, n12255, n11637, n12223, n12222, n12225, n11638,
    n12204, n12203, n12206, n12217, n11639, n12032, n12031, n11641, n12038,
    n11640, n11643, n11642, n11924, n11645, n11644, n11648, n11647, n11932,
    n11650, n14887, n11649, n11651, n11670, n12186, n12240, n12239, n12242,
    n11654, n12228, n12227, n12230, n11656, n12209, n12208, n12211, n11658,
    n12029, n12028, n11661, n11660, n11667, n11666, n11665, n15261, n11663,
    n14882, n12924, n11668, n11937, n11669, n11679, n11673, n11672, n11677,
    n11674, n11676, n11678, n11681, n11680, n12951, n11682, n11685, n11684,
    n11687, n11688, n11703, n11701, n11690, n11734, n11694, n11712, n11695,
    n11698, n11697, n11699, n11700, n11702, n11705, n11704, n11707, n11706,
    n11709, n11708, n11711, n11710, n11713, n11779, n11716, n11715, n11756,
    n11754, n11717, n11729, n11718, n11722, n11720, n11746, n11744, n11723,
    n11725, n13276, n11727, n11726, n11728, n11731, n11730, n11736, n11735,
    n11738, n11737, n11741, n11740, n11743, n11742, n13479, n11747, n11750,
    n11749, n11752, n11753, n11767, n11765, n11757, n11761, n11760, n11763,
    n11764, n11766, n11769, n11768, n11771, n11770, n11773, n11772, n11775,
    n11774, n11777, n11776, n11781, n11780, n11783, n11782, n11785, n11784,
    n11787, n11786, n11790, n11789, n11796, n11792, n11791, n11794, n11793,
    n11795, n11798, n11797, n11800, n11799, n11802, n11801, n11811, n11806,
    n11805, n11809, n11808, n11810, n11815, n11817, n11816, n11819, n11818,
    n11821, n11820, n11824, n11823, n11826, n11825, n11828, n11827, n11830,
    n11829, n11833, n11832, n11835, n11834, n11837, n11840, n11839, n11842,
    n11841, n11849, n12630, n17087, n11847, n11848, n11850, n11918, n11855,
    n11854, n11863, n11858, n11861, n11860, n11862, n11865, n11864, n11866,
    n11868, n11867, n11870, n11869, n11872, n11871, n11874, n11873, n11876,
    n11875, n11878, n11877, n11880, n11879, n11882, n11881, n11884, n11883,
    n11886, n11885, n11887, n11889, n11888, n11891, n11890, n11893, n11892,
    n11895, n11894, n11897, n11896, n11899, n11898, n11901, n11900, n11903,
    n11902, n11906, n11909, n11908, n11916, n11914, n11913, n11915, n11917,
    n12672, n11919, n11921, n11920, n13550, n11922, n11949, n11931, n12126,
    n11923, n12260, n12259, n12262, n11925, n12056, n11929, n11928, n12055,
    n12054, n11930, n12127, n11953, n11933, n11947, n11943, n12121, n11936,
    n12265, n12264, n12267, n11938, n12062, n11940, n11939, n11941, n12060,
    n11942, n11963, n11945, n11946, n11948, n11951, n11950, n13513, n11952,
    n11961, n11959, n11956, n11955, n12089, n11957, n11958, n11960, n11970,
    n11966, n12082, n11968, n11969, n12107, n11972, n11973, n11986, n11978,
    n11976, n11980, n11979, n11982, n13570, n11984, n11983, n11985, n11988,
    n11987, n11990, n11989, n11992, n11991, n11994, n11993, n11997, n11996,
    n11999, n11998, n12003, n12019, n12010, n15970, n12011, n12013, n12012,
    n13093, n13094, n16498, n12016, n12015, n12017, n12022, n12018, n12024,
    n12023, n12026, n12025, n12613, n12027, n12037, n12030, n12035, n12033,
    n12034, n12036, n12040, n12039, n12052, n12045, n12042, n12044, n12050,
    n12048, n12047, n12049, n12051, n13199, n12053, n12069, n12058, n12057,
    n12059, n12067, n12061, n12063, n12065, n12066, n12068, n12072, n12071,
    n12074, n12073, n12076, n12075, n12079, n12078, n12081, n12080, n13640,
    n12085, n12086, n12087, n12097, n12095, n12092, n12301, n12093, n12094,
    n12096, n12099, n12098, n13819, n12100, n12114, n12471, n12470, n12103,
    n12102, n12104, n12112, n12109, n12478, n12110, n12111, n12113, n12116,
    n12115, n12119, n12118, n13289, n12122, n12124, n12125, n12134, n12132,
    n12128, n12917, n12130, n12131, n12133, n12137, n12136, n12141, n12143,
    n12142, n12145, n12144, n12148, n12147, n12150, n12149, n12152, n12151,
    n12155, n12179, n16558, n12168, n12276, n12159, n12161, n12160, n12166,
    n12162, n12164, n12163, n12165, n12170, n12520, n12169, n12525, n12176,
    n12172, n12171, n12519, n12174, n12173, n12175, n12177, n12183, n12178,
    n12185, n12184, n12191, n12189, n12188, n12190, n12192, n12196, n12194,
    n12193, n12195, n12201, n12198, n12197, n12199, n12200, n12401, n12202,
    n12216, n12205, n12207, n12214, n12210, n12212, n12213, n12215, n12219,
    n12218, n12221, n12220, n12235, n12224, n12226, n12233, n12229, n12231,
    n12232, n12234, n12238, n12237, n12241, n12243, n12245, n12244, n12254,
    n12252, n12248, n12250, n12251, n12253, n12257, n12256, n13015, n12258,
    n12272, n12261, n12263, n12270, n12266, n12268, n12269, n12271, n12275,
    n12274, n12287, n16975, n12936, n12277, n12279, n12278, n12942, n12280,
    n12284, n12283, n12285, n12288, n12286, n12290, n12289, n12292, n12291,
    n12294, n12293, n12297, n13771, n12296, n12299, n12298, n14165, n12300,
    n12316, n12304, n12576, n12305, n12314, n12310, n12312, n12313, n12315,
    n12318, n12317, n12322, n12333, n12324, n12323, n12331, n12328, n12329,
    n12330, n12332, n12336, n12420, n12335, n12358, n15972, n12337, n12339,
    n12340, n12344, n12342, n12341, n12343, n12349, n12815, n12347, n12348,
    n12811, n12350, n12807, n12355, n12353, n12352, n12354, n12356, n12359,
    n12357, n12361, n12360, n12379, n12363, n12367, n12365, n12364, n12366,
    n12444, n12368, n12369, n12371, n12439, n12438, n14935, n12375, n12374,
    n12376, n12377, n12380, n12378, n12382, n12381, n12394, n12392, n12384,
    n12385, n12387, n12390, n12389, n12391, n12393, n12396, n12395, n12398,
    n12397, n12404, n12400, n12399, n12402, n12403, n12411, n12409, n12407,
    n12408, n12410, n12413, n12412, n12426, n12417, n12419, n12424, n12422,
    n12421, n12423, n12425, n12430, n12428, n12429, n12432, n12431, n12434,
    n12433, n12437, n12436, n12443, n12441, n12440, n12442, n12445, n12446,
    n12448, n12447, n12465, n12450, n12455, n12453, n12452, n12454, n12458,
    n12790, n12457, n12788, n12462, n12801, n12460, n12459, n12461, n12463,
    n12466, n12464, n12468, n12467, n12473, n12476, n12475, n12491, n12482,
    n12481, n12485, n12484, n12487, n12486, n13853, n12489, n12488, n12490,
    n12493, n12492, n12515, n12494, n12499, n12497, n12496, n12498, n12715,
    n12504, n12503, n12714, n12512, n12508, n12507, n12707, n12510, n12509,
    n12511, n12513, n12516, n12514, n12518, n12517, n12531, n12524, n12523,
    n12526, n12527, n12529, n12528, n12530, n12533, n12532, n12536, n12535,
    n12546, n12540, n12541, n12544, n12543, n12545, n12548, n12547, n12567,
    n12963, n12558, n12552, n12551, n12556, n12554, n12555, n12557, n12962,
    n12564, n12972, n12562, n12561, n12563, n12565, n12568, n12566, n12570,
    n12569, n12574, n14243, n12575, n12591, n12579, n12580, n12589, n12585,
    n12587, n12588, n12590, n12593, n12592, n12609, n15975, n12595, n12598,
    n13047, n12597, n12602, n12600, n12599, n12601, n13058, n13053, n12604,
    n12603, n12605, n12607, n12606, n12610, n12608, n12612, n12611, n12614,
    n12616, n12615, n12623, n12620, n12621, n12622, n12625, n12624, n12627,
    n12626, n12636, n12634, n12632, n12631, n12633, n12635, n12638, n12637,
    n12641, n12639, n12640, n12643, n12642, n12645, n12648, n12647, n12660,
    n12653, n12652, n12654, n12658, n12656, n12655, n12657, n12659, n12662,
    n12661, n12679, n12665, n12667, n12677, n12670, n12669, n12675, n12673,
    n12674, n12676, n12678, n12683, n12682, n12685, n12684, n12703, n12686,
    n12853, n12690, n12859, n12688, n12689, n12701, n12847, n12699, n12693,
    n12692, n12698, n12696, n12697, n12856, n12700, n12704, n12702, n12706,
    n12705, n12713, n12709, n12708, n12711, n12710, n12712, n12719, n13829,
    n12716, n12717, n12718, n12725, n12723, n12722, n12724, n12727, n12729,
    n12728, n12734, n12732, n12733, n12744, n12737, n12736, n12742, n12740,
    n12741, n12743, n12747, n12746, n12750, n12752, n12760, n12754, n12753,
    n12758, n12756, n12757, n12759, n12762, n12761, n12765, n12764, n12773,
    n12771, n12769, n12768, n12770, n12772, n12787, n12820, n12778, n12777,
    n12784, n12782, n12783, n12785, n12786, n12800, n15608, n12798, n12793,
    n12792, n12796, n12795, n12797, n12799, n12803, n12802, n12805, n12804,
    n12814, n12809, n12808, n12810, n12812, n12813, n12817, n12816, n12833,
    n12821, n12831, n12824, n12823, n12829, n12827, n12828, n12830, n12832,
    n12837, n12839, n12838, n12841, n12840, n12844, n12843, n12846, n12845,
    n12852, n12850, n12849, n12851, n12864, n12854, n12861, n12857, n12858,
    n12860, n12862, n12863, n12884, n13085, n12868, n12867, n12872, n12870,
    n12871, n13073, n12881, n12875, n12874, n13070, n12879, n13072, n12877,
    n12878, n12880, n12882, n12885, n12883, n12887, n12886, n12909, n13143,
    n12894, n12892, n12891, n12893, n12898, n12896, n12897, n13139, n12903,
    n12901, n12902, n13137, n12905, n12904, n12906, n12907, n12910, n12908,
    n12912, n12911, n12916, n12918, n12931, n12923, n12925, n12927, n12929,
    n12928, n12930, n12933, n12932, n12935, n12941, n12937, n12939, n12938,
    n12940, n12946, n12943, n12944, n12945, n12950, n12948, n12947, n12949,
    n12952, n12954, n12953, n12961, n12958, n12959, n12960, n12971, n12967,
    n12965, n12964, n12966, n12969, n12968, n12970, n12974, n12973, n14187,
    n12975, n12982, n12980, n12977, n12978, n12979, n12981, n12992, n12985,
    n12989, n12987, n12990, n12991, n13010, n13039, n12998, n12996, n12995,
    n12997, n13002, n13000, n13001, n13044, n13038, n13005, n13004, n13006,
    n13008, n13007, n13009, n13013, n13012, n13016, n13019, n13018, n13031,
    n13029, n13027, n13023, n13025, n13026, n13028, n13030, n13035, n13034,
    n13037, n13036, n13043, n13041, n13040, n13042, n13046, n13045, n13057,
    n13049, n13048, n13052, n13051, n13055, n13054, n13056, n13060, n13059,
    n13062, n13061, n13064, n13063, n13067, n13066, n13069, n13068, n13084,
    n13074, n13082, n13077, n13076, n13080, n13079, n13081, n13083, n13087,
    n13086, n13089, n13088, n13092, n13090, n13091, n13098, n13096, n13095,
    n13097, n16617, n13099, n13101, n13370, n13103, n13105, n13222, n13112,
    n13109, n13108, n13110, n13359, n13162, n13111, n13128, n13115, n13374,
    n16613, n13116, n16899, n13119, n13118, n13120, n13125, n13123, n13122,
    n13124, n13127, n13126, n13129, n13136, n13134, n13132, n13131, n13133,
    n13135, n13141, n13138, n13140, n13142, n13148, n13146, n13145, n13150,
    n13149, n13154, n13151, n13153, n13159, n13157, n13156, n13158, n13168,
    n13164, n13161, n13163, n13165, n13167, n13171, n13170, n13177, n13175,
    n13174, n13194, n13179, n13178, n13183, n13181, n13182, n13186, n13187,
    n13395, n13190, n13188, n13393, n13189, n13191, n13192, n13193, n13198,
    n13200, n13202, n13201, n13213, n13211, n13205, n13207, n13209, n13208,
    n13210, n13212, n13215, n13214, n13219, n13238, n13217, n13216, n13218,
    n13236, n13588, n13590, n13220, n13221, n13224, n13589, n13237, n13233,
    n13226, n13340, n13227, n13232, n13230, n13229, n13231, n13234, n13235,
    n13246, n13242, n13240, n13239, n13241, n13243, n13245, n13249, n13248,
    n13255, n13253, n13252, n13254, n13259, n13257, n13258, n13262, n13261,
    n13263, n13264, n13270, n13437, n13268, n13267, n13272, n13271, n13275,
    n13284, n13277, n13279, n13278, n13282, n13281, n13283, n13287, n13286,
    n13290, n13292, n13291, n13304, n13302, n13300, n13296, n13298, n13299,
    n13301, n13303, n13306, n13305, n13308, n13307, n13316, n13490, n13314,
    n13311, n13310, n13313, n13315, n13326, n13321, n13319, n13318, n13320,
    n13324, n13322, n13323, n13494, n13325, n13328, n13327, n13333, n13331,
    n13330, n13332, n13339, n13337, n13336, n13338, n13341, n16991, n13348,
    n13344, n13343, n13346, n13345, n13347, n13363, n13349, n13351, n16910,
    n13580, n13352, n13356, n13354, n13353, n13355, n13357, n13610, n13408,
    n13360, n13361, n13362, n13382, n13434, n13369, n13367, n13426, n13368,
    n13380, n13423, n13378, n13373, n13372, n13377, n13375, n13376, n13379,
    n13381, n13385, n13384, n13389, n13392, n13391, n13403, n13394, n13398,
    n13400, n13402, n13406, n13405, n13416, n13412, n13410, n13409, n13411,
    n13413, n13415, n13419, n13418, n13422, n13421, n13433, n13431, n13429,
    n13427, n13428, n13430, n13432, n13436, n13435, n13447, n13440, n13439,
    n13441, n13445, n13444, n13446, n13450, n13449, n13454, n13457, n13456,
    n13470, n13460, n13464, n13463, n13466, n13468, n13467, n13469, n13472,
    n13471, n13478, n13476, n13475, n13477, n13480, n13482, n13481, n13489,
    n13487, n13488, n13499, n13492, n13491, n13493, n13502, n13505, n17093,
    n13504, n13507, n13506, n13510, n13509, n13512, n13511, n13514, n13516,
    n13515, n13527, n13525, n13523, n13519, n13521, n13522, n13526, n13528,
    n13544, n13533, n13534, n13542, n13539, n13540, n13541, n13546, n13545,
    n13562, n13551, n13553, n13552, n13560, n13557, n13558, n13559, n13564,
    n13563, n13579, n13567, n13569, n13577, n13571, n13573, n13572, n13575,
    n13574, n13576, n13578, n13781, n13582, n13585, n13584, n13586, n13591,
    n13789, n13788, n13609, n13605, n13603, n13602, n13604, n13607, n13606,
    n13613, n13793, n13658, n13612, n13615, n13617, n13624, n13622, n13621,
    n13623, n13636, n13632, n13630, n13629, n13631, n13634, n13633, n13639,
    n13671, n13638, n13641, n13644, n13643, n13651, n13647, n13649, n13652,
    n13655, n13666, n13662, n13660, n13659, n13661, n13669, n13679, n13675,
    n13673, n13672, n13674, n13682, n13685, n13684, n13687, n13686, n13694,
    n13739, n13692, n13691, n13693, n13704, n13698, n13697, n13699, n13703,
    n13706, n13711, n13716, n13714, n13713, n13736, n13718, n13724, n13721,
    n13722, n13723, n13733, n13726, n13725, n13727, n13748, n13744, n13742,
    n13741, n13751, n13755, n13754, n13756, n14528, n13758, n13769, n13767,
    n13764, n13762, n13765, n13766, n13768, n13780, n13777, n13775, n13778,
    n13779, n13801, n13785, n13784, n13786, n13791, n13790, n13798, n13794,
    n13795, n13831, n13796, n13797, n13799, n13804, n13807, n13809, n13828,
    n13816, n13813, n13814, n13815, n13824, n13822, n13820, n13821, n13823,
    n13825, n13835, n13833, n13836, n13841, n13839, n13838, n13840, n13843,
    n13863, n13849, n13848, n13850, n13851, n13859, n13854, n13857, n13856,
    n13858, n13860, n13868, n13870, n13872, n13871, n13887, n13879, n13881,
    n13880, n13883, n14449, n13885, n13884, n13888, n13898, n13891, n13901,
    n13904, n13903, n13905, n13912, n13913, n13933, n13914, n13919, n13922,
    n13926, n13925, n13929, n13928, n13930, n13935, n13934, n13936, n13939,
    n13941, n13945, n13948, n13951, n13950, n13959, n13953, n13956, n13954,
    n13964, n13962, n13966, n14131, n13967, n13970, n13969, n14025, n13976,
    n13975, n13977, n13980, n13987, n13984, n13990, n13989, n13991, n13998,
    n13999, n14000, n14009, n14004, n14003, n14006, n14013, n14019, n14022,
    n14033, n14029, n14027, n14028, n14036, n14040, n14039, n14041, n14044,
    n14043, n14046, n14045, n14056, n14055, n14057, n14059, n14065, n14064,
    n14066, n14075, n14076, n14084, n14081, n14085, n14089, n14088, n14090,
    n14097, n14100, n14105, n14107, n14111, n14114, n14118, n14124, n14127,
    n14135, n14134, n14280, n14138, n14137, n14140, n14139, n14141, n16671,
    n14143, n16653, n14145, n16650, n14265, n14153, n14152, n14154, n14295,
    n14160, n14179, n14166, n14169, n14168, n14177, n14174, n14249, n14172,
    n14173, n14180, n14196, n14185, n14192, n14190, n14188, n14189, n14191,
    n14193, n14200, n14199, n14201, n14210, n14213, n14224, n14220, n14219,
    n14222, n14221, n14223, n14231, n14232, n14392, n14238, n14240, n14260,
    n14244, n14246, n14245, n14258, n14250, n14253, n14254, n14262, n14346,
    n14268, n14286, n14269, n14272, n14271, n14273, n14276, n14282, n14281,
    n14356, n14285, n14481, n14289, n14292, n14304, n14298, n14297, n14307,
    n14309, n14315, n14313, n14312, n14314, n14324, n14322, n14327, n14326,
    n14341, n14332, n14330, n14335, n14334, n14337, n14546, n14339, n14338,
    n14342, n14345, n14351, n14350, n14352, n14361, n14359, n14360, n14372,
    n14366, n14364, n14363, n14365, n14367, n14374, n14373, n14379, n14382,
    n14389, n14400, n14394, n14393, n14403, n14406, n14405, n14407, n14410,
    n14412, n14414, n14423, n14559, n14558, n14418, n14417, n14419, n14420,
    n14431, n14564, n14563, n14428, n14427, n14429, n14430, n14446, n14438,
    n14441, n14454, n14450, n14452, n14451, n14453, n14455, n14460, n14465,
    n14468, n14473, n14472, n14474, n14477, n14483, n14604, n14487, n14490,
    n14493, n14499, n14497, n14496, n14498, n14514, n14507, n14556, n14509,
    n14508, n14512, n14511, n14513, n14521, n14533, n14531, n14529, n14530,
    n14532, n14534, n14537, n14552, n14550, n14548, n14545, n14547, n14549,
    n14551, n14553, n14555, n14571, n14867, n14874, n14572, n14579, n14578,
    n14580, n14587, n14584, n14586, n14588, n14668, n14595, n14594, n14596,
    n14602, n14607, n14683, n14611, n14614, n14798, n14616, n14626, n14624,
    n14618, n14630, n14621, n14619, n14622, n14636, n14629, n14633, n14631,
    n14634, n14635, n14648, n14641, n14866, n14644, n14643, n14646, n14645,
    n14649, n14652, n14653, n14660, n14663, n14662, n14730, n14672, n14671,
    n14673, n14675, n14678, n14677, n14679, n14685, n14747, n14696, n14699,
    n14710, n14713, n14727, n14721, n14720, n14723, n14722, n14725, n16877,
    n17012, n14907, n14734, n14733, n14735, n14737, n14741, n14740, n14742,
    n14750, n14923, n14755, n14761, n14764, n14773, n14772, n14774, n14778,
    n14782, n14781, n14785, n14793, n14805, n14803, n14801, n14799, n14800,
    n14802, n14806, n14816, n14819, n14824, n14821, n14851, n14832, n14829,
    n14838, n14843, n14861, n14857, n14855, n14854, n14856, n14858, n14865,
    n14886, n14872, n14869, n14880, n14877, n14888, n14903, n14897, n14896,
    n14899, n16311, n14898, n14901, n17014, n14967, n14911, n14910, n14912,
    n14914, n14918, n14917, n14919, n14926, n14932, n14939, n14942, n14956,
    n14954, n14950, n14949, n14951, n14959, n14960, n14964, n15370, n14963,
    n14965, n17016, n15153, n14971, n14970, n14972, n15158, n14988, n14985,
    n14999, n15006, n15004, n15007, n15021, n15015, n15014, n15017, n15016,
    n15019, n15026, n15050, n15033, n15032, n15034, n15038, n15042, n15041,
    n15045, n15058, n15061, n15064, n15073, n15071, n15074, n15079, n15096,
    n15090, n15089, n15091, n15093, n15102, n15124, n15107, n15106, n15108,
    n15112, n15117, n15116, n15126, n15132, n15135, n15150, n15144, n15143,
    n15146, n15145, n15148, n15147, n15297, n15156, n15162, n15305, n15164,
    n15192, n15168, n15176, n15178, n15188, n15187, n15193, n15196, n15199,
    n15200, n16520, n15204, n15760, n15207, n15206, n15740, n15219, n15208,
    n15216, n15215, n16836, n15220, n15221, n15228, n15237, n15233, n15232,
    n15234, n15238, n15243, n15249, n15252, n15255, n15260, n15259, n16411,
    n15962, n15262, n15835, n15377, n15263, n15264, n15462, n16018, n15273,
    n15277, n15479, n15280, n15279, n15284, n15286, n15290, n15294, n15391,
    n16857, n15302, n15301, n15303, n15307, n15401, n15329, n15310, n15317,
    n15315, n15318, n15324, n15332, n15330, n15333, n15340, n15339, n15347,
    n15345, n15348, n15356, n15354, n15357, n15366, n15364, n15367, n15373,
    n15376, n15378, n15388, n15386, n15389, n15392, n16864, n17026, n15592,
    n15398, n15397, n15399, n15403, n15601, n15428, n15413, n15415, n15425,
    n15431, n15429, n15432, n15437, n15447, n15441, n15440, n15443, n15442,
    n15444, n15458, n15456, n15459, n15560, n15942, n15470, n15469, n15477,
    n15475, n15474, n15476, n15480, n15545, n15498, n15489, n15501, n15499,
    n15502, n15507, n15520, n15518, n15514, n15513, n15515, n15541, n15534,
    n15533, n15537, n15536, n15538, n16030, n15546, n15551, n15664, n15555,
    n15706, n15866, n15570, n15567, n15571, n15589, n15580, n15583, n15586,
    n15633, n15597, n15596, n15603, n15644, n15627, n15606, n15614, n15612,
    n15611, n15630, n15628, n15631, n16947, n15734, n15638, n15637, n15678,
    n15641, n15649, n15668, n15666, n15669, n15681, n15679, n15682, n15701,
    n15693, n15692, n15694, n15698, n15823, n16406, n16414, n16022, n15715,
    n15714, n15783, n15721, n15726, n16861, n15735, n15737, n17064, n16951,
    n17023, n15744, n15742, n15741, n15798, n15746, n15750, n15753, n15749,
    n15757, n15755, n15754, n15756, n15772, n15767, n15786, n15784, n15787,
    n15797, n15799, n15803, n15802, n15808, n15807, n15818, n15814, n15813,
    n15815, n15819, n15827, n16499, n15842, n15947, n15831, n15838, n15836,
    n15837, n15841, n16509, n15844, n15843, n15856, n15851, n15862, n15864,
    n15880, n15878, n15871, n15870, n15874, n15873, n15875, n16462, n16305,
    n15885, n15886, n15911, n15896, n15898, n15900, n15903, n15908, n16308,
    n15921, n15923, n15927, n15933, n15937, n15939, n15944, n15950, n15956,
    n15951, n15952, n15957, n15963, n16463, n16041, n15964, n16482, n16033,
    n15974, n15973, n15980, n15978, n15979, n15982, n15983, n15985, n15987,
    n15990, n15991, n15993, n15995, n15999, n15998, n16000, n16002, n16004,
    n16005, n16007, n16009, n16011, n16013, n16015, n16017, n16035, n16034,
    n16047, n16040, n16042, n16050, n16049, n16052, n16058, n16055, n16057,
    n16059, n16060, n16065, n16064, n16066, n16069, n16068, n16100, n16072,
    n16075, n16074, n16092, n16077, n16078, n16089, n16083, n16086, n16085,
    n16099, n16088, n16098, n16096, n16105, n16094, n16095, n16097, n16103,
    n16101, n16107, n16123, n16109, n16108, n16122, n16121, n16113, n16112,
    n16114, n16139, n16118, n16117, n16119, n16120, n16131, n16129, n16127,
    n16126, n16128, n16130, n16159, n16133, n16134, n16138, n16137, n16142,
    n16140, n16141, n16157, n16144, n16155, n16149, n16153, n16152, n16154,
    n16156, n16158, n16172, n16163, n16162, n16182, n16170, n16168, n16167,
    n16169, n16171, n16187, n16174, n16173, n16179, n16178, n16210, n16184,
    n16183, n16185, n16186, n16218, n16191, n16190, n16193, n16197, n16196,
    n16202, n16200, n16201, n16216, n16204, n16208, n16207, n16214, n16211,
    n16213, n16215, n16224, n16222, n16221, n16223, n16234, n16228, n16227,
    n16232, n16231, n16237, n16233, n16242, n16236, n16235, n16240, n16239,
    n16241, n16258, n16246, n16245, n16250, n16249, n16256, n16254, n16253,
    n16255, n16262, n16261, n16269, n16264, n16263, n16271, n16267, n16268,
    n16276, n16274, n16283, n16278, n16281, n16284, n16282, n16288, n16286,
    n16287, n16289, n16291, n16307, n16297, n16295, n16296, n16304, n16301,
    n16300, n16303, n16315, n16310, n16309, n16313, n16314, n16327, n16330,
    n16320, n16319, n16318, n16326, n16324, n16323, n16325, n16344, n16332,
    n16331, n16336, n16335, n16340, n16339, n16343, n16357, n16346, n16345,
    n16349, n16352, n16361, n16360, n16371, n16365, n16364, n16369, n16368,
    n16377, n16384, n16381, n16380, n16402, n16389, n16388, n16397, n16395,
    n16394, n16396, n16404, n16440, n16438, n16407, n16419, n16409, n16408,
    n16428, n16412, n16418, n16416, n16445, n16424, n16420, n16421, n16435,
    n16431, n16430, n16433, n16448, n16437, n16441, n16456, n16460, n16475,
    n16470, n16473, n16476, n16480, n16484, n16483, n16485, n16497, n16490,
    n16489, n16495, n16493, n16494, n16496, n16507, n16508, n16515, n16513,
    n16512, n16518, n16517, n16519, n16522, n16521, n16800, n16526, n16525,
    n16821, n16533, n16688, n16532, n16536, n16542, n16539, n16538, n16541,
    n16550, n16551, n16556, n16555, n16557, n16560, n16559, n16566, n16571,
    n16564, n16565, n16578, n16570, n16573, n17038, n16572, n16576, n16575,
    n16577, n16586, n16580, n16584, n16582, n16583, n16585, n16594, n16588,
    n16587, n16592, n16591, n16593, n16602, n16893, n16597, n16600, n16900,
    n16599, n16601, n16608, n16604, n16603, n16605, n16607, n16612, n16610,
    n16611, n16615, n16907, n16614, n16621, n16619, n16618, n16620, n16623,
    n16622, n16626, n16625, n16635, n16633, n16631, n16630, n16632, n16634,
    n16642, n16636, n16638, n16640, n16639, n16641, n16646, n16644, n16647,
    n16649, n16652, n16651, n16665, n16654, n16655, n16681, n16658, n16663,
    n16662, n16664, n16670, n16667, n16669, n16675, n16674, n16676, n16679,
    n16682, n16683, n16686, n16685, n16691, n16690, n16695, n16694, n16703,
    n16702, n16704, n16710, n16715, n16714, n16719, n16718, n16722, n16725,
    n16724, n16730, n16733, n16740, n16743, n16742, n16751, n16750, n16761,
    n16753, n16755, n16766, n16769, n16773, n16772, n16774, n16780, n16779,
    n16784, n16783, n16809, n16791, n16790, n16789, n16792, n16793, n16795,
    n16797, n16802, n16833, n16954, n16826, n16831, n16828, n16838, n17036,
    n17031, n16850, n16848, n16852, n16966, n16855, n16858, n16871, n16876,
    n16927, n16883, n17004, n16882, n16930, n16886, n17008, n16889, n16895,
    n16891, n16894, n16898, n16932, n16897, n16906, n16904, n16902, n16903,
    n16905, n16908, n16909, n16911, n16913, n16912, n16917, n16916, n16918,
    n16920, n16921, n16923, n16924, n16925, n16926, n16928, n17048, n16942,
    n16938, n16933, n16936, n16937, n16939, n16941, n16943, n16944, n16948,
    n16952, n16968, n17083, n16970, n16973, n16978, n17040, n16977, n16980,
    n16982, n16984, n16986, n16988, n16990, n16992, n16993, n16995, n16997,
    n16999, n17001, n17003, n17006, n17007, n17009, n17011, n17015, n17017,
    n17019, n17039, n17042, n17044, n17045, n17047, n17068, n17074, n17082,
    n17085, n17101, n17088, n17090, n17095, n17094, n17098, n17097, n17099,
    n17100, n17105, n17113, n17129, n17140, n17134, n17133, n17138, n17137,
    n17139, n17141, n17152, n17151;
  assign n15720 = ~n15488;
  assign n15434 = ~n11243 | ~n11244;
  assign n15465 = ~n15462 & ~n15461;
  assign n17063 = ~n15199 | ~n15198;
  assign n15298 = ~n15297 | ~n15296;
  assign n16449 = ~n15256 | ~n15255;
  assign n11236 = ~n11235 & ~n11234;
  assign n15154 = ~n15153 | ~n17016;
  assign n11075 = ~n11070 | ~n11069;
  assign n14968 = n14967 | n17014;
  assign n16854 = ~n16524;
  assign n16503 = ~n15260 | ~n15259;
  assign n14908 = ~n14907 & ~n16877;
  assign n14669 = ~n14668 & ~n16887;
  assign n11217 = ~n14518 | ~n14516;
  assign n14590 = n14470 & n16885;
  assign n14470 = ~n14268 | ~n14286;
  assign n14225 = ~n13956 | ~n16996;
  assign n14997 = ~n11098 & ~n11097;
  assign n14048 = ~n10563 | ~n10562;
  assign n16302 = ~n11092 | ~n11632;
  assign n13952 = ~n13582 | ~n16637;
  assign n15914 = ~n10236 | ~n10235;
  assign n14510 = ~n10617 | ~n10616;
  assign n14447 = ~n10570 & ~n10569;
  assign n13350 = ~n13119 & ~n16985;
  assign n13117 = ~n13374 & ~n16983;
  assign n10922 = ~n13206 | ~n13204;
  assign n13206 = ~n10917 | ~n13022;
  assign n13024 = ~n12649 & ~n10912;
  assign n12651 = ~n12619 | ~n10908;
  assign n12618 = ~n10903 & ~n10902;
  assign n11296 = ~n10887 & ~n10886;
  assign n9179 = ~n9175 ^ n17107;
  assign n9035 = ~n9040;
  assign n15212 = ~n9183;
  assign n16491 = n10640 ^ P2_IR_REG_22__SCAN_IN;
  assign n10630 = ~n10611 | ~P2_IR_REG_31__SCAN_IN;
  assign n10586 = n14404 & n16487;
  assign n10639 = ~n10632 | ~n10635;
  assign n10239 = ~n14961 | ~P2_IR_REG_31__SCAN_IN;
  assign n10632 = ~n10564 & ~n10190;
  assign n9106 = ~n9105 & ~n9733;
  assign n10237 = ~n10227 | ~n10226;
  assign n10209 = ~n10232 | ~n10205;
  assign n9304 = ~n9189 & ~P1_IR_REG_2__SCAN_IN;
  assign n9092 = ~n9053 & ~n9052;
  assign n9044 = ~P1_IR_REG_0__SCAN_IN;
  assign n9093 = ~P1_IR_REG_9__SCAN_IN & ~P1_IR_REG_8__SCAN_IN;
  assign n10261 = ~P2_IR_REG_0__SCAN_IN;
  assign n11222 = ~n14637 & ~n14638;
  assign n13555 = ~n10927 | ~n13295;
  assign n10973 = ~n10951 | ~n14252;
  assign n11232 = ~n11228 | ~n14890;
  assign n11251 = ~n11250 & ~n15524;
  assign n11212 = ~n11206 & ~n11205;
  assign n11012 = ~n10979 | ~n10978;
  assign n11227 = ~n14718 | ~n14715;
  assign n11238 = ~n15140 | ~n15138;
  assign n10891 = n12351 ^ n11296;
  assign n10278 = ~n10276 & ~n10275;
  assign n10940 = ~n13648;
  assign n15395 = ~n15392 & ~n16857;
  assign n15634 = ~n15633 | ~n17054;
  assign n10224 = ~n9170;
  assign P1_U3520 = ~n15803 | ~n15802;
  assign P1_U3552 = ~n15808 | ~n15807;
  assign n15739 = ~n15737 ^ n17023;
  assign n12522 = ~n12542;
  assign n14731 = ~n14730 | ~n16879;
  assign n14266 = ~n14346 | ~n16940;
  assign n9169 = ~n9183 & ~n9162;
  assign n16976 = ~n16563;
  assign n13581 = ~n13580 | ~n16915;
  assign n10768 = ~n12553 & ~n16969;
  assign n10771 = ~n12449 | ~n16888;
  assign n10769 = ~n16896;
  assign n10772 = ~n12362 | ~n12373;
  assign n15960 = ~n15965;
  assign n9666 = ~n13852 | ~n9630;
  assign n16048 = ~n11295 & ~n11294;
  assign n10578 = ~n14048 | ~n16001;
  assign n15160 = ~n9953 | ~n9952;
  assign n16778 = ~n16782;
  assign n12043 = ~n9072 | ~n14583;
  assign n15201 = ~n15257 | ~n15212;
  assign n17018 = ~n17051 | ~n16771;
  assign n10796 = ~n17073 | ~n17037;
  assign n9112 = ~n9111 & ~P2_RD_REG_SCAN_IN;
  assign n9915 = ~n9898 | ~n9897;
  assign n11207 = ~n11023 & ~n11022;
  assign n11315 = ~n9035 | ~n15724;
  assign n11191 = ~n9035 | ~n15529;
  assign n11121 = ~n9035 | ~n15040;
  assign n16502 = ~n12855 | ~n10883;
  assign n14216 = ~n14131 | ~n14130;
  assign n16124 = ~n10309 & ~n10308;
  assign n15961 = ~n15373 & ~n15372;
  assign n15850 = ~n12004 | ~n11612;
  assign n15845 = ~n15720 | ~n15272;
  assign n11089 = ~n9034;
  assign n16957 = ~n17063;
  assign n15763 = ~n15745 | ~n13968;
  assign n15867 = ~n10965 | ~n15850;
  assign n15488 = ~n10728 & ~n15725;
  assign n15369 = ~n11075 ^ n11074;
  assign n13390 = P2_U3152 | n11635;
  assign n11613 = ~n11612 | ~n11611;
  assign n12117 = ~n10175 | ~n10174;
  assign n10309 = ~n10305 | ~n10304;
  assign n9209 = n9205 ^ n17107;
  assign n9205 = ~n9204 | ~n9203;
  assign n9138 = ~n12534 | ~n17104;
  assign n12534 = ~n9076 | ~n9043;
  assign n11807 = ~n11061 & ~n14576;
  assign n10256 = ~n10476 | ~P2_REG2_REG_0__SCAN_IN;
  assign n9033 = ~n11274;
  assign n9180 = ~n9179;
  assign n12537 = ~n9178 | ~n9179;
  assign n12806 = ~n10888;
  assign n15733 = ~n15722 | ~n15721;
  assign n15722 = ~n15783 | ~n15720;
  assign n15782 = ~n15781 & ~n15780;
  assign n16481 = ~n16047 | ~n16046;
  assign n15732 = ~n15731 & ~n15730;
  assign n16477 = n16475 | n16470;
  assign n15781 = ~n15775 & ~n16498;
  assign n17081 = ~n17077 & ~n17076;
  assign n15490 = ~n15477 & ~n15476;
  assign n16037 = ~n16034 | ~n16038;
  assign n15573 = ~n15572 & ~n15571;
  assign n17080 = ~n17079 & ~n17089;
  assign n15703 = ~n15688 | ~n10132;
  assign n16046 = ~n16045 & ~n16044;
  assign n15663 = ~n15658 & ~n15657;
  assign n17077 = ~n17034 & ~n17073;
  assign n15572 = ~n15658 & ~n15563;
  assign n16467 = ~n16460 | ~n16459;
  assign n17076 = ~n17075 & ~n17074;
  assign n17034 = ~n17033 & ~n17037;
  assign n16840 = ~n16835 | ~n16834;
  assign n16045 = ~n16482 & ~n16391;
  assign n16044 = ~n16043 | ~n16042;
  assign n15496 = ~n15491 & ~n16498;
  assign n16036 = ~n16035 | ~n16472;
  assign n15543 = ~n15528 | ~n15527;
  assign n15368 = ~n15366 | ~n15800;
  assign n15449 = ~n15438 | ~n15527;
  assign n15522 = ~n15508 | ~n10132;
  assign n15349 = ~n15347 | ~n16514;
  assign n15485 = ~n15478 | ~n10644;
  assign n16835 = ~n16831 | ~n16830;
  assign n15346 = ~n15347 | ~n16510;
  assign n15295 = ~n15293 | ~n15720;
  assign n16846 = ~n16845 | ~n16844;
  assign n15591 = ~n15577 | ~n10132;
  assign n15365 = ~n15366 | ~n15804;
  assign n16043 = ~n16041 | ~n16040;
  assign n15136 = ~n15134 | ~n16510;
  assign n17032 = ~n17031 | ~n17030;
  assign n15677 = ~n15676 & ~n15675;
  assign n15253 = ~n15251 | ~n16510;
  assign n15618 = ~n15607 | ~n15606;
  assign n16834 = ~n16833 | ~n16832;
  assign n15655 = ~n15654 & ~n15653;
  assign n15123 = ~n15113 | ~n15112;
  assign n16965 = ~n16964 | ~n16963;
  assign n15133 = ~n15134 | ~n16514;
  assign n15774 = ~n15747 | ~n15746;
  assign n16845 = ~n16841 | ~n16688;
  assign n15293 = ~n15292 | ~n15291;
  assign n15250 = ~n15251 | ~n16514;
  assign n17071 = ~n17069 | ~n17068;
  assign n16459 = ~n16458 | ~n16457;
  assign n16466 = ~n16465 | ~n16464;
  assign n15251 = ~n15248 | ~n15247;
  assign n16849 = ~n17036 & ~n17093;
  assign n15134 = ~n15131 | ~n15130;
  assign n15223 = ~n15222 & ~n15221;
  assign n16964 = ~n16961 | ~n17070;
  assign n15344 = ~n15336 | ~n15335;
  assign n15654 = ~n15671 & ~n15758;
  assign n17069 = ~n17036 & ~n17035;
  assign n15292 = ~n15336 | ~n15273;
  assign n11204 = ~n11184 | ~n11183;
  assign n15747 = ~n15798 | ~n15745;
  assign n16464 = ~n16463 | ~n16391;
  assign n15966 = ~n15965 & ~n15964;
  assign n15358 = ~n15356 | ~n15800;
  assign n16961 = ~n16960 | ~n16959;
  assign n15222 = ~n16839 & ~n15763;
  assign n15574 = ~n15556 | ~n15555;
  assign n15355 = ~n15356 | ~n15804;
  assign n11184 = ~n15242 | ~n14047;
  assign n15059 = ~n15060 | ~n16514;
  assign n16457 = ~n16463 | ~n16461;
  assign n15248 = ~n15242 | ~n15335;
  assign n15433 = ~n15431 | ~n15800;
  assign n17070 = ~n16842;
  assign n15131 = ~n15111 & ~n15110;
  assign n15840 = ~n15833 | ~n15832;
  assign n15122 = ~n15121 & ~n15120;
  assign n15420 = ~n15416 | ~n15415;
  assign n15049 = ~n15039 | ~n15038;
  assign n15390 = ~n15388 | ~n16510;
  assign n15062 = ~n15060 | ~n16510;
  assign n15656 = ~n15642 | ~n15641;
  assign n15387 = ~n15388 | ~n16514;
  assign n15241 = ~n15229 | ~n10132;
  assign n15430 = ~n15431 | ~n15804;
  assign n15617 = ~n15616 & ~n15615;
  assign n16029 = ~n16028 & ~n16027;
  assign n17030 = ~n17029 & ~n17028;
  assign n15129 = ~n15124 & ~n16498;
  assign n15111 = ~n15124 & ~n14769;
  assign n15965 = ~n16462 | ~n15952;
  assign n16960 = ~n16955 | ~n16954;
  assign n15416 = ~n15428 | ~n15414;
  assign n16465 = ~n16462 | ~n16461;
  assign n15642 = ~n15678 | ~n15745;
  assign n16458 = ~n16462 | ~n16391;
  assign n16839 = ~n16836;
  assign n16455 = ~n16454 | ~n16453;
  assign n15556 = ~n15664 | ~n15720;
  assign n16842 = ~n16836 & ~n16837;
  assign n15380 = ~n15379 & ~n15378;
  assign n17145 = ~n17144 | ~n17143;
  assign n15048 = ~n15047 & ~n15046;
  assign n16806 = ~n16805 & ~n16804;
  assign n16454 = ~n16451 | ~n16450;
  assign n16958 = ~n16956;
  assign n16423 = ~n16422 & ~n16421;
  assign n9968 = ~n9942 & ~n15226;
  assign n15334 = ~n15332 | ~n15804;
  assign n15056 = ~n15055 & ~n15054;
  assign n15453 = ~n15961 & ~n15451;
  assign n16447 = ~n16446 | ~n16445;
  assign n15968 = ~n15961;
  assign n15057 = ~n15037 & ~n15036;
  assign n15379 = ~n15961 & ~n15848;
  assign n15210 = ~n15209 & ~n15208;
  assign n15419 = ~n15418 & ~n15417;
  assign n15321 = ~n15311 | ~n15310;
  assign n15266 = ~n15265 & ~n15264;
  assign n15959 = ~n15958 | ~n15957;
  assign n16824 = ~n16823 & ~n16822;
  assign n15331 = ~n15332 | ~n15800;
  assign n15037 = ~n15050 & ~n14769;
  assign n16832 = n16827 & n16826;
  assign n15640 = ~n15635 & ~n15738;
  assign n15055 = ~n15050 & ~n16498;
  assign n15217 = ~n16957 | ~n15760;
  assign n15183 = ~n15169 | ~n15168;
  assign n15418 = ~n15421 & ~n15608;
  assign n15771 = ~n15770 | ~n15769;
  assign n15830 = ~n15947 | ~n15829;
  assign n15008 = ~n15006 | ~n16510;
  assign n15958 = ~n15956 | ~n15955;
  assign n15209 = ~n16957 & ~n15763;
  assign n15405 = ~n15421 & ~n15404;
  assign n15265 = ~n16432 & ~n15848;
  assign n15351 = ~n16957 & ~n15422;
  assign n11140 = ~n11131 & ~n11130;
  assign n15796 = ~n15795 | ~n15794;
  assign n15005 = ~n15006 | ~n16514;
  assign n16027 = ~n16026 | ~n16025;
  assign n15711 = ~n15710 | ~n15829;
  assign n14966 = ~n15213 | ~n11059;
  assign n15197 = ~n15195 | ~n15804;
  assign n17144 = ~n17125 | ~n17124;
  assign n16451 = ~n16432 | ~n16452;
  assign n15554 = ~n15548 & ~n15547;
  assign n15194 = ~n15195 | ~n15800;
  assign n15152 = ~n15141 | ~n15527;
  assign n16805 = ~n16800 & ~n16799;
  assign n16830 = ~n16829 | ~n16828;
  assign n16956 = ~n16953 | ~n17064;
  assign n16446 = ~n16444 | ~n16443;
  assign n16953 = ~n16952 | ~n17059;
  assign n15320 = ~n15319 & ~n15318;
  assign n15855 = ~n15854 | ~n15853;
  assign n15955 = ~n16449 & ~n15954;
  assign n11083 = ~n15369 & ~n14384;
  assign n17121 = ~n17148 | ~n17120;
  assign n17067 = ~n17061 & ~n17060;
  assign n15195 = ~n15192 | ~n15191;
  assign n17149 = ~n17148 & ~n17147;
  assign n15213 = ~n15369;
  assign n16799 = ~n16798 & ~n16797;
  assign n17025 = ~n17023 | ~n17022;
  assign n15795 = ~n15792 | ~n15791;
  assign n15375 = ~n16449 & ~n15374;
  assign n16443 = ~n16442 | ~n16441;
  assign n16506 = ~n16505 | ~n16504;
  assign n15769 = ~n15768 & ~n15767;
  assign n15730 = ~n15729 | ~n15728;
  assign n15653 = ~n15652 | ~n15651;
  assign n15002 = ~n15001 | ~n15000;
  assign n11342 = n11341 & n11340;
  assign n15792 = ~n15761 & ~n15760;
  assign n15098 = ~n15084 | ~n10132;
  assign n11065 = ~n11060 & ~n14094;
  assign n16417 = ~n16416 & ~n16415;
  assign n15291 = ~n15342 & ~n15290;
  assign n16529 = ~n16528 | ~n16527;
  assign n15308 = ~n15322 & ~n15404;
  assign n15319 = ~n15322 & ~n15608;
  assign n16798 = ~n16796 | ~n16795;
  assign n15483 = ~n15481 & ~n15547;
  assign n17060 = ~n17059;
  assign n11058 = ~n11060 & ~n14384;
  assign n16444 = ~n16438 | ~n16437;
  assign n15853 = ~n15852 & ~n15851;
  assign n17061 = ~n17058 & ~n17057;
  assign n11139 = ~n11138 | ~n11137;
  assign n15675 = ~n15674 | ~n15673;
  assign n15182 = ~n15181 & ~n15180;
  assign n15728 = ~n15727 & ~n15726;
  assign n15780 = ~n15779 | ~n15778;
  assign n15949 = ~n15948 & ~n16414;
  assign n15374 = ~n16411 | ~n15846;
  assign n17124 = ~n17123 & ~n17147;
  assign n16528 = ~n16523 & ~n16950;
  assign n15256 = ~n15254 | ~n10310;
  assign n11322 = ~n11324 & ~n11321;
  assign n16505 = ~n16501 | ~n16500;
  assign n11129 = ~n14994 | ~n10644;
  assign n17143 = ~n17142 & ~n17141;
  assign n15481 = ~n15545 ^ n16020;
  assign n15400 = ~n15396 | ~n15592;
  assign n16801 = ~n17064;
  assign n15023 = ~n15013 | ~n15527;
  assign n17058 = ~n16862 | ~n16861;
  assign n16823 = ~n16820 & ~n16819;
  assign n15001 = ~n14994 | ~n14993;
  assign n15651 = ~n15650 & ~n15649;
  assign n11203 = ~n11202 & ~n11201;
  assign n15674 = ~n15672 | ~n15791;
  assign n15181 = ~n15184 & ~n15608;
  assign n11340 = ~n11339 & ~n11338;
  assign n11338 = ~n11337 | ~n11336;
  assign n15672 = ~n15648 & ~n15759;
  assign n15282 = ~n15278 | ~n15832;
  assign n14817 = ~n14818 | ~n16510;
  assign n14789 = ~n14779 | ~n14778;
  assign n16504 = ~n16503 | ~n16502;
  assign n15165 = ~n15170 | ~n15163;
  assign n15396 = ~n15394 & ~n15738;
  assign n14820 = ~n14818 | ~n16514;
  assign n15184 = ~n15170;
  assign n11344 = ~n11323 & ~n15861;
  assign n15948 = ~n16503 & ~n16410;
  assign n17142 = ~n17127 & ~n17126;
  assign n15075 = ~n15073 | ~n15800;
  assign n17120 = ~n17122 & ~n17147;
  assign n14958 = ~n14946 | ~n10132;
  assign n17115 = ~n17114 | ~n17113;
  assign n16794 = ~n16950;
  assign n15953 = ~n16503 | ~n16410;
  assign n16425 = ~n16414;
  assign n17123 = ~n17122;
  assign n15072 = ~n15073 | ~n15804;
  assign n17108 = ~n17106 | ~n17105;
  assign n15083 = ~n15079 & ~n15078;
  assign n15779 = ~n15776 | ~n16500;
  assign n15414 = ~n15413 & ~n15412;
  assign n14711 = ~n14712 | ~n16514;
  assign n15615 = ~n15614 | ~n15613;
  assign n15394 = ~n15395 & ~n17026;
  assign n14714 = ~n14712 | ~n16510;
  assign n17057 = ~n17056 & ~n17055;
  assign n17122 = ~n17119 & ~n17118;
  assign n11066 = n11068 ^ n11067;
  assign n15648 = n15647 & n17110;
  assign n14991 = ~n14990 & ~n14989;
  assign n15759 = ~n15647 & ~n17110;
  assign n14807 = ~n14794 | ~n10132;
  assign n15613 = ~n15612 & ~n15611;
  assign n15879 = ~n15878 & ~n15877;
  assign n15304 = ~n15300 | ~n10774;
  assign n14940 = ~n14941 | ~n15804;
  assign n15859 = ~n11301 & ~n11324;
  assign n15069 = ~n15068 & ~n15789;
  assign n14814 = ~n14813 & ~n14812;
  assign n11068 = ~n11051 | ~n11050;
  assign n14943 = ~n14941 | ~n15800;
  assign n15821 = ~n15820 & ~n15819;
  assign n11200 = ~n11189 | ~n15832;
  assign n14863 = ~n14849 | ~n10132;
  assign n10741 = ~n10737 | ~n10736;
  assign n15624 = ~n15623 | ~n15622;
  assign n10172 = ~n10171 & ~n10170;
  assign n14788 = ~n14787 & ~n14786;
  assign n15643 = ~n16854 | ~n17135;
  assign n14813 = ~n14808 & ~n16498;
  assign n15662 = ~n15661 | ~n15660;
  assign n15167 = ~n15157 | ~n15156;
  assign n17020 = ~n17054 | ~n17019;
  assign n16776 = ~n16775 | ~n16774;
  assign n14777 = ~n14808 & ~n14769;
  assign n14709 = ~n14706 & ~n14705;
  assign n10736 = ~n10735 & ~n10734;
  assign n17117 = ~n10082 | ~n10081;
  assign n15946 = ~n15945 | ~n15944;
  assign n10059 = ~n10058 | ~n10057;
  assign n15110 = ~n15109 | ~n15108;
  assign n10170 = ~n10169 | ~n10168;
  assign n15820 = ~n15818 | ~n15817;
  assign n15623 = ~n15621 | ~n15791;
  assign n14992 = ~n14976 | ~n14975;
  assign n16403 = ~n16402 | ~n16401;
  assign n15877 = ~n15876 | ~n15875;
  assign n15569 = ~n15568 | ~n15567;
  assign n15257 = n14575 ^ n14574;
  assign n16775 = ~n16770 | ~n16769;
  assign n15661 = ~n15659 | ~n16500;
  assign n14937 = ~n14936 | ~n14935;
  assign n15070 = ~n15067 | ~n15066;
  assign n16401 = ~n16400 & ~n16399;
  assign n15157 = ~n15155 | ~n10774;
  assign n15686 = ~n15685 & ~n15684;
  assign n14765 = ~n14763 | ~n15800;
  assign n15702 = ~n15701 & ~n15700;
  assign n15705 = ~n15704 & ~n16436;
  assign n14575 = n11306 & n11046;
  assign n15645 = ~n16524 | ~n16853;
  assign n15876 = ~n16436 | ~n15867;
  assign n11301 = ~n11297 & ~n11298;
  assign n15817 = ~n15816 & ~n15815;
  assign n14929 = ~n14922 & ~n14921;
  assign n14706 = ~n14701 & ~n16498;
  assign n14762 = ~n14763 | ~n15804;
  assign n11268 = ~n11292 | ~n11290;
  assign n15109 = ~n15105 | ~n15832;
  assign n15424 = ~n15410 & ~n15609;
  assign n16020 = ~n15467 | ~n15466;
  assign n14922 = ~n14915 & ~n14914;
  assign n15410 = ~n15409 | ~n15791;
  assign n14469 = ~n14467 | ~n16514;
  assign n11288 = ~n11287 | ~n11286;
  assign n15471 = ~n15470 | ~n15469;
  assign n14466 = ~n14467 | ~n16510;
  assign n15943 = ~n15941 & ~n15940;
  assign n11292 = ~n11265 | ~n11264;
  assign n17050 = ~n16874 & ~n16873;
  assign n16808 = ~n16790 | ~n16789;
  assign n15685 = n10032 & n10031;
  assign n15180 = ~n15179 | ~n15178;
  assign n15036 = ~n15035 | ~n15034;
  assign n10685 = ~n10729 | ~n10644;
  assign n17024 = ~n15299 | ~n16863;
  assign n16436 = ~n16048;
  assign n15495 = ~n15494 | ~n15493;
  assign n15700 = ~n15699 | ~n15698;
  assign n11305 = ~n11304 | ~n11303;
  assign n16814 = ~n16788;
  assign n9998 = ~n9997 | ~n9996;
  assign n14752 = ~n14745 & ~n14744;
  assign n15542 = ~n15541 & ~n15540;
  assign n15341 = ~n15340 | ~n15339;
  assign n16400 = ~n16389 | ~n16388;
  assign n14390 = ~n14387 & ~n14386;
  assign n14915 = ~n14934 & ~n15218;
  assign n11044 = ~n11304;
  assign n15299 = ~n16857;
  assign n15179 = ~n15177 & ~n15176;
  assign n14759 = ~n14758 | ~n14935;
  assign n14938 = ~n14934 & ~n14933;
  assign n11286 = ~n11285 & ~n11284;
  assign n14973 = ~n14969 & ~n15738;
  assign n15494 = ~n15492 | ~n16500;
  assign n11183 = ~n11182 & ~n11181;
  assign n15035 = ~n15029 | ~n15832;
  assign n15699 = ~n15695 & ~n15694;
  assign n15326 = ~n15325 | ~n15324;
  assign n14697 = ~n14698 | ~n15804;
  assign n15590 = ~n15589 & ~n15588;
  assign n15316 = ~n15315 | ~n15314;
  assign n14700 = ~n14698 | ~n15800;
  assign n15559 = ~n15558 & ~n15557;
  assign n15189 = ~n15188 | ~n15187;
  assign n15565 = ~n15558 & ~n15468;
  assign n11006 = ~n10996 | ~n10995;
  assign n15245 = ~n15244 | ~n15243;
  assign n15561 = ~n16392 & ~n16393;
  assign n15695 = ~n16778 & ~n17126;
  assign n14554 = ~n14543 | ~n10132;
  assign n15066 = n15065 & n15064;
  assign n14464 = ~n14457 | ~n15335;
  assign n14197 = ~n14385;
  assign n14989 = ~n14988 | ~n14987;
  assign n15325 = ~n15323 | ~n15791;
  assign n11182 = ~n15244 & ~n14079;
  assign n15588 = ~n15587 | ~n15586;
  assign n15558 = ~n16392;
  assign n11128 = ~n11127 & ~n11126;
  assign n14745 = ~n14738 & ~n14737;
  assign n15464 = ~n16386;
  assign n15288 = ~n15287 | ~n15286;
  assign n15408 = ~n16778 | ~n15312;
  assign n15540 = ~n15539 | ~n15538;
  assign n15289 = ~n15284 & ~n15338;
  assign n11304 = ~n11037 | ~n11036;
  assign n15448 = ~n15447 & ~n15446;
  assign n15338 = ~n15468 | ~n16500;
  assign n11037 = ~n11034 | ~n11033;
  assign n14694 = ~n14693 | ~n14935;
  assign n14101 = ~n14098 & ~n14097;
  assign n14687 = ~n14682 & ~n14681;
  assign n15938 = ~n15531 | ~n16379;
  assign n14615 = ~n14613 | ~n15804;
  assign n11127 = ~n11116 & ~n15547;
  assign n15587 = ~n15584 & ~n15583;
  assign n15186 = ~n15173 | ~n15172;
  assign n14760 = ~n14757 & ~n14756;
  assign n14913 = ~n14909 | ~n10774;
  assign n14538 = ~n14535 & ~n14534;
  assign n15521 = ~n15520 & ~n15519;
  assign n14612 = ~n14613 | ~n15800;
  assign n16386 = ~n15531 | ~n15463;
  assign n14665 = n14661 & n14660;
  assign n15065 = ~n15063 | ~n15791;
  assign n10860 = ~n10850 | ~n10849;
  assign n14535 = ~n14526 & ~n17147;
  assign n15063 = ~n14984 & ~n14983;
  assign n14212 = ~n14209 | ~n14208;
  assign n14776 = ~n14775 | ~n14774;
  assign n15584 = ~n15581 | ~n15580;
  assign n15519 = ~n15518 | ~n15517;
  assign n16382 = ~n16378 | ~n16379;
  assign n16763 = ~n16761 & ~n16760;
  assign n14456 = n14446 & n14445;
  assign n16771 = ~n15697 | ~n15175;
  assign n16373 = ~n16365 & ~n16364;
  assign n15274 = ~n15934;
  assign n15531 = ~n16378;
  assign n15446 = ~n15445 | ~n15444;
  assign n14682 = ~n14676 & ~n14675;
  assign n14661 = ~n14658 | ~n14657;
  assign n15936 = ~n16378 | ~n15463;
  assign n14037 = ~n14095;
  assign n11034 = ~n10065 | ~n10064;
  assign n16378 = ~n11249 & ~n11248;
  assign n11031 = ~n11030 | ~n11029;
  assign n14609 = ~n14656 | ~n14935;
  assign n14126 = ~n14123 | ~n14122;
  assign n15151 = ~n15150 & ~n15149;
  assign n14488 = ~n14489 | ~n15804;
  assign n14491 = ~n14489 | ~n15800;
  assign n15517 = ~n15516 & ~n15515;
  assign n15312 = ~n15579 & ~n15171;
  assign n14209 = ~n14203 | ~n15335;
  assign n15175 = ~n15579;
  assign n13949 = ~n13946 & ~n13945;
  assign n17051 = ~n15509 | ~n15579;
  assign n15934 = ~n16362 & ~n16367;
  assign n10987 = ~n10986 | ~n10985;
  assign n14987 = ~n14986 & ~n14985;
  assign n15283 = ~n16362 & ~n11177;
  assign n16760 = ~n16759 & ~n16758;
  assign n14775 = ~n14771 | ~n15832;
  assign n13942 = ~n13940 & ~n13939;
  assign n14736 = ~n14732 | ~n10774;
  assign n15240 = ~n15239 & ~n15238;
  assign n14695 = ~n14692 & ~n14691;
  assign n16359 = ~n16346 & ~n16345;
  assign n11160 = ~n15930;
  assign n15239 = ~n15237 | ~n15236;
  assign n16865 = ~n15511 & ~n15159;
  assign n15128 = ~n15127 | ~n15126;
  assign n14692 = ~n14674 | ~n14673;
  assign n14658 = ~n14654 & ~n14653;
  assign n14504 = ~n14501 & ~n14500;
  assign n14123 = ~n14121 & ~n14120;
  assign n16362 = ~n16366;
  assign n14921 = ~n14920 | ~n14919;
  assign n14525 = ~n9722 | ~n9721;
  assign n16342 = ~n16332 | ~n16331;
  assign n10062 = ~n10046 & ~n10045;
  assign n14610 = ~n14654 & ~n14603;
  assign n11005 = ~n11004 & ~n11003;
  assign n14113 = ~n14110 | ~n14109;
  assign n15149 = ~n15148 | ~n15147;
  assign n16768 = ~n16762;
  assign n10023 = ~n13943;
  assign n15268 = ~n16366 | ~n16367;
  assign n10684 = ~n10683 & ~n10682;
  assign n14062 = ~n14050 & ~n14049;
  assign n15932 = ~n16366 & ~n16363;
  assign n15120 = ~n15119 | ~n15118;
  assign n9940 = ~n9939;
  assign n11161 = ~n16358;
  assign n14110 = ~n14074 & ~n14073;
  assign n10683 = ~n10672 & ~n15547;
  assign n13810 = ~n13808 & ~n13807;
  assign n15022 = ~n15021 & ~n15020;
  assign n15161 = ~n15160 & ~n15159;
  assign n14443 = ~n14436 | ~n14435;
  assign n14485 = ~n14502 | ~n14935;
  assign n15227 = ~n9937 & ~n9936;
  assign n14109 = ~n14108 & ~n14107;
  assign n15118 = ~n15117 & ~n15116;
  assign n10875 = ~n10874 | ~n10873;
  assign n16358 = ~n16348 & ~n16347;
  assign n14933 = ~n14932 | ~n14931;
  assign n14195 = ~n14194 & ~n14193;
  assign n14654 = ~n14597 | ~n14596;
  assign n15511 = ~n15160;
  assign n14121 = ~n14116 & ~n15657;
  assign n14463 = ~n14462 & ~n14461;
  assign n14049 = ~n15563 & ~n14116;
  assign n14320 = ~n14317 & ~n14316;
  assign n15236 = ~n15235 & ~n15234;
  assign n14092 = ~n14091 & ~n14090;
  assign n14501 = ~n14494 & ~n14493;
  assign n16762 = ~n15582 & ~n15160;
  assign n14674 = ~n14670 | ~n10774;
  assign n9909 = ~n9908 & ~n15078;
  assign n15930 = ~n16348 | ~n15030;
  assign n15097 = ~n15096 & ~n15095;
  assign n15127 = ~n15125 | ~n16500;
  assign n10980 = ~n14436 | ~n14434;
  assign n11115 = ~n16010;
  assign n14194 = ~n14186 & ~n17147;
  assign n11113 = ~n11112 & ~n11111;
  assign n13937 = ~n13931 & ~n13930;
  assign n11164 = ~n13805 & ~n9036;
  assign n15020 = ~n15019 | ~n15018;
  assign n9937 = ~n15231 & ~n9934;
  assign n10859 = ~n10858 & ~n10857;
  assign n15046 = ~n15045 | ~n15044;
  assign n11147 = ~n15926;
  assign n16351 = ~n16336 & ~n16335;
  assign n9908 = ~n15081 & ~n15080;
  assign n14021 = ~n14018 | ~n14017;
  assign n14108 = ~n14103 & ~n16498;
  assign n15095 = ~n15094 | ~n15093;
  assign n14462 = ~n11002 | ~n11001;
  assign n14597 = ~n14593 | ~n10774;
  assign n16754 = ~n16869;
  assign n15054 = ~n15053 | ~n15052;
  assign n16348 = ~n15115;
  assign n14074 = ~n14067 | ~n14066;
  assign n15235 = ~n15231 & ~n17126;
  assign n16747 = ~n16737 & ~n16736;
  assign n14317 = ~n14310 & ~n14309;
  assign n10874 = ~n10866 | ~n10132;
  assign n14486 = ~n14492 & ~n14479;
  assign n9911 = ~n15081 | ~n15080;
  assign n14435 = ~n14434 | ~n14433;
  assign n14756 = ~n14755 | ~n14754;
  assign n11137 = ~n11136 & ~n11135;
  assign n14263 = ~n14260 & ~n14259;
  assign n14287 = ~n14318 | ~n14935;
  assign n14181 = ~n14179 & ~n14178;
  assign n11002 = ~n10998 | ~n15832;
  assign n15053 = ~n15051 | ~n16500;
  assign n14001 = ~n14010 & ~n13999;
  assign n15076 = ~n14945 | ~n14944;
  assign n14008 = ~n14007 & ~n14006;
  assign n11146 = ~n15924;
  assign n13707 = ~n13705 & ~n17084;
  assign n13712 = ~n13710 & ~n16492;
  assign n14103 = ~n14102;
  assign n11234 = ~n15010;
  assign n14982 = ~n14981 & ~n14980;
  assign n14492 = ~n14475 | ~n14474;
  assign n15094 = ~n15092 & ~n15091;
  assign n14208 = ~n14207 & ~n14206;
  assign n14904 = ~n14903 & ~n14902;
  assign n15115 = ~n11151 & ~n11150;
  assign n16869 = ~n14981 & ~n14906;
  assign n14288 = ~n14308 & ~n14278;
  assign n14381 = ~n14378 | ~n14377;
  assign n16737 = ~n16552 & ~n16551;
  assign n14017 = ~n14016 & ~n14015;
  assign n13921 = ~n13918 | ~n13917;
  assign n16010 = ~n11107 & ~n11106;
  assign n10969 = ~n10954 | ~n10953;
  assign n13805 = ~n10011 ^ n10010;
  assign n14980 = ~n15087 | ~n14916;
  assign n14981 = ~n9922 | ~n9921;
  assign n16741 = ~n14924 | ~n15087;
  assign n14945 = ~n15078;
  assign n14377 = ~n14376 & ~n14375;
  assign n14239 = ~n14398 | ~n14238;
  assign n14957 = ~n14956 & ~n14955;
  assign n14401 = ~n14398 | ~n14397;
  assign n14308 = ~n14274 | ~n14273;
  assign n15000 = ~n14999 & ~n14998;
  assign n9951 = ~n13708;
  assign n14207 = ~n10856 | ~n10855;
  assign n14369 = ~n14368 & ~n14367;
  assign n14475 = ~n14471 | ~n10774;
  assign n16552 = ~n16547 & ~n16546;
  assign n14902 = ~n14901 | ~n14900;
  assign n14378 = ~n14358 & ~n14357;
  assign n14728 = ~n14727 & ~n14726;
  assign n16328 = ~n16319 & ~n16318;
  assign n9903 = ~n9902 | ~n9901;
  assign n10011 = ~n9984 | ~n9983;
  assign n14010 = ~n13996 | ~n13995;
  assign n14178 = ~n14177 | ~n14176;
  assign n14016 = ~n14011 & ~n16498;
  assign n14259 = ~n14258 | ~n14257;
  assign n13918 = ~n13927;
  assign n14592 = ~n14668 & ~n14591;
  assign n15087 = ~n16738;
  assign n14305 = ~n14302 | ~n14301;
  assign n14161 = ~n14302 | ~n14160;
  assign n13927 = ~n13910 | ~n13909;
  assign n13708 = n9981 ^ n9950;
  assign n14955 = ~n14954 | ~n14953;
  assign n16317 = ~n16301 | ~n16300;
  assign n16546 = ~n16732 & ~n16545;
  assign n14357 = ~n14371 & ~n15404;
  assign n14398 = ~n14235 & ~n14234;
  assign n14726 = ~n14725 | ~n14724;
  assign n13995 = ~n14005 | ~n10644;
  assign n14944 = ~n9907 | ~n9906;
  assign n13827 = ~n13826 & ~n13825;
  assign n10856 = ~n10852 | ~n15832;
  assign n14847 = ~n14846 | ~n14845;
  assign n14786 = ~n14785 | ~n14784;
  assign n14812 = ~n14811 | ~n14810;
  assign n14274 = ~n14270 | ~n10774;
  assign n13899 = ~n13896 | ~n13895;
  assign n14122 = ~n14058 & ~n14057;
  assign n15078 = ~n9907 & ~n9906;
  assign n14358 = ~n14353 | ~n14352;
  assign n16316 = ~n16298 & ~n16299;
  assign n14691 = ~n14690 | ~n14689;
  assign n14767 = ~n15916;
  assign n11094 = ~n16298 | ~n16299;
  assign n14058 = ~n14054 & ~n15547;
  assign n16732 = ~n16542 | ~n16541;
  assign n13981 = ~n13978 & ~n13977;
  assign n13895 = n13894 & n13893;
  assign n14301 = ~n14300 & ~n14299;
  assign n13826 = ~n13817 & ~n17147;
  assign n9920 = ~n13508;
  assign n13996 = ~n13992 & ~n13991;
  assign n13680 = ~n13677 | ~n13676;
  assign n16321 = ~n14997;
  assign n14270 = ~n14269 | ~n14470;
  assign n14034 = ~n14031 | ~n14030;
  assign n14175 = ~n14174 & ~n14173;
  assign n14953 = ~n14952 & ~n14951;
  assign n13917 = ~n13916 & ~n13915;
  assign n14715 = ~n11223 | ~n11224;
  assign n13910 = ~n13906 & ~n13905;
  assign n11226 = ~n11223;
  assign n14302 = ~n14157 & ~n14156;
  assign n14163 = ~n14142 & ~n14141;
  assign n14603 = ~n14651 | ~n14602;
  assign n11145 = ~n13508 & ~n9036;
  assign n14234 = ~n14233 | ~n14232;
  assign n16738 = ~n9900 | ~n9899;
  assign n11141 = ~n14997 | ~n15031;
  assign n14746 = ~n14948 | ~n14850;
  assign n14255 = ~n14250 & ~n14249;
  assign n9947 = ~n9944 | ~n9943;
  assign n14030 = ~n14029 & ~n14028;
  assign n14157 = ~n14155 | ~n14154;
  assign n14845 = ~n9857 | ~n9856;
  assign n14233 = ~n14231 & ~n14230;
  assign n14353 = ~n14349 | ~n10774;
  assign n14651 = ~n14601 | ~n14739;
  assign n13894 = ~n13732 & ~n13731;
  assign n13677 = ~n13628 & ~n13627;
  assign n16292 = ~n16061 & ~n16060;
  assign n13978 = ~n13972 & ~n15218;
  assign n16879 = ~n14948 | ~n15088;
  assign n13992 = ~n13987 & ~n13986;
  assign n9906 = ~n9882 | ~n9881;
  assign n9880 = ~n9879 | ~n9878;
  assign n13817 = ~n13816 & ~n13815;
  assign n11174 = ~n16302 | ~n14783;
  assign n14156 = ~n14294 & ~n15404;
  assign n16298 = ~n16302;
  assign n16290 = ~n16067 & ~n16066;
  assign n13676 = ~n13675 & ~n13674;
  assign n14948 = ~n14748;
  assign n13896 = ~n13892 & ~n13891;
  assign n13972 = ~n14026 & ~n13971;
  assign n14539 = ~n9794 | ~n9793;
  assign n10849 = ~n10848 & ~n10847;
  assign n14916 = ~n14748 & ~n14739;
  assign n14053 = ~n14052 | ~n14051;
  assign n14705 = ~n14704 | ~n14703;
  assign n13334 = ~n11096;
  assign n14155 = ~n14150 | ~n10774;
  assign n11098 = ~n11096 & ~n9036;
  assign n11221 = ~n11220 & ~n11219;
  assign n14479 = ~n14478 | ~n14477;
  assign n14071 = ~n14069 | ~n14068;
  assign n14608 = ~n16878 | ~n14667;
  assign n14889 = ~n14886 & ~n14885;
  assign n14069 = ~n13985 | ~n13984;
  assign n13909 = ~n13908 | ~n15832;
  assign n9853 = ~n9852 | ~n9851;
  assign n14739 = ~n16530 | ~n14600;
  assign n9858 = ~n9855 | ~n9854;
  assign n11220 = ~n11218;
  assign n14026 = ~n13959 | ~n13958;
  assign n16887 = ~n14667 | ~n14666;
  assign n14461 = ~n14460 | ~n14459;
  assign n16878 = ~n16530 | ~n16534;
  assign n11085 = ~n11084 | ~n15913;
  assign n14206 = ~n14205 | ~n14204;
  assign n14748 = ~n9869 | ~n9868;
  assign n10995 = ~n10994 & ~n10993;
  assign n14397 = ~n14396 & ~n14395;
  assign n16537 = ~n16530 | ~n16531;
  assign n10602 = ~n16003 | ~n16051;
  assign n14348 = ~n14346 | ~n14345;
  assign n14540 = ~n9791 | ~n9792;
  assign n14149 = ~n14265 | ~n16672;
  assign n14484 = ~n14591 & ~n16881;
  assign n13667 = ~n13664 | ~n13663;
  assign n13844 = ~n13841 & ~n13840;
  assign n14515 = ~n11216 | ~n11215;
  assign n11091 = ~n13155 | ~n11089;
  assign n14844 = ~n14841 & ~n14840;
  assign n11087 = ~n15914 | ~n14506;
  assign n14667 = ~n16548 | ~n16531;
  assign n13958 = ~n13957 | ~n14225;
  assign n14783 = ~n15914 & ~n11134;
  assign n14885 = ~n14884 | ~n14883;
  assign n14228 = ~n14227 & ~n14226;
  assign n13670 = ~n13620 | ~n13619;
  assign n14235 = ~n14391 & ~n15404;
  assign n14600 = ~n14598 & ~n14797;
  assign n13749 = ~n13746 | ~n13745;
  assign n14883 = ~n14882 | ~n14881;
  assign n14840 = ~n14839 | ~n14838;
  assign n14480 = ~n16712 | ~n16713;
  assign n13500 = ~n13497 | ~n13496;
  assign n14516 = ~n11213 | ~n11214;
  assign n14031 = ~n14024 | ~n14935;
  assign n13745 = ~n13744 & ~n13743;
  assign n16540 = ~n16728 | ~n16544;
  assign n14792 = ~n9824 | ~n9823;
  assign n14227 = ~n14225;
  assign n14267 = ~n16885;
  assign n9788 = ~n9787 | ~n9786;
  assign n13664 = ~n13601 & ~n13600;
  assign n14524 = ~n14523 & ~n14522;
  assign n14598 = ~n16712 | ~n14476;
  assign n14573 = ~n14571 & ~n14570;
  assign n13719 = ~n13616 & ~n13614;
  assign n9792 = ~n9790 | ~n9789;
  assign n9822 = ~n9821 | ~n9820;
  assign n10627 = ~n14510 | ~n11788;
  assign n13497 = ~n13494 & ~n13493;
  assign n14024 = ~n14131 | ~n13967;
  assign n14523 = ~n9759 & ~n9758;
  assign n13737 = ~n13702 | ~n13701;
  assign n13802 = ~n13832 | ~n13799;
  assign n10662 = ~n13729 & ~n15899;
  assign n14570 = ~n14569 | ~n14568;
  assign n16885 = ~n16716 | ~n16713;
  assign n16880 = ~n16716 & ~n16713;
  assign n13616 = ~n13618 & ~n16220;
  assign n13955 = ~n13956 & ~n16996;
  assign n9893 = ~n9865 | ~n9864;
  assign n14839 = ~n14851 & ~n14835;
  assign n14666 = ~n14797 | ~n16544;
  assign n13404 = ~n13401 | ~n13400;
  assign n16881 = ~n14797 & ~n16544;
  assign n15881 = ~n14510 & ~n14642;
  assign n10731 = ~n14510;
  assign n14522 = ~n9756 & ~n9757;
  assign n13401 = ~n13398 & ~n13397;
  assign n14841 = ~n14826 & ~n14825;
  assign n9759 = ~n9756;
  assign n13663 = ~n13662 & ~n13661;
  assign n16056 = ~n16053;
  assign n14343 = ~n14341 & ~n14340;
  assign n14879 = ~n14878 & ~n14877;
  assign n14355 = ~n14354;
  assign n13701 = ~n13700 & ~n13699;
  assign n14568 = ~n14567 | ~n14882;
  assign n14835 = ~n14834 & ~n14833;
  assign n14884 = ~n14873 | ~n11932;
  assign n13417 = ~n13414 | ~n13413;
  assign n11022 = ~n11021 | ~n11020;
  assign n14354 = ~n14347 | ~n16884;
  assign n14878 = ~n14875 & ~n14874;
  assign n13832 = ~n13787 & ~n13786;
  assign n10661 = ~n13625 & ~n15988;
  assign n11021 = ~n14439 | ~n11016;
  assign n13396 = ~n13183 & ~n13182;
  assign n13830 = ~n13791 & ~n13790;
  assign n11011 = ~n14440 | ~n11010;
  assign n16699 = ~n16684 & ~n16683;
  assign n14283 = ~n16687 | ~n16689;
  assign n13414 = ~n13358 & ~n13357;
  assign n10590 = ~n12680 & ~n9036;
  assign n9753 = ~n9751 | ~n9750;
  assign n9834 = ~n9831 | ~n9830;
  assign n14831 = ~n14830 | ~n14829;
  assign n16940 = ~n17002 & ~n14344;
  assign n14871 = ~n14870 & ~n14869;
  assign n9757 = ~n9755 | ~n9754;
  assign n14279 = ~n17000;
  assign n14440 = ~n11013 | ~n14437;
  assign n14476 = ~n16692 & ~n14362;
  assign n14870 = ~n14868 & ~n14867;
  assign n14822 = ~n14633 | ~n14632;
  assign n14439 = ~n11013;
  assign n13960 = ~n13788 | ~n13599;
  assign n9831 = ~n9800 | ~n9799;
  assign n9720 = ~n10863;
  assign n14830 = ~n14621 | ~n14620;
  assign n16279 = ~n15882;
  assign n16884 = ~n16692 | ~n16689;
  assign n14565 = ~n14563 & ~n14562;
  assign n17002 = ~n16692 & ~n16689;
  assign n11016 = ~n11015 | ~n14437;
  assign n16272 = ~n14447 | ~n16277;
  assign n13244 = ~n13232 & ~n13231;
  assign n15905 = ~n15996 & ~n16251;
  assign n15882 = ~n14447 & ~n16277;
  assign n9629 = ~n13847 & ~n13845;
  assign n14106 = ~n14083 & ~n14082;
  assign n14620 = ~n14618 | ~n14617;
  assign n11020 = ~n11019 | ~n11018;
  assign n10844 = ~n14447 | ~n14082;
  assign n10577 = ~n14447 | ~n16285;
  assign n14632 = ~n14629 | ~n14628;
  assign n14560 = ~n14558 & ~n14557;
  assign n10665 = ~n14104 | ~n16265;
  assign n14362 = ~n16700 | ~n14275;
  assign n14129 = ~n14264;
  assign n14617 = ~n14332 | ~n14331;
  assign n14628 = ~n14324 | ~n14323;
  assign n13847 = ~n9630 | ~n9626;
  assign n9738 = ~n9731 | ~n15212;
  assign n9715 = ~n9714 | ~n9713;
  assign n16922 = n14264 & n16672;
  assign n10862 = n9718 & n9717;
  assign n10562 = ~n16270;
  assign n9668 = ~n9667;
  assign n16931 = ~n14226 & ~n16680;
  assign n9731 = ~n12427;
  assign n10978 = ~n10977 | ~n10976;
  assign n16270 = ~n16266 & ~n16265;
  assign n14323 = ~n14322 | ~n14321;
  assign n13597 = ~n13593 | ~n13592;
  assign n9626 = ~n9625 | ~n9624;
  assign n14331 = ~n14330 | ~n14329;
  assign n14082 = ~n16266 & ~n14080;
  assign n14264 = ~n14296 | ~n16701;
  assign n14344 = ~n14296 & ~n16701;
  assign n10570 = ~n12427 & ~n9036;
  assign n16700 = ~n14296;
  assign n16998 = ~n14215 | ~n16672;
  assign n10666 = ~n16266 | ~n10956;
  assign n9663 = ~n9662 | ~n9661;
  assign n13593 = ~n13589 | ~n13588;
  assign n9630 = ~n9622 | ~n9623;
  assign n14132 = ~n14217 | ~n14151;
  assign n14226 = ~n14148 | ~n14147;
  assign n10977 = ~n10974;
  assign n14321 = ~n13777 | ~n13776;
  assign n14329 = ~n13764 | ~n13763;
  assign n13866 = ~P2_REG2_REG_15__SCAN_IN & ~n13865;
  assign n14080 = ~n16243 | ~n14002;
  assign n14184 = n9665 & n9664;
  assign n16680 = ~n16657 & ~n14151;
  assign n13548 = ~n10835 & ~n13387;
  assign n13763 = ~n13761 | ~n13760;
  assign n10664 = ~n16247 | ~n16244;
  assign n13776 = ~n13773 | ~n13772;
  assign n15994 = ~n16251 & ~n16252;
  assign n13867 = ~n13874 & ~n13864;
  assign n14275 = ~n16657 & ~n14236;
  assign n10948 = ~n14251 & ~n14247;
  assign n9700 = ~n12295 | ~n15212;
  assign n13772 = ~P1_REG2_REG_15__SCAN_IN | ~n13455;
  assign n16919 = n16671 & n16661;
  assign n9619 = ~n9618 | ~n9617;
  assign n13876 = ~P2_REG1_REG_15__SCAN_IN & ~n13875;
  assign n13225 = ~n13222 | ~n13221;
  assign n14251 = ~n10950 & ~n10949;
  assign n14252 = ~n10950 | ~n10949;
  assign n13845 = ~n9628 & ~n9627;
  assign n9623 = ~n9621 | ~n9620;
  assign n10835 = ~n13386 & ~n13388;
  assign n13846 = ~n9628 | ~n9627;
  assign n10529 = ~n10528 | ~n14167;
  assign n13760 = ~P1_REG1_REG_15__SCAN_IN | ~n13462;
  assign n14130 = ~n14159 | ~n14146;
  assign n13877 = ~n13874 & ~n13873;
  assign n9724 = ~n9675 | ~n9674;
  assign n15992 = ~n13718 | ~n13717;
  assign n10537 = ~n12146 | ~n10310;
  assign n14002 = ~n13911 & ~n14261;
  assign n16252 = ~n14261 & ~n14167;
  assign n13982 = ~n14261 | ~n14167;
  assign n13388 = ~n10834 & ~n13196;
  assign n13538 = ~n13537 & ~n13536;
  assign n14159 = ~n16668;
  assign n9650 = ~n12146 | ~n15212;
  assign n9591 = ~n9590 | ~n9589;
  assign n13759 = ~n13460 | ~n13459;
  assign n10834 = ~n13195 & ~n13197;
  assign n9627 = ~n9593 | ~n9592;
  assign n13963 = ~n13962 | ~n13961;
  assign n16643 = ~n16661;
  assign n13537 = ~n12923 & ~n12922;
  assign n14171 = ~n10947 | ~n10946;
  assign n10511 = ~n16225 | ~n16226;
  assign n13106 = ~n13370 | ~n13103;
  assign n14247 = ~n10947 & ~n10946;
  assign n13566 = ~n9557 | ~n9556;
  assign n13532 = ~n13531 & ~n13530;
  assign n12922 = ~n12921 & ~n12920;
  assign n14144 = ~n13973 & ~n13961;
  assign n15839 = ~n15838 & ~n15837;
  assign n16225 = ~n16229;
  assign n13720 = ~n13637 & ~n16188;
  assign n13565 = ~n9555 | ~n9554;
  assign n16661 = ~n13973 | ~n13961;
  assign n14158 = ~n13974 & ~n13973;
  assign n13459 = ~n12989 | ~n12988;
  assign n9606 = ~n12077 | ~n15212;
  assign n13717 = ~n16229 | ~n16226;
  assign n13453 = ~n13452 & ~n13451;
  assign n15902 = ~n16229 & ~n16226;
  assign n12988 = ~n12985 | ~n12984;
  assign n10653 = ~n12869 & ~n16110;
  assign n10833 = ~n12834 & ~n12836;
  assign n15598 = ~n15597 & ~n15596;
  assign n13518 = ~n10938 | ~n10937;
  assign n13645 = ~n10944 | ~n10943;
  assign n15716 = ~n15715 & ~n15714;
  assign n15988 = ~n13614 & ~n16220;
  assign n13451 = ~n12977 | ~n12976;
  assign n15989 = ~n13689 & ~n15895;
  assign n9469 = ~n9468 | ~n9467;
  assign n10468 = ~n16175;
  assign n12976 = ~n12483 | ~n12482;
  assign n9556 = ~n9553 | ~n9552;
  assign n13614 = ~n16203 & ~n16192;
  assign n9503 = ~n9502 | ~n9501;
  assign n15986 = ~n13311 & ~n13310;
  assign n12584 = ~n12583 & ~n12582;
  assign n15834 = ~n15868;
  assign n12915 = ~n12914 & ~n12913;
  assign n9579 = ~n11995 | ~n15212;
  assign n13517 = ~n10935 | ~n10936;
  assign n9551 = ~n9550 | ~n9549;
  assign n13688 = ~n16176 & ~n13309;
  assign n13554 = ~n10933 & ~n10932;
  assign n9633 = ~n9598 | ~n9597;
  assign n10938 = ~n10935;
  assign n13974 = ~n13793 | ~n13792;
  assign n12984 = ~n12474 | ~n12473;
  assign n13646 = ~n10941 | ~n10942;
  assign n13485 = ~n9505 | ~n9504;
  assign n16637 = ~n13792 | ~n13818;
  assign n16934 = ~n13349 | ~n16616;
  assign n16987 = ~n13588 | ~n13590;
  assign n13595 = ~n13611;
  assign n15895 = ~n16205 & ~n13642;
  assign n16914 = ~n13837 | ~n13598;
  assign n12583 = ~n12310 & ~n12309;
  assign n15752 = ~n17112;
  assign n10934 = ~n10933;
  assign n13309 = ~n13185 | ~n13184;
  assign n10832 = ~n12571 & ~n12573;
  assign n12483 = ~n12481 & ~n12480;
  assign n10392 = ~n15981;
  assign n12474 = ~n12472 & ~n12471;
  assign n16220 = ~n16188 & ~n16189;
  assign n16203 = ~n16188;
  assign n16175 = ~n16205 & ~n16195;
  assign n10932 = ~n10931 & ~n10930;
  assign n9466 = ~n9463 | ~n9462;
  assign n12472 = ~n12470 & ~n12469;
  assign n9461 = ~n9460 | ~n9459;
  assign n15563 = ~n14047;
  assign n15890 = ~n16199 | ~n16177;
  assign n13022 = ~n10916 | ~n10915;
  assign n13203 = ~n10921 | ~n10920;
  assign n12309 = ~n12308 & ~n12307;
  assign n10933 = ~n10928 & ~n10929;
  assign n10445 = ~n16199 | ~n16209;
  assign n12578 = ~n12577 & ~n12576;
  assign n11316 = n11315 & n11314;
  assign n12480 = ~n12479 & ~n12478;
  assign n13185 = ~n13266 & ~n13443;
  assign n13173 = ~n15984;
  assign n15281 = ~n15280 & ~n15279;
  assign n10831 = ~n12319 & ~n12321;
  assign n9486 = ~n11831 | ~n15212;
  assign n13266 = ~n13003 | ~n13032;
  assign n15566 = ~n15848;
  assign n9539 = ~n11822 | ~n15212;
  assign n14047 = ~n15845 | ~n10841;
  assign n15984 = ~n10656 | ~n10657;
  assign n12469 = ~n12102 | ~n12101;
  assign n15486 = ~n16405 & ~n15713;
  assign n12577 = ~n12304 & ~n12303;
  assign n12308 = ~n12085 & ~n12084;
  assign n12479 = ~n12109 & ~n12108;
  assign n15888 = ~n16176 | ~n16209;
  assign n15865 = ~n15530;
  assign n13295 = ~n10926 | ~n10925;
  assign n12372 = ~n10786 | ~n10785;
  assign n10456 = ~n11831 | ~n10310;
  assign n10475 = ~n11822 | ~n10310;
  assign n10163 = ~n10159 & ~n10158;
  assign n12101 = ~n11978 | ~n11977;
  assign n12108 = ~n12107 & ~n12106;
  assign n9561 = ~n9559;
  assign n15848 = ~n15720 | ~n15285;
  assign n15847 = ~n13071;
  assign n10965 = ~n10964 | ~n15285;
  assign n10159 = ~n12041 & ~n17128;
  assign n10078 = ~n16853 | ~n17111;
  assign n13294 = ~n10923 | ~n10924;
  assign n11329 = ~n9035 | ~n11327;
  assign n12084 = ~n12083 & ~n12082;
  assign n13003 = ~n12873 & ~n12876;
  assign n15724 = ~n11327 & ~n11313;
  assign n16606 = ~n13116 & ~n16899;
  assign n16405 = ~n15704;
  assign n12303 = ~n12302 & ~n12301;
  assign n11225 = ~n11224;
  assign n16393 = ~n15557;
  assign n16367 = ~n16363;
  assign n16265 = ~n10956;
  assign n16853 = ~n10077 | ~n10076;
  assign n9476 = ~n9473 | ~n9512;
  assign n16135 = ~n13265 | ~n13288;
  assign n10376 = ~n13020 | ~n13251;
  assign n9450 = ~n11778 | ~n15212;
  assign n12646 = ~n13251;
  assign n15030 = ~n16347;
  assign n15031 = ~n16322;
  assign n16248 = ~n16244;
  assign n16609 = ~n13223 & ~n13366;
  assign n10830 = ~n12138 & ~n12140;
  assign n12106 = ~n11972 | ~n11971;
  assign n11977 = ~n11976 | ~n11975;
  assign n10882 = ~n12334 & ~n10881;
  assign n13988 = ~n14167;
  assign n16338 = ~n16334;
  assign n15869 = ~n15535;
  assign n16054 = ~n16051;
  assign n12083 = ~n11966 & ~n11965;
  assign n12302 = ~n12092 & ~n12091;
  assign n16379 = ~n15463;
  assign n15913 = ~n14506;
  assign n10657 = ~n16160 | ~n13317;
  assign n14642 = ~n11788;
  assign n16164 = ~n16160 & ~n16161;
  assign n15557 = ~n11263 | ~n11262;
  assign n11971 = ~n11762 | ~n11761;
  assign n11975 = ~n11751 | ~n11750;
  assign n16160 = ~n10410 | ~n10409;
  assign n11788 = ~n10624 | ~n10623;
  assign n11278 = ~n15564 | ~n9035;
  assign n10963 = ~n10960 | ~n11612;
  assign n12091 = ~n12090 & ~n12089;
  assign n11965 = ~n11964 & ~n11963;
  assign n16209 = ~n10444 & ~n10443;
  assign n16816 = ~n16787;
  assign n10156 = ~n10154 | ~n10153;
  assign n12334 = ~n10960 & ~n12004;
  assign n10956 = ~n10561 & ~n10560;
  assign n16347 = ~n11158 | ~n11157;
  assign n15452 = ~n15962 & ~n15835;
  assign n16511 = ~n12021 | ~n12009;
  assign n11313 = ~P2_REG3_REG_28__SCAN_IN & ~n11312;
  assign n16516 = ~n12021 | ~n12020;
  assign n11262 = n11261 & n11260;
  assign n9473 = ~n9472 | ~n9471;
  assign n17126 = ~n15578;
  assign n10623 = n10622 & n10621;
  assign n10829 = ~n12000 & ~n12002;
  assign n11170 = n11169 & n11168;
  assign n11104 = n11103 & n11102;
  assign n10678 = n10677 & n10676;
  assign n16787 = ~n10041 | ~n10040;
  assign n11260 = ~n9035 | ~n15473;
  assign n10728 = ~n12008 & ~n10727;
  assign n10598 = n10597 & n10596;
  assign n11122 = n11121 & n11120;
  assign n11196 = n11192 & n11191;
  assign n11312 = n11311 & P2_REG3_REG_27__SCAN_IN;
  assign n12090 = ~n11956 & ~n11955;
  assign n11964 = ~n11943 | ~n12123;
  assign n11157 = n11156 & n11155;
  assign n10252 = n10251 & n10250;
  assign n15689 = ~n17132;
  assign n13443 = ~n13265;
  assign n10345 = n10341 & n10340;
  assign n15762 = ~n15174;
  assign n10483 = ~n10482 | ~n10481;
  assign n11751 = ~n11748 & ~n11747;
  assign n10073 = ~n12041 & ~n15610;
  assign n11762 = ~n11758 & ~n11757;
  assign n10466 = ~n10462 | ~n10461;
  assign n16087 = ~n16069 | ~n16068;
  assign n10544 = ~n10540 | ~n10539;
  assign n11748 = ~n11745 & ~n11744;
  assign n11758 = ~n11755 & ~n11754;
  assign n16781 = ~n10009 | ~n10008;
  assign n15509 = ~n15697;
  assign n9379 = ~n9372 | ~n15212;
  assign n15758 = ~n15745 | ~n14655;
  assign n12002 = ~n10828 & ~n11813;
  assign n13020 = ~n13032;
  assign n10250 = ~n9035 | ~n14640;
  assign n10676 = ~n9035 | ~n14780;
  assign n11103 = ~n9035 | ~n14895;
  assign n11156 = ~n9035 | ~n15142;
  assign n11169 = ~n9035 | ~n15439;
  assign n11277 = ~n11276 & ~n11275;
  assign n11311 = ~n11270 & ~n11279;
  assign n16452 = ~n11794 | ~n11793;
  assign n15967 = ~n11809 | ~n11808;
  assign n10727 = ~n11464 | ~n10726;
  assign n17147 = ~n10132;
  assign n9990 = ~n15697 | ~n17111;
  assign n15578 = ~n10136 | ~n15766;
  assign n10253 = n10243 & n10242;
  assign n11745 = ~n11719 | ~n11718;
  assign n10828 = ~n11812 & ~n11814;
  assign n9350 = ~n9349 | ~n9348;
  assign n11755 = ~n11714 & ~n11713;
  assign n11195 = n11194 & n11193;
  assign n10525 = ~n10524 | ~n10523;
  assign n10508 = ~n10507 | ~n10506;
  assign n13317 = ~n10418 & ~n10417;
  assign n11270 = ~n11259 | ~P2_REG3_REG_25__SCAN_IN;
  assign n12009 = ~n12020;
  assign n12005 = ~n16486 & ~n12004;
  assign n15745 = ~n10766 | ~n15766;
  assign n15725 = ~n15850;
  assign n11954 = ~n11931 | ~n12129;
  assign n10751 = ~n10140 & ~n10139;
  assign n9208 = ~n9207 & ~n9206;
  assign n12539 = ~n9177 & ~n9176;
  assign n12120 = ~n11942 & ~n11941;
  assign n11259 = n11190 & P2_REG3_REG_24__SCAN_IN;
  assign n16544 = ~n14605;
  assign n10287 = n10286 & n10285;
  assign n11719 = ~n11686 | ~n11685;
  assign n11714 = ~n11696 & ~n11695;
  assign n9309 = ~n9293 | ~n15212;
  assign n10474 = n10473 & n10472;
  assign n10553 = n10552 & n10551;
  assign n10569 = ~n10568 | ~n10567;
  assign n10536 = n10535 & n10534;
  assign n10070 = ~n10034 & ~n15690;
  assign n9040 = ~n10412;
  assign n10589 = ~n10588 | ~n10587;
  assign n11814 = ~n10827 & ~n10826;
  assign n14906 = ~n15512;
  assign n9274 = ~n9273 & ~n9272;
  assign n10147 = ~n10749 & ~n11369;
  assign n10315 = ~n9036 & ~n11386;
  assign n15512 = ~n9930 | ~n9929;
  assign n10497 = ~n10496 & ~n10495;
  assign n13366 = ~n13228;
  assign n11686 = ~n11683 | ~n11682;
  assign n10034 = ~n10002 | ~P1_REG3_REG_24__SCAN_IN;
  assign n10616 = ~n10615 & ~n10614;
  assign n10720 = ~P2_D_REG_1__SCAN_IN & ~n11611;
  assign n10235 = ~n10234 & ~n10233;
  assign n16534 = ~n9850 | ~n9849;
  assign n10455 = ~n10454 & ~n10453;
  assign n10430 = ~n10429 & ~n10428;
  assign n15806 = ~n12182 | ~n12181;
  assign n10409 = ~n10408 & ~n10407;
  assign n15801 = ~n12182 | ~n12180;
  assign n16713 = ~n16717;
  assign n10826 = ~n11733 & ~n11732;
  assign n15360 = ~n16837 & ~n15740;
  assign n11190 = n11167 & P2_REG3_REG_23__SCAN_IN;
  assign n13818 = ~n9548 | ~n9547;
  assign n16739 = ~n9891 | ~n9890;
  assign n15088 = ~n9877 | ~n9876;
  assign n10764 = ~n10763 & ~n12158;
  assign n10644 = ~n14769;
  assign n15789 = ~n14935;
  assign n15258 = ~n15371;
  assign n12181 = ~n12180;
  assign n16837 = ~n11623 & ~n11622;
  assign n11294 = ~n15371 & ~n14198;
  assign n10008 = ~n10007 & ~n10006;
  assign n10040 = ~n10039 & ~n10038;
  assign n9849 = ~n9848 & ~n9847;
  assign n15335 = ~n14769 | ~n16498;
  assign n10002 = n9972 & P1_REG3_REG_23__SCAN_IN;
  assign n9978 = ~n9977 & ~n9976;
  assign n11255 = ~n15371 & ~n14096;
  assign n9818 = ~n9817 & ~n9816;
  assign n9588 = ~n9583 & ~n9582;
  assign n13474 = ~n9458 | ~n9457;
  assign n9960 = ~n9959 & ~n9958;
  assign n15372 = ~n15371 & ~n15370;
  assign n11248 = ~n15371 & ~n13944;
  assign n9876 = ~n9875 & ~n9874;
  assign n11097 = ~n15371 & ~n13335;
  assign n13228 = ~n9427 | ~n9426;
  assign n9339 = ~n9332 | ~n15212;
  assign n15451 = ~n16502;
  assign n9929 = ~n9928 & ~n9927;
  assign n11733 = ~n10825 & ~n10824;
  assign n11150 = ~n15371 & ~n11149;
  assign n11144 = ~n15371 & ~n11143;
  assign n17062 = ~n11677 & ~n11676;
  assign n11318 = ~n11296;
  assign n9890 = ~n9889 & ~n9888;
  assign n11163 = ~n15371 & ~n11162;
  assign n11167 = n11154 & P2_REG3_REG_22__SCAN_IN;
  assign n11154 = n11119 & P2_REG3_REG_21__SCAN_IN;
  assign n15832 = ~n15547;
  assign n9972 = n9954 & P1_REG3_REG_22__SCAN_IN;
  assign n9202 = ~n9198 & ~n9197;
  assign n10824 = ~n11544 & ~n11543;
  assign n14825 = ~n11423 | ~n11492;
  assign n11373 = ~n11372;
  assign P1_U3083 = ~n10225 | ~P1_STATE_REG_SCAN_IN;
  assign n10765 = ~n12154;
  assign n15404 = ~n15163;
  assign n10120 = ~n11364 | ~n10118;
  assign n16474 = ~n16473 | ~n16472;
  assign n15713 = ~n15549;
  assign n11119 = n11101 & P2_REG3_REG_20__SCAN_IN;
  assign n9954 = n9923 & P1_REG3_REG_21__SCAN_IN;
  assign n12855 = ~n15285;
  assign n10887 = ~n10885;
  assign n9290 = ~n9331 | ~n9330;
  assign n10642 = ~n10885 & ~n10641;
  assign n9616 = ~n9611 & ~n9610;
  assign n9749 = ~n9745 & ~n9744;
  assign n9660 = ~n9655 & ~n9654;
  assign n11544 = ~n10823 & ~n10822;
  assign n9712 = ~n9708 & ~n9707;
  assign n10721 = ~n13806;
  assign n11101 = n10675 & P2_REG3_REG_19__SCAN_IN;
  assign P1_U4006 = ~n12117;
  assign n10774 = ~n15738;
  assign n11364 = ~n10117;
  assign n9449 = ~n9448 & ~n9447;
  assign n15766 = ~n10761 | ~n12156;
  assign n9217 = n9216 & n9215;
  assign n9342 = n9037 & P1_REG2_REG_5__SCAN_IN;
  assign n9538 = ~n9537 & ~n9536;
  assign n9699 = ~n9698 & ~n9697;
  assign n9842 = ~n9841 & ~n9840;
  assign n12934 = ~n12282;
  assign n9737 = ~n9736 & ~n9735;
  assign n9776 = n9775 & n9774;
  assign n9649 = ~n9648 & ~n9647;
  assign n11967 = ~n12088;
  assign n9578 = ~n9577 & ~n9576;
  assign n10550 = ~n10549 | ~P2_IR_REG_31__SCAN_IN;
  assign n9485 = ~n9484 & ~n9483;
  assign n10822 = ~n11436 & ~n11435;
  assign n9923 = n9884 & P1_REG3_REG_20__SCAN_IN;
  assign n10225 = ~n11417 | ~n10224;
  assign n9285 = ~n9282 | ~n9281;
  assign n12088 = ~n10451 & ~n10470;
  assign n10761 = ~n11369;
  assign n10050 = ~n15214 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n9037 = ~n9957;
  assign n9899 = ~n15214 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n15594 = ~n17091;
  assign n11417 = ~n10223 | ~n17086;
  assign n10217 = ~n10715 & ~n10716;
  assign n10549 = ~n10548 | ~n10547;
  assign n9884 = ~n9870 & ~n14827;
  assign n10675 = n10620 & P2_REG3_REG_18__SCAN_IN;
  assign n9952 = ~n15214 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n11436 = ~n10821 | ~n10820;
  assign n17091 = n10141 & n11423;
  assign n14876 = ~n10613 & ~n10612;
  assign n9870 = ~n9844 | ~P1_REG3_REG_18__SCAN_IN;
  assign n15595 = ~n15636;
  assign n10760 = ~n10141 | ~n17089;
  assign n9038 = ~n9041;
  assign n11369 = ~n11416 | ~n10174;
  assign n10715 = ~n13947;
  assign n10620 = ~n10593 & ~n10249;
  assign n9521 = ~n9520 & ~n9519;
  assign n10470 = ~n10450 & ~P2_IR_REG_10__SCAN_IN;
  assign n11365 = ~n14038 | ~n13938;
  assign n13968 = ~n10135 & ~n17073;
  assign n14099 = ~n10716;
  assign n15793 = ~n15422;
  assign n15791 = ~n15185;
  assign n11671 = ~n12043;
  assign n10175 = ~n11416;
  assign n9844 = ~n9812 & ~n14336;
  assign n10114 = ~n10111 | ~P1_B_REG_SCAN_IN;
  assign n10638 = ~n10637 | ~n10636;
  assign n10450 = ~n10449;
  assign n10220 = ~n10218 | ~P2_IR_REG_23__SCAN_IN;
  assign n11944 = ~n10427 | ~n10447;
  assign n9520 = ~n9518 | ~n9517;
  assign n14038 = ~n10119;
  assign n16967 = ~n17073 & ~n13329;
  assign n11378 = ~n10819 & ~n10818;
  assign n16847 = ~n13503 | ~n14836;
  assign n10593 = ~n10557 | ~P2_REG3_REG_15__SCAN_IN;
  assign n9266 = ~n9263 | ~n9262;
  assign n13461 = ~n9696 | ~n9695;
  assign n9128 = ~n10796;
  assign n10533 = ~n10532 | ~n10531;
  assign n17092 = ~n17086;
  assign n10557 = ~n10538 & ~n10957;
  assign n10042 = ~n10044 | ~n10022;
  assign n10113 = ~n13753 | ~n10112;
  assign n9597 = ~n9596;
  assign n9671 = ~n9674 | ~n9642;
  assign n9594 = ~n9570 & ~n9596;
  assign n11046 = ~n11045;
  assign n12135 = ~n10406 & ~n10405;
  assign n10449 = ~n10447 | ~P2_IR_REG_31__SCAN_IN;
  assign n9438 = ~n9440 | ~n9407;
  assign n9805 = ~n9773 | ~P1_IR_REG_31__SCAN_IN;
  assign n9812 = ~n9741 | ~P1_REG3_REG_16__SCAN_IN;
  assign n9726 = ~n9725;
  assign n10227 = ~n10229;
  assign n9632 = ~n9631;
  assign n10538 = ~n10248 | ~P2_REG3_REG_13__SCAN_IN;
  assign n10634 = ~n10633 | ~P2_IR_REG_31__SCAN_IN;
  assign n9232 = ~n9229 | ~n9228;
  assign n10491 = ~n10486 | ~n10485;
  assign n9407 = ~n9406 | ~SI_8_;
  assign n9596 = ~n9569 & ~SI_12_;
  assign n9562 = ~n9531 & ~SI_11_;
  assign n11532 = ~n9305 | ~n9374;
  assign n9517 = ~n9516 | ~n9515;
  assign n11363 = ~n10817 & ~n10816;
  assign n11846 = ~n11423;
  assign n10045 = ~n10044;
  assign n9569 = ~n9568;
  assign n9861 = n9863 ^ SI_19_;
  assign n9980 = n9982 ^ SI_23_;
  assign n11935 = ~n10352 & ~n10351;
  assign n9570 = ~n9568 & ~n9567;
  assign n9400 = ~n9399 | ~SI_7_;
  assign n9440 = ~n9405 | ~n9404;
  assign n9524 = ~n9523 | ~SI_10_;
  assign n9532 = ~n9530 & ~n9529;
  assign n9892 = n9894 ^ SI_20_;
  assign n9368 = ~n9367 | ~SI_6_;
  assign n9864 = ~n9863 | ~SI_19_;
  assign n11033 = n11035 ^ SI_27_;
  assign n9482 = ~n9480 | ~P1_IR_REG_31__SCAN_IN;
  assign n10061 = n10063 ^ SI_26_;
  assign n9762 = n9764 ^ SI_16_;
  assign n9680 = ~n9679;
  assign n9704 = ~n9652 | ~n9651;
  assign n9772 = ~n9694 & ~P1_IR_REG_15__SCAN_IN;
  assign n10131 = ~n10129 | ~n10128;
  assign n11042 = ~n11041;
  assign n11043 = ~n11041 & ~n11040;
  assign n9830 = n9832 ^ SI_18_;
  assign n9635 = n9634 & SI_13_;
  assign n9796 = n9798 ^ SI_17_;
  assign n9863 = ~n9836 | ~n9835;
  assign n9284 = ~n9283 | ~SI_4_;
  assign n9945 = ~n9919 | ~n9918;
  assign n9634 = ~n9600 | ~n9599;
  assign n9289 = ~n9288 | ~SI_5_;
  assign n9640 = ~n9638 & ~n9637;
  assign n9530 = ~n9528 & ~n9527;
  assign n9399 = ~n9371 | ~n9370;
  assign n9367 = ~n9292 | ~n9291;
  assign n9568 = ~n9566 & ~n9565;
  assign n9894 = ~n9867 | ~n9866;
  assign n9231 = ~n9230 | ~SI_2_;
  assign n9405 = ~n9403 & ~n9402;
  assign n9764 = ~n9729 | ~n9728;
  assign n11067 = ~n11053 | ~n11052;
  assign n9798 = ~n9768 | ~n9767;
  assign n9265 = ~n9264 | ~SI_3_;
  assign n9652 = ~n9584 & ~n11981;
  assign n14388 = ~n14585;
  assign n10129 = ~n10126 | ~P1_IR_REG_23__SCAN_IN;
  assign n9186 = ~n9153 | ~SI_0_;
  assign n9832 = ~n9802 | ~n9801;
  assign n9694 = ~n9689 | ~n9688;
  assign n9080 = ~n9077 | ~P1_IR_REG_24__SCAN_IN;
  assign n10066 = ~n11089 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n9566 = ~n11089 & ~n9571;
  assign n9283 = ~n9268 | ~n9267;
  assign n14582 = ~n14384;
  assign n11038 = ~n11089 & ~n14409;
  assign n10564 = n10196;
  assign n9835 = ~n11089 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n10718 = ~n10713 & ~n10712;
  assign n11059 = n11089 & P2_U3152;
  assign n9801 = ~n11089 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n10126 = ~n10125 | ~P1_IR_REG_31__SCAN_IN;
  assign n10018 = n11089 & P1_DATAO_REG_25__SCAN_IN;
  assign n10499 = ~n10480 & ~n10479;
  assign n9077 = ~n10130 | ~P1_IR_REG_31__SCAN_IN;
  assign n9479 = ~n9446 | ~P1_IR_REG_31__SCAN_IN;
  assign n9866 = ~n11089 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n9600 = ~n11089 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n10404 = ~n10399 & ~n10398;
  assign n9602 = ~n9684 & ~P1_IR_REG_12__SCAN_IN;
  assign n9288 = ~n9287 | ~n9286;
  assign n9230 = ~n9188 | ~n9187;
  assign n14577 = ~n14962;
  assign n9638 = n11089 & P1_DATAO_REG_14__SCAN_IN;
  assign n9494 = ~n9491 & ~n11724;
  assign n9684 = ~n9573 | ~n9572;
  assign n9099 = ~n9098 & ~n9097;
  assign n9188 = ~n10016 | ~P1_DATAO_REG_2__SCAN_IN;
  assign n9491 = ~n9421 | ~P1_REG3_REG_8__SCAN_IN;
  assign n10436 = ~n10432 & ~n10247;
  assign n10432 = ~n10385 | ~P2_REG3_REG_7__SCAN_IN;
  assign n9097 = ~n9096 | ~n9095;
  assign n9421 = ~n9418 & ~n11524;
  assign n9034 = ~n10016;
  assign n10189 = ~n10188 & ~P2_IR_REG_18__SCAN_IN;
  assign n9096 = ~n9094 & ~P1_IR_REG_20__SCAN_IN;
  assign n10385 = ~n10365 & ~n10364;
  assign n9113 = ~n9110 & ~P2_ADDR_REG_19__SCAN_IN;
  assign n9418 = ~n9318 | ~P1_REG3_REG_6__SCAN_IN;
  assign n10398 = ~n10397 | ~n10396;
  assign n10179 = ~n10178 | ~n10349;
  assign n10188 = ~n10187 | ~n10186;
  assign n9318 = ~n9315 & ~n9314;
  assign n10203 = ~n10202 | ~n10201;
  assign n10193 = ~n10192 | ~n10191;
  assign n10128 = ~n10127 | ~P1_IR_REG_31__SCAN_IN;
  assign n9079 = ~n9078 | ~P1_IR_REG_31__SCAN_IN;
  assign n9089 = ~n9093 | ~n9481;
  assign n9124 = ~n9123 | ~P1_IR_REG_31__SCAN_IN;
  assign n10365 = ~n10246 | ~P2_REG3_REG_4__SCAN_IN;
  assign n9056 = ~n9095 | ~n9055;
  assign n10207 = ~n10210 | ~P2_IR_REG_31__SCAN_IN;
  assign n10226 = ~P2_IR_REG_27__SCAN_IN;
  assign n9683 = ~P2_DATAO_REG_15__SCAN_IN;
  assign n9111 = ~P2_ADDR_REG_19__SCAN_IN | ~P1_ADDR_REG_19__SCAN_IN;
  assign n9109 = ~P1_RD_REG_SCAN_IN;
  assign n9703 = ~P1_REG3_REG_15__SCAN_IN | ~P1_REG3_REG_14__SCAN_IN;
  assign n9123 = ~P1_IR_REG_19__SCAN_IN;
  assign n9733 = ~P1_IR_REG_31__SCAN_IN;
  assign n10606 = ~P2_IR_REG_18__SCAN_IN;
  assign n10608 = ~P2_IR_REG_31__SCAN_IN;
  assign n9063 = ~P1_IR_REG_28__SCAN_IN;
  assign n9643 = ~P2_DATAO_REG_14__SCAN_IN;
  assign n9060 = ~P1_IR_REG_24__SCAN_IN & ~P1_IR_REG_23__SCAN_IN;
  assign n10182 = ~P2_IR_REG_9__SCAN_IN & ~P2_IR_REG_7__SCAN_IN;
  assign n10181 = ~P2_IR_REG_8__SCAN_IN & ~P2_IR_REG_6__SCAN_IN;
  assign n9061 = ~P1_IR_REG_26__SCAN_IN & ~P1_IR_REG_25__SCAN_IN;
  assign n9639 = ~SI_14_;
  assign n10210 = ~P2_IR_REG_26__SCAN_IN;
  assign n10247 = ~P2_REG3_REG_8__SCAN_IN | ~P2_REG3_REG_9__SCAN_IN;
  assign n10201 = ~P2_IR_REG_19__SCAN_IN & ~P2_IR_REG_18__SCAN_IN;
  assign n10202 = ~P2_IR_REG_22__SCAN_IN & ~P2_IR_REG_20__SCAN_IN;
  assign n10192 = ~P2_IR_REG_24__SCAN_IN & ~P2_IR_REG_23__SCAN_IN;
  assign n10127 = ~P1_IR_REG_23__SCAN_IN;
  assign n10197 = ~P2_IR_REG_23__SCAN_IN & ~P2_IR_REG_21__SCAN_IN;
  assign n10810 = ~P1_ADDR_REG_19__SCAN_IN;
  assign n9119 = ~P1_IR_REG_22__SCAN_IN;
  assign n10015 = ~P2_DATAO_REG_25__SCAN_IN;
  assign n10249 = ~P2_REG3_REG_16__SCAN_IN | ~P2_REG3_REG_17__SCAN_IN;
  assign n9651 = P1_REG3_REG_13__SCAN_IN & P1_REG3_REG_12__SCAN_IN;
  assign n10403 = ~P2_IR_REG_8__SCAN_IN;
  assign n9101 = ~P1_IR_REG_21__SCAN_IN;
  assign n10019 = ~SI_25_;
  assign n10629 = ~P2_IR_REG_19__SCAN_IN | ~P2_IR_REG_31__SCAN_IN;
  assign n10485 = ~P2_IR_REG_11__SCAN_IN & ~P2_IR_REG_10__SCAN_IN;
  assign n9300 = ~P1_IR_REG_5__SCAN_IN;
  assign n10198 = ~P2_IR_REG_25__SCAN_IN & ~P2_IR_REG_24__SCAN_IN;
  assign n10635 = ~P2_IR_REG_21__SCAN_IN;
  assign n15858 = ~n15844 | ~n15843;
  assign n15857 = ~n15856 & ~n15855;
  assign n15785 = ~n15786 | ~n16510;
  assign n15788 = ~n15786 | ~n16514;
  assign n15667 = ~n15668 | ~n16510;
  assign n15670 = ~n15668 | ~n16514;
  assign n16479 = ~n16477 | ~n16476;
  assign n15503 = ~n15501 | ~n16514;
  assign n15731 = ~n15775 & ~n15845;
  assign n15719 = ~n15775 & ~n14769;
  assign n15822 = ~n15811 | ~n10132;
  assign n15500 = ~n15501 | ~n16510;
  assign n16851 = ~n16850 | ~n16849;
  assign n15665 = ~n15663 & ~n15662;
  assign n15826 = ~n15823 & ~n16022;
  assign n15773 = ~n15772 & ~n15771;
  assign n15497 = ~n15496 & ~n15495;
  assign n15680 = ~n15681 | ~n15800;
  assign n10033 = ~n15687 & ~n15685;
  assign n15487 = ~n15485 | ~n15484;
  assign n17075 = ~n17078 & ~n17072;
  assign n15472 = ~n15491 & ~n15845;
  assign n15683 = ~n15681 | ~n15804;
  assign n15491 = ~n15478;
  assign n17033 = ~n17032 ^ n17072;
  assign n15790 = ~n15757 | ~n15756;
  assign n17078 = ~n17071 | ~n17070;
  assign n15562 = ~n15560 & ~n15559;
  assign n11250 = ~n15526;
  assign n15629 = ~n15630 | ~n15800;
  assign n15632 = ~n15630 | ~n15804;
  assign n15607 = ~n15627 | ~n15745;
  assign n16963 = ~n17036 & ~n16962;
  assign n16844 = ~n17070 | ~n16843;
  assign n15460 = ~n15458 | ~n16514;
  assign n15457 = ~n15458 | ~n16510;
  assign n16434 = ~n16433 | ~n16451;
  assign n16032 = ~n16030 | ~n16029;
  assign n15676 = ~n15671 & ~n15789;
  assign n15113 = ~n15131 | ~n15720;
  assign n15362 = ~n15361 & ~n15360;
  assign n15224 = ~n15359 | ~n15762;
  assign n15626 = ~n15625 & ~n15624;
  assign n15130 = ~n15129 & ~n15128;
  assign n15718 = ~n15717 | ~n15716;
  assign n16825 = ~n16807 | ~n16806;
  assign n15363 = ~n15359 | ~n15791;
  assign n15361 = ~n16839 & ~n15422;
  assign n15381 = ~n15450 | ~n15847;
  assign n15455 = ~n15450 | ~n16500;
  assign n15717 = ~n15712 | ~n15832;
  assign n15060 = ~n15057 | ~n15056;
  assign n15454 = ~n15453 & ~n15452;
  assign n15616 = ~n15620 & ~n15608;
  assign n16959 = ~n16958 | ~n16957;
  assign n15625 = ~n15620 & ~n15619;
  assign n15604 = ~n15620 & ~n15404;
  assign n15121 = ~n15124 & ~n15845;
  assign n15748 = ~n15646 | ~n15645;
  assign n15039 = ~n15057 | ~n15720;
  assign n16807 = ~n16791 | ~n16808;
  assign n15505 = ~n9968 & ~n9967;
  assign n15269 = ~n11172 | ~n16016;
  assign n17028 = ~n17027 | ~n17026;
  assign n16955 = ~n16956 | ~n17063;
  assign n15352 = ~n15351 & ~n15360;
  assign n16426 = ~n16445;
  assign n15384 = ~n15383 & ~n15452;
  assign n15427 = ~n15426 & ~n15425;
  assign n15267 = ~n15382 | ~n15847;
  assign n15353 = ~n15350 | ~n15791;
  assign n17066 = ~n17065 | ~n17064;
  assign n15047 = ~n15050 & ~n15845;
  assign n16786 = ~n16821 | ~n16776;
  assign n15211 = ~n15350 | ~n15762;
  assign n16422 = ~n16432 & ~n16452;
  assign n15426 = ~n15421 & ~n15619;
  assign n15385 = ~n15382 | ~n16500;
  assign n15383 = ~n16432 & ~n15451;
  assign n15311 = ~n15329 | ~n15745;
  assign n17027 = ~n17025 & ~n17024;
  assign n15605 = ~n15599 | ~n15598;
  assign n11131 = ~n15003 & ~n15488;
  assign n15169 = ~n15192 | ~n15745;
  assign n15484 = ~n15483 & ~n15482;
  assign n15770 = ~n15792 | ~n15762;
  assign n16025 = ~n16024 & ~n16023;
  assign n15328 = ~n15327 & ~n15326;
  assign n16804 = ~n16803 | ~n16802;
  assign n16432 = ~n16449;
  assign n16827 = ~n17063 | ~n16688;
  assign n17035 = ~n17063 & ~n17062;
  assign n17125 = ~n17148;
  assign n15343 = ~n15342 & ~n15341;
  assign n15406 = ~n15400 | ~n15399;
  assign n15191 = ~n15190 & ~n15189;
  assign n15599 = ~n15593 | ~n10774;
  assign n16023 = ~n16022 | ~n16021;
  assign n15327 = ~n15322 & ~n15619;
  assign n17148 = n17116 ^ n17115;
  assign n15003 = ~n11129 | ~n11128;
  assign n9938 = ~n9912 | ~n9911;
  assign n15190 = ~n15184 & ~n15619;
  assign n15342 = ~n15282 | ~n15281;
  assign n11138 = ~n14994 | ~n14078;
  assign n15166 = ~n15165 | ~n15164;
  assign n15854 = ~n16501 | ~n15847;
  assign n17059 = ~n16951 & ~n16950;
  assign n15652 = ~n15672 | ~n15762;
  assign n15768 = ~n15764 & ~n15763;
  assign n15761 = ~n15764 & ~n15759;
  assign n11341 = ~n11324 | ~n11344;
  assign n17116 = ~n17108 ^ n17107;
  assign n15852 = ~n16411 & ~n15848;
  assign n9910 = ~n9883 | ~n14944;
  assign n17022 = ~n17021 & ~n17020;
  assign n11321 = ~n11323 | ~n15527;
  assign n15650 = ~n17127 & ~n15763;
  assign n15247 = ~n15246 & ~n15245;
  assign n16862 = ~n16860 | ~n16947;
  assign n16413 = ~n16406;
  assign n15825 = ~n15824 & ~n15834;
  assign n16024 = n16503 ^ n16427;
  assign n11202 = ~n15246 & ~n15488;
  assign n15727 = ~n15824 & ~n15848;
  assign n15794 = ~n16520 | ~n15793;
  assign n15729 = ~n15776 | ~n15847;
  assign n16950 = ~n17110 & ~n15752;
  assign n17102 = n17119 ^ n17117;
  assign n15673 = ~n17110 | ~n15793;
  assign n14779 = ~n14815 | ~n15720;
  assign n15778 = ~n15777 | ~n16502;
  assign n15246 = ~n11200 | ~n11199;
  assign n15309 = ~n15304 | ~n15303;
  assign n15846 = ~n15777 & ~n15723;
  assign n17106 = ~n17110 | ~n17111;
  assign n14818 = ~n14815 | ~n14814;
  assign n16860 = ~n16859 | ~n16858;
  assign n9883 = ~n15077;
  assign n17021 = n17110 ^ n17112;
  assign n17114 = ~n17110 | ~n17109;
  assign n17119 = n10080 ^ n17107;
  assign n14589 = ~n15257 | ~n14582;
  assign n14712 = ~n14709 | ~n14708;
  assign n14581 = ~n15257 | ~n11059;
  assign n14990 = ~n15068 & ~n15758;
  assign n14815 = ~n14777 & ~n14776;
  assign n14905 = ~n14894 | ~n15527;
  assign n15412 = ~n15411 | ~n15745;
  assign n17118 = ~n17117;
  assign n16527 = ~n16526 | ~n16525;
  assign n14408 = ~n15202 | ~n11059;
  assign n15411 = ~n15424 | ~n17072;
  assign n16946 = ~n16945 | ~n17051;
  assign n15647 = ~n16854 | ~n15609;
  assign n14787 = ~n14808 & ~n15845;
  assign n11308 = ~n15202 | ~n10310;
  assign n11324 = ~n11300 & ~n11299;
  assign n14941 = ~n14938 | ~n14937;
  assign n14413 = ~n15202 | ~n14582;
  assign n16021 = ~n16020 & ~n16019;
  assign n10080 = ~n10079 | ~n10078;
  assign n10737 = ~n14707 | ~n15720;
  assign n10082 = ~n16524 | ~n17111;
  assign n15622 = ~n16524 | ~n15793;
  assign n17054 = ~n16524 ^ n16853;
  assign n17056 = ~n16864 | ~n16863;
  assign n15568 = ~n15659 | ~n15847;
  assign n15660 = ~n16436 | ~n16502;
  assign n10169 = ~n16524 | ~n15578;
  assign n16945 = ~n17050 | ~n16944;
  assign n16439 = ~n16050 | ~n16049;
  assign n14729 = ~n14719 | ~n15527;
  assign n14928 = ~n14936 | ~n14927;
  assign n14707 = ~n10685 | ~n10684;
  assign n10079 = ~n16524 | ~n17109;
  assign n14976 = ~n15067 | ~n15745;
  assign n10735 = ~n14701 & ~n15845;
  assign n15417 = ~n16814 & ~n15763;
  assign n14763 = ~n14760 | ~n14759;
  assign n15575 = ~n9999 | ~n9998;
  assign n15707 = ~n16405 & ~n16048;
  assign n15816 = ~n16814 & ~n17126;
  assign n14979 = ~n14977 | ~n17014;
  assign n10057 = ~n10056 | ~n10055;
  assign n15723 = ~n15565 | ~n16048;
  assign n10054 = ~n10053 | ~n10052;
  assign n15067 = ~n14973 & ~n14972;
  assign n16856 = ~n16787 & ~n16814;
  assign n15684 = ~n10032 & ~n10031;
  assign n15423 = ~n16814 & ~n15422;
  assign n15945 = ~n15704 | ~n16048;
  assign n15828 = ~n15704 & ~n16048;
  assign n16019 = ~n16018 | ~n16017;
  assign n15600 = ~n16816 | ~n16814;
  assign n16810 = ~n16780 | ~n16779;
  assign n14202 = ~n14197 | ~n11059;
  assign n10052 = ~n16788 | ~n17109;
  assign n15409 = ~n16788 | ~n15408;
  assign n14467 = ~n14464 | ~n14463;
  assign n15602 = ~n16787 | ~n16788;
  assign n10055 = ~n16788 | ~n17111;
  assign n15609 = ~n16788 & ~n15408;
  assign n14751 = ~n14758 | ~n14927;
  assign n15493 = ~n15558 | ~n16502;
  assign n14650 = ~n14639 | ~n15527;
  assign n11290 = ~n11267 | ~n11266;
  assign n16398 = ~n16387 | ~n16386;
  assign n15296 = ~n17018;
  assign n16863 = ~n16781 | ~n16778;
  assign n16788 = ~n10051 | ~n10050;
  assign n15940 = ~n16392 & ~n15557;
  assign n14698 = ~n14695 | ~n14694;
  assign n14934 = ~n14913 | ~n14912;
  assign n15177 = ~n15186 & ~n15174;
  assign n16376 = ~n16375 | ~n16374;
  assign n11285 = ~n16392 & ~n14448;
  assign n9999 = ~n9995 | ~n9994;
  assign n14387 = ~n14385 & ~n14384;
  assign n16383 = ~n16385 | ~n16382;
  assign n10028 = ~n10027 | ~n10026;
  assign n10996 = ~n14457 | ~n14047;
  assign n10031 = ~n10030 | ~n10029;
  assign n14738 = ~n14757 & ~n15218;
  assign n15314 = ~n16782 | ~n15313;
  assign n14214 = ~n14212 | ~n16510;
  assign n16764 = ~n16763 & ~n16762;
  assign n16868 = ~n16929;
  assign n14686 = ~n14693 | ~n14927;
  assign n16874 = ~n16771 | ~n16768;
  assign n10029 = ~n16782 | ~n17111;
  assign n10026 = ~n16782 | ~n17109;
  assign n15402 = ~n16781 | ~n16782;
  assign n15539 = ~n15531 | ~n15867;
  assign n14520 = ~n14519 | ~n15527;
  assign n14211 = ~n14212 | ~n16514;
  assign n14042 = ~n14037 | ~n14582;
  assign n15287 = ~n15531 | ~n15285;
  assign n16385 = ~n16381 | ~n16380;
  assign n16370 = ~n16373 | ~n16372;
  assign n14098 = ~n14095 & ~n14094;
  assign n11181 = ~n11180 | ~n11179;
  assign n9991 = ~n9990 | ~n9989;
  assign n14757 = ~n14736 | ~n14735;
  assign n9996 = ~n9993 | ~n9992;
  assign n16782 = ~n10025 | ~n10024;
  assign n14128 = ~n14126 | ~n16514;
  assign n15935 = ~n15933 & ~n15932;
  assign n15337 = ~n15283 & ~n16378;
  assign n14125 = ~n14126 | ~n16510;
  assign n15173 = ~n15312;
  assign n16929 = ~n16870 | ~n16866;
  assign n15100 = ~n16014;
  assign n14613 = ~n14610 | ~n14609;
  assign n15468 = ~n15283 | ~n16378;
  assign n14115 = ~n14113 | ~n16510;
  assign n16870 = ~n16865;
  assign n15172 = ~n15579 | ~n15171;
  assign n9992 = ~n15579 | ~n17111;
  assign n15306 = ~n15697 | ~n15579;
  assign n9989 = ~n15579 | ~n17109;
  assign n15445 = ~n16362 | ~n15867;
  assign n14112 = ~n14113 | ~n16514;
  assign n15581 = ~n15579 | ~n15578;
  assign n15276 = ~n15932;
  assign n14657 = ~n14656 | ~n14655;
  assign n11176 = ~n16362 | ~n11177;
  assign n14676 = ~n14692 & ~n15218;
  assign n16355 = ~n16359 | ~n16349;
  assign n14445 = ~n14444 | ~n15527;
  assign n14093 = ~n14077 | ~n14076;
  assign n15506 = ~n9970 | ~n9969;
  assign n13946 = ~n13943 & ~n14094;
  assign n14986 = ~n15511 & ~n15763;
  assign n10986 = ~n10981 | ~n15527;
  assign n15516 = ~n15511 & ~n17126;
  assign n9964 = ~n9963 | ~n9962;
  assign n15171 = ~n15511 | ~n14982;
  assign n14983 = ~n15511 & ~n14982;
  assign n15579 = ~n9988 | ~n9987;
  assign n14077 = ~n14110 | ~n15720;
  assign n14489 = ~n14486 | ~n14485;
  assign n13940 = ~n13943 & ~n14384;
  assign n11030 = ~n11025 | ~n15527;
  assign n16341 = ~n16351 | ~n16350;
  assign n16366 = ~n11164 & ~n11163;
  assign n14023 = ~n14021 | ~n16514;
  assign n14290 = ~n14291 | ~n15804;
  assign n14020 = ~n14021 | ~n16510;
  assign n14293 = ~n14291 | ~n15800;
  assign n14503 = ~n14502 | ~n14927;
  assign n9970 = ~n15160 | ~n17111;
  assign n11004 = ~n14462 & ~n15488;
  assign n15929 = ~n15927 & ~n15926;
  assign n15119 = ~n15125 | ~n15847;
  assign n9939 = ~n9933 ^ n17107;
  assign n9963 = ~n15160 | ~n17109;
  assign n14494 = ~n14492 & ~n15218;
  assign n13920 = ~n13921 | ~n16514;
  assign n9933 = ~n9932 | ~n9931;
  assign n14370 = ~n14361 | ~n14360;
  assign n13923 = ~n13921 | ~n16510;
  assign n14380 = ~n14381 | ~n15800;
  assign n15928 = ~n15115 | ~n16347;
  assign n14744 = ~n14743 | ~n14742;
  assign n14291 = ~n14288 | ~n14287;
  assign n11177 = ~n15114 | ~n15115;
  assign n13808 = ~n13805 & ~n14094;
  assign n13752 = ~n13805;
  assign n16353 = ~n16350;
  assign n14383 = ~n14381 | ~n15804;
  assign n10858 = ~n14207 & ~n15488;
  assign n15052 = ~n16333 | ~n16502;
  assign n14310 = ~n14308 & ~n15218;
  assign n14399 = ~n15800 | ~n14401;
  assign n14067 = ~n14102 | ~n10644;
  assign n15081 = ~n9903 ^ n17107;
  assign n16866 = ~n14981 | ~n14906;
  assign n16736 = ~n16735 | ~n16879;
  assign n14402 = ~n15804 | ~n14401;
  assign n16745 = ~n16741 | ~n16740;
  assign n15044 = ~n15051 | ~n15847;
  assign n9932 = ~n14981 | ~n17109;
  assign n14978 = ~n14981 | ~n15512;
  assign n15018 = ~n15867 | ~n16333;
  assign n15114 = ~n16333 & ~n15043;
  assign n14061 = ~n14060 | ~n14059;
  assign n16350 = ~n16340 | ~n16339;
  assign n14717 = ~n14716 | ~n14715;
  assign n15924 = ~n16337 & ~n16334;
  assign n13897 = ~n16514 | ~n13899;
  assign n14060 = ~n14122 | ~n15720;
  assign n14306 = ~n15804 | ~n14305;
  assign n11148 = ~n16337 | ~n16338;
  assign n10953 = ~n15527 | ~n10952;
  assign n13900 = ~n16510 | ~n13899;
  assign n14162 = ~n14161 | ~n15745;
  assign n16735 = ~n16734 | ~n16733;
  assign n15092 = ~n15087 & ~n17126;
  assign n14303 = ~n15800 | ~n14305;
  assign n13705 = ~n13708 & ~n14384;
  assign n15080 = ~n9905 | ~n9904;
  assign n13710 = ~n13708 & ~n14094;
  assign n16333 = ~n16337;
  assign n14368 = ~n14371 & ~n15608;
  assign n14035 = ~n15800 | ~n14034;
  assign n11135 = ~n13071 & ~n14996;
  assign n14176 = ~n15527 | ~n14175;
  assign n14376 = ~n14371 & ~n15619;
  assign n16008 = ~n14767 | ~n14766;
  assign n16744 = ~n16743 & ~n16742;
  assign n9901 = ~n16738 | ~n17109;
  assign n14257 = ~n14256 | ~n15527;
  assign n9904 = ~n16738 | ~n17111;
  assign n15922 = ~n16321 | ~n15031;
  assign n16867 = ~n14924 & ~n16738;
  assign n16547 = ~n16536 | ~n16875;
  assign n14716 = ~n11226 | ~n11225;
  assign n15043 = ~n11175 | ~n14997;
  assign n14032 = ~n15804 | ~n14034;
  assign n16734 = ~n16731 | ~n16730;
  assign n14073 = ~n14072 & ~n15547;
  assign n17010 = ~n16879 | ~n16875;
  assign n14810 = ~n16298 | ~n16502;
  assign n14846 = ~n9859 | ~n9858;
  assign n14811 = ~n14809 | ~n16500;
  assign n15919 = ~n15917 & ~n15916;
  assign n9907 = ~n9880 ^ n17107;
  assign n15920 = ~n14997 | ~n16322;
  assign n14998 = ~n14997 & ~n15451;
  assign n15917 = ~n15915 | ~n16308;
  assign n11223 = n16302 ^ n11296;
  assign n13916 = ~n13932 & ~n16498;
  assign n14766 = ~n16302 | ~n16299;
  assign n14300 = ~n14294 & ~n15619;
  assign n16535 = ~n16549 & ~n16534;
  assign n13906 = ~n13932 & ~n14769;
  assign n14690 = ~n14688 | ~n15791;
  assign n14952 = ~n14948 & ~n17126;
  assign n14142 = ~n14294 & ~n15608;
  assign n9879 = ~n14748 | ~n17109;
  assign n13732 = ~n13728 | ~n13727;
  assign n13986 = ~n14069 | ~n15832;
  assign n9882 = ~n14748 | ~n17111;
  assign n16875 = ~n14748 | ~n14850;
  assign n10734 = ~n10733 | ~n10732;
  assign n14749 = ~n14748 | ~n15088;
  assign n16549 = ~n16533 | ~n16532;
  assign n14601 = ~n14599 & ~n15185;
  assign n14230 = ~n14229 & ~n15738;
  assign n13728 = ~n13890 | ~n10644;
  assign n11111 = ~n16006;
  assign n16720 = ~n16723 | ~n16722;
  assign n14248 = ~n10945 | ~n13645;
  assign n14704 = ~n14702 | ~n16500;
  assign n11092 = ~n11091 | ~n11090;
  assign n13812 = ~n9042 | ~n13846;
  assign n14599 = ~n16530 & ~n14600;
  assign n16723 = ~n16715 | ~n16714;
  assign n16543 = ~n16539 | ~n16538;
  assign n16530 = ~n16548;
  assign n14684 = ~n16548 | ~n16534;
  assign n9855 = ~n16548 | ~n17111;
  assign n9852 = ~n16548 | ~n17109;
  assign n16721 = ~n16711 | ~n16710;
  assign n14396 = ~n14391 & ~n15619;
  assign n9791 = ~n9788 ^ n17107;
  assign n11134 = ~n10731 | ~n10992;
  assign n16711 = ~n16707 | ~n16706;
  assign n13957 = ~n15738 & ~n13955;
  assign n13746 = ~n13737;
  assign n13731 = ~n13730 & ~n15547;
  assign n15909 = ~n15906 | ~n15905;
  assign n9790 = ~n16716 | ~n17111;
  assign n14482 = ~n16716 | ~n16717;
  assign n10236 = ~n13065 | ~n10310;
  assign n15906 = ~n15904 | ~n15903;
  assign n10992 = ~n16056 & ~n10844;
  assign n9824 = ~n14797 | ~n17111;
  assign n9787 = ~n16716 | ~n17109;
  assign n9821 = ~n14797 | ~n17109;
  assign n14606 = ~n14797 | ~n14605;
  assign n16706 = ~n16705 | ~n16704;
  assign n15904 = ~n15901 | ~n15900;
  assign n15883 = ~n16053 | ~n16051;
  assign n11208 = n16053 ^ n11296;
  assign n10600 = ~n16053 | ~n16054;
  assign n13627 = ~n13626 & ~n15547;
  assign n9756 = n9753 ^ n9752;
  assign n13600 = ~n13657 & ~n15404;
  assign n13700 = ~n13698 | ~n13697;
  assign n13787 = ~n15738 & ~n13782;
  assign n13448 = ~n13445 | ~n13444;
  assign n15907 = ~n14051 | ~n16272;
  assign n14347 = ~n17002;
  assign n13690 = ~n10446 | ~n10445;
  assign n14875 = ~n14565 & ~n14564;
  assign n16001 = ~n16272 | ~n16279;
  assign n14284 = ~n16692 | ~n16693;
  assign n9751 = ~n16692 | ~n17109;
  assign n9755 = ~n16692 | ~n17111;
  assign n14051 = ~n15997 | ~n10666;
  assign n15997 = ~n10665 | ~n14068;
  assign n16280 = ~n14447;
  assign n11015 = ~n11019 | ~n14433;
  assign n14562 = ~n14427 | ~n14426;
  assign n10863 = n9715 ^ n9752;
  assign n13442 = ~n13259 | ~n13258;
  assign n11013 = n14447 ^ n11296;
  assign n17000 = ~n14129 & ~n14344;
  assign n16257 = ~n16256 & ~n16255;
  assign n14070 = ~n10665 | ~n10666;
  assign n15891 = ~n15889 | ~n15888;
  assign n14868 = ~n14560 & ~n14559;
  assign n16677 = ~n16659 | ~n16658;
  assign n11010 = ~n11014 | ~n11017;
  assign n14426 = ~n13870 | ~n13869;
  assign n16659 = ~n16656 | ~n16655;
  assign n9797 = ~n9766 | ~n9765;
  assign n15996 = ~n10666 | ~n10664;
  assign n9667 = ~n9663 ^ n17107;
  assign n11014 = n16266 ^ n11318;
  assign n9714 = ~n14296 | ~n17109;
  assign n14557 = ~n14417 | ~n14416;
  assign n13869 = ~n13867 & ~n13866;
  assign n13994 = ~n14068 | ~n10664;
  assign n9718 = ~n14296 | ~n17111;
  assign n16260 = ~n16246 | ~n16245;
  assign n14416 = ~n13879 | ~n13878;
  assign n10394 = ~n13250 | ~n10392;
  assign n10972 = n10974 ^ n10975;
  assign n14068 = ~n16243 | ~n16248;
  assign n10545 = ~n16243 | ~n16244;
  assign n10974 = n16247 ^ n11296;
  assign n9622 = n9619 ^ n9752;
  assign n16645 = ~n16642 | ~n16641;
  assign n13878 = ~n13877 & ~n13876;
  assign n10554 = ~n12295 | ~n10310;
  assign n14148 = ~n16919 | ~n14145;
  assign n16672 = ~n16657 | ~n14151;
  assign n9662 = ~n16657 | ~n17109;
  assign n16996 = ~n14130 | ~n13954;
  assign n10663 = ~n16252;
  assign n13864 = ~n13539 & ~n13538;
  assign n9727 = ~n9724 | ~n9723;
  assign n9618 = ~n16668 | ~n17109;
  assign n16994 = ~n16660 | ~n16661;
  assign n13770 = ~n13454 & ~n13453;
  assign n13873 = ~n13533 & ~n13532;
  assign n13911 = ~n16225 | ~n13720;
  assign n10517 = ~n12077 | ~n10310;
  assign n9508 = ~n9507;
  assign n13197 = ~n10833 & ~n12835;
  assign n13637 = ~n13738 | ~n13688;
  assign n16198 = ~n16194 & ~n16175;
  assign n16989 = ~n16637 | ~n16914;
  assign n12921 = ~n12585 & ~n12584;
  assign n13531 = ~n12916 & ~n12915;
  assign n15553 = ~n15552 | ~n15551;
  assign n9555 = n9551 ^ n17107;
  assign n13102 = ~n13100 | ~n13099;
  assign n16624 = ~n16935 | ~n16915;
  assign n9507 = n9503 ^ n17107;
  assign n9468 = ~n9465;
  assign n10498 = ~n11995 | ~n10310;
  assign n12869 = ~n10652 | ~n16143;
  assign n12836 = ~n10832 & ~n12572;
  assign n13599 = ~n13792 | ~n13598;
  assign n16935 = ~n13595 | ~n13783;
  assign n12914 = ~n12579 & ~n12578;
  assign n13738 = ~n16205;
  assign n16915 = ~n13611 | ~n13594;
  assign n9550 = ~n13837 | ~n17109;
  assign n15894 = ~n16188 & ~n16192;
  assign n9467 = ~n9466;
  assign n12573 = ~n10831 & ~n12320;
  assign n14448 = ~n15867;
  assign n12694 = ~n10651 | ~n10650;
  assign n16427 = ~n11331 | ~n11330;
  assign n13837 = ~n9539 | ~n9538;
  assign n16985 = ~n16616 | ~n16617;
  assign n9363 = ~n9362 | ~n9361;
  assign n16983 = ~n16606;
  assign n15736 = ~n17131;
  assign n16151 = ~n16132 | ~n16146;
  assign n14078 = ~n15845;
  assign n15977 = ~n10375 | ~n10376;
  assign n11330 = n11329 & n11328;
  assign n14079 = ~n15720 | ~n16038;
  assign n15861 = ~n15527;
  assign n17131 = ~n12050 | ~n12049;
  assign n11201 = ~n15720 & ~P2_REG2_REG_24__SCAN_IN;
  assign n15971 = ~n12889;
  assign n15482 = ~n16379 & ~n16488;
  assign n9362 = ~n9358 | ~n12780;
  assign n12321 = ~n10830 & ~n12139;
  assign n9354 = ~n12781 | ~n9353;
  assign n15976 = ~n12695;
  assign n16148 = ~n13443 | ~n13017;
  assign n11130 = ~n15720 & ~P2_REG2_REG_21__SCAN_IN;
  assign n16146 = ~n13020 | ~n12646;
  assign n10431 = ~n11778 | ~n10310;
  assign n12873 = ~n12899 | ~n16115;
  assign n9393 = ~n9391 | ~n9390;
  assign n9389 = ~n9388 | ~n9387;
  assign n9360 = ~n9359;
  assign n17128 = ~n10156 | ~n15765;
  assign n16514 = ~n16516;
  assign n13184 = ~n16160;
  assign n16510 = ~n16511;
  assign n15532 = ~n15872;
  assign n16132 = ~n13032 | ~n13251;
  assign n16110 = ~n13014 & ~n13078;
  assign n12994 = ~n13014;
  assign n16226 = ~n10509 & ~n10508;
  assign n14796 = ~n14853;
  assign n16244 = ~n10544 & ~n10543;
  assign n14506 = ~n10253 | ~n10252;
  assign n16277 = ~n10576 | ~n10575;
  assign n16192 = ~n10484 & ~n10483;
  assign n14167 = ~n10526 & ~n10525;
  assign n10077 = ~n10073 & ~n10072;
  assign n15849 = ~P2_REG3_REG_28__SCAN_IN | ~n11312;
  assign n16051 = ~n10599 | ~n10598;
  assign n13642 = ~n10466 & ~n10465;
  assign n13424 = ~n13364;
  assign n10894 = ~n10893 | ~n10892;
  assign n13288 = ~n10391 | ~n10390;
  assign n12140 = ~n10829 & ~n12001;
  assign n15765 = ~P1_REG3_REG_28__SCAN_IN | ~n10155;
  assign n12779 = ~n9329 | ~n9328;
  assign n10526 = ~n10522 | ~n10521;
  assign n10153 = ~n10155;
  assign n15313 = ~n15763;
  assign n9327 = ~n9326 | ~n9325;
  assign n10509 = ~n10505 | ~n10504;
  assign n12502 = ~n10783 | ~n10782;
  assign n12501 = ~n16971;
  assign n10444 = ~n10440 | ~n10439;
  assign n10410 = ~n11739 | ~n10310;
  assign n12876 = ~n13078;
  assign n10877 = ~n11464 | ~n12020;
  assign n12007 = ~n12006 | ~n12005;
  assign n9511 = ~n9439 & ~n9438;
  assign n16979 = ~n16890 | ~n16598;
  assign n10155 = ~n10152 & ~n10151;
  assign n15696 = ~n17136;
  assign n10679 = n10674 & n10673;
  assign n12819 = ~n9352 | ~n9351;
  assign n17041 = ~n16579;
  assign n16115 = ~n12687;
  assign n10152 = ~n10070 | ~P1_REG3_REG_26__SCAN_IN;
  assign n10726 = ~n12020 & ~n16486;
  assign n11464 = ~n12006;
  assign n11664 = ~n11646 | ~P2_STATE_REG_SCAN_IN;
  assign n15800 = ~n15801;
  assign n15804 = ~n15806;
  assign n11646 = ~n11635 | ~n11634;
  assign n10766 = ~n10765 | ~n10764;
  assign n10465 = ~n10464 | ~n10463;
  assign n12687 = ~n10336 | ~n10335;
  assign n10484 = ~n10478 | ~n10477;
  assign n9240 = ~n9239 | ~n9238;
  assign n11105 = n11100 & n11099;
  assign n11102 = ~n11804 | ~P2_REG2_REG_21__SCAN_IN;
  assign n10516 = n10515 & n10514;
  assign n11123 = n11118 & n11117;
  assign n10673 = ~n11804 | ~P2_REG2_REG_20__SCAN_IN;
  assign n10288 = n10284 & n10283;
  assign n11168 = ~n11804 | ~P2_REG2_REG_24__SCAN_IN;
  assign n11155 = ~n11804 | ~P2_REG2_REG_23__SCAN_IN;
  assign n11120 = ~n11804 | ~P2_REG2_REG_22__SCAN_IN;
  assign n10588 = ~n15258 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n10568 = ~n15258 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n13783 = ~n9500 | ~n9499;
  assign n13855 = ~n9588 | ~n9587;
  assign n14605 = ~n9819 | ~n9818;
  assign n10723 = ~n11611 & ~P2_D_REG_0__SCAN_IN;
  assign n11635 = ~n10221 | ~n13709;
  assign n11307 = ~n15258 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n13121 = ~n13104;
  assign n16568 = ~n12671;
  assign n10749 = ~n10765 | ~n10123;
  assign n10300 = ~n10297 | ~n10296;
  assign n10234 = ~n15371 & ~n10231;
  assign n16666 = ~n9616 | ~n9615;
  assign n16678 = ~n9660 | ~n9659;
  assign n14527 = ~n9712 | ~n9711;
  assign n16717 = ~n9785 | ~n9784;
  assign n9369 = ~n9366 | ~n9365;
  assign n10123 = ~n12158 & ~n12180;
  assign n11611 = ~n10717 | ~n14099;
  assign n13104 = ~n9386 | ~n9385;
  assign n10615 = ~n15371 & ~n10604;
  assign n16693 = ~n9749 | ~n9748;
  assign n10717 = ~n10715 | ~n10714;
  assign n10880 = ~n10724 | ~n11631;
  assign n10722 = ~n10721 & ~n14099;
  assign n12157 = ~n12156 & ~n12155;
  assign n10233 = ~n11632 & ~n16038;
  assign n10552 = ~n13874 | ~n10586;
  assign n9132 = ~n9131 & ~n9130;
  assign n10614 = ~n14566 & ~n11632;
  assign n12794 = ~n12668;
  assign n9036 = ~n10310;
  assign n10724 = ~n9039 | ~n16038;
  assign n10122 = ~n11364 | ~n10121;
  assign n15407 = ~n15766;
  assign n12668 = ~n9270 | ~n9269;
  assign n11372 = ~n11364 & ~n11369;
  assign n10714 = ~P2_B_REG_SCAN_IN ^ n13806;
  assign n9172 = ~n9169 & ~n9168;
  assign n11007 = ~n10595 & ~n10620;
  assign n15549 = n11631 & n14404;
  assign n12153 = ~n10761 | ~n10760;
  assign n16492 = ~n13709 & ~P2_U3152;
  assign n14833 = ~n11417 | ~n11410;
  assign n10719 = ~n13947 & ~n14099;
  assign n9147 = ~n9143 & ~n9142;
  assign n9921 = ~n15214 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n9194 = ~n9839 & ~n9193;
  assign n10137 = ~n15793 & ~n10141;
  assign n10471 = ~n10470 & ~n10608;
  assign n9868 = ~n15214 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n15203 = ~n15214 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n12311 = ~n10493 | ~n10492;
  assign n9987 = ~n15214 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n16471 = ~n16031;
  assign n14655 = ~n10791 | ~n10790;
  assign n10024 = ~n15214 | ~P2_DATAO_REG_25__SCAN_IN;
  assign n11368 = ~n14038 | ~n13753;
  assign n14424 = ~n12681;
  assign n16478 = n10631 ^ P2_IR_REG_20__SCAN_IN;
  assign n10223 = ~n11416 | ~n10222;
  assign n10548 = ~n10533 | ~P2_IR_REG_31__SCAN_IN;
  assign n10115 = ~n10114 | ~n10113;
  assign n10215 = ~n10218;
  assign n10141 = ~n10222;
  assign n15619 = ~n16843 | ~n17073;
  assign n11303 = ~n11302;
  assign n9672 = ~n9671;
  assign n10513 = ~n10532 & ~n10608;
  assign n9682 = ~n9723;
  assign n10212 = ~n10208 | ~n10207;
  assign n17084 = ~n17086 & ~P1_U3084;
  assign n9518 = ~n9513 | ~n9512;
  assign n9560 = ~n9532 & ~n9562;
  assign n10532 = ~n10491 & ~P2_IR_REG_12__SCAN_IN;
  assign n16843 = ~n13503 & ~n17072;
  assign n14836 = ~n17072;
  assign n10637 = ~n10634 | ~P2_IR_REG_21__SCAN_IN;
  assign n10111 = ~n13938 | ~n13753;
  assign n9950 = ~n9980;
  assign n9646 = ~n9645 & ~n9733;
  assign n9642 = ~n9641 | ~SI_14_;
  assign n10208 = ~n10206 | ~P2_IR_REG_26__SCAN_IN;
  assign n9837 = ~n9861;
  assign n9803 = ~n9830;
  assign n9730 = ~n9762;
  assign n10022 = ~n10021 | ~SI_25_;
  assign n9741 = ~n9704 & ~n9703;
  assign n9083 = ~n9080 | ~n9079;
  assign n10010 = n10012 ^ SI_24_;
  assign n10486 = ~n10426 & ~P2_IR_REG_9__SCAN_IN;
  assign n9943 = n9945 ^ SI_22_;
  assign n9086 = ~n9084;
  assign n9631 = n9634 ^ SI_13_;
  assign n11036 = ~n11035 | ~SI_27_;
  assign n10211 = ~n10209;
  assign n9681 = ~n9679 & ~n9678;
  assign n9512 = ~n9514 | ~SI_9_;
  assign n9519 = ~n9523 ^ SI_10_;
  assign n11423 = n9106 ^ P1_IR_REG_28__SCAN_IN;
  assign n9913 = n9915 ^ SI_21_;
  assign n9127 = ~n9125 | ~n9124;
  assign n10064 = ~n10063 | ~SI_26_;
  assign n9120 = ~n9118 | ~P1_IR_REG_31__SCAN_IN;
  assign n9228 = n9230 ^ SI_2_;
  assign n9125 = ~n9122 | ~P1_IR_REG_19__SCAN_IN;
  assign n9514 = ~n9442 | ~n9441;
  assign n9523 = ~n9475 | ~n9474;
  assign n9185 = ~n9184 | ~SI_1_;
  assign n10519 = ~n10499 | ~P2_REG3_REG_12__SCAN_IN;
  assign n9103 = ~n9102 & ~n9101;
  assign n9262 = n9264 ^ SI_3_;
  assign n10426 = ~n10404 | ~n10403;
  assign n11049 = ~n11048 | ~n11047;
  assign n9644 = ~n9602 & ~n9733;
  assign n14094 = ~n11059;
  assign n9090 = ~n9121;
  assign n9371 = ~n11089 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n9918 = ~n11089 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n9948 = ~n11089 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n9442 = ~n11089 | ~P1_DATAO_REG_9__SCAN_IN;
  assign n10017 = ~n11089 & ~n10015;
  assign n9153 = ~n9152 | ~n9151;
  assign n9676 = ~n11089 & ~n9683;
  assign n9677 = n11089 & P1_DATAO_REG_15__SCAN_IN;
  assign n9985 = ~n11089 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n9292 = ~n11089 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n9122 = ~n9121 | ~P1_IR_REG_31__SCAN_IN;
  assign n9528 = ~n11089 & ~n9533;
  assign n9897 = ~n11089 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n9475 = ~n11089 | ~P1_DATAO_REG_10__SCAN_IN;
  assign n9584 = ~n9494 | ~P1_REG3_REG_10__SCAN_IN;
  assign n9728 = ~n11089 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n10047 = ~n11089 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n9264 = ~n9234 | ~n9233;
  assign n9403 = ~n11089 & ~n9408;
  assign n9767 = ~n11089 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n9637 = ~n11089 & ~n9643;
  assign n9100 = ~n9445 | ~n9099;
  assign n9267 = ~n9034 | ~P2_DATAO_REG_4__SCAN_IN;
  assign n9867 = ~n9034 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n9527 = ~n9034 & ~n9526;
  assign n9402 = ~n9034 & ~n10395;
  assign n9729 = ~n9034 | ~P2_DATAO_REG_16__SCAN_IN;
  assign n10048 = ~n9034 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n11090 = ~n9034 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n9534 = ~n9573 & ~n9733;
  assign n9565 = ~n9034 & ~n10494;
  assign n9898 = ~n9034 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n14962 = ~n9034 | ~P2_U3152;
  assign n9768 = ~n9034 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n9291 = ~n9034 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n9986 = ~n9034 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n9286 = ~n9034 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n10480 = ~n10436 | ~P2_REG3_REG_10__SCAN_IN;
  assign n9599 = ~n9034 | ~P2_DATAO_REG_13__SCAN_IN;
  assign n9802 = ~n9034 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n9836 = ~n9034 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n9919 = ~n9034 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n9233 = ~n9034 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n10067 = ~n9034 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n9370 = ~n9034 | ~P2_DATAO_REG_7__SCAN_IN;
  assign n9474 = ~n9034 | ~P2_DATAO_REG_10__SCAN_IN;
  assign n9949 = ~n9034 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n9441 = ~n9034 | ~P2_DATAO_REG_9__SCAN_IN;
  assign n9234 = ~n10016 | ~P1_DATAO_REG_3__SCAN_IN;
  assign n9152 = ~n10016 | ~n9149;
  assign n10124 = ~n9409 & ~n9059;
  assign n9287 = ~n10016 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n9268 = ~n10016 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n10190 = ~n10189 | ~n10199;
  assign n10204 = ~n10200 | ~n10199;
  assign n10200 = n10198 & n10197;
  assign n10289 = ~n10271 | ~n10261;
  assign n9046 = ~n9045 | ~n9300;
  assign n9062 = n9061 & n9060;
  assign n9053 = ~n9049 | ~n9048;
  assign n10180 = ~n10177 | ~n10176;
  assign n9057 = ~n9093 | ~n9054;
  assign n10183 = ~n10182 | ~n10181;
  assign n9164 = ~P1_IR_REG_1__SCAN_IN;
  assign n9163 = ~P1_IR_REG_31__SCAN_IN | ~P1_IR_REG_0__SCAN_IN;
  assign n10214 = ~P2_IR_REG_23__SCAN_IN;
  assign n10312 = ~P2_IR_REG_3__SCAN_IN;
  assign n9085 = ~P1_IR_REG_31__SCAN_IN | ~P1_IR_REG_25__SCAN_IN;
  assign n9050 = ~P1_IR_REG_17__SCAN_IN & ~P1_IR_REG_18__SCAN_IN;
  assign P1_U3084 = ~P1_STATE_REG_SCAN_IN;
  assign n10565 = ~P2_IR_REG_16__SCAN_IN;
  assign n10270 = ~P2_IR_REG_31__SCAN_IN | ~P2_IR_REG_0__SCAN_IN;
  assign P2_U3152 = ~P2_STATE_REG_SCAN_IN;
  assign n12666 = ~n12664 & ~n12663;
  assign n14583 = n9066 ^ P1_IR_REG_29__SCAN_IN;
  assign n10310 = n11632 & n11089;
  assign n16969 = ~n10767 & ~n10781;
  assign n9039 = ~n16478;
  assign n17104 = ~n9271 & ~n14237;
  assign n11061 = ~n10239 ^ P2_IR_REG_30__SCAN_IN;
  assign n17110 = ~n15204 | ~n15203;
  assign n9934 = ~n11416 | ~n9128;
  assign n9072 = ~n9064 ^ P1_IR_REG_30__SCAN_IN;
  assign n12014 = ~n16031 | ~n16491;
  assign n16080 = n16491 & n16472;
  assign n12388 = ~n16070;
  assign n12346 = n16070 ^ n12351;
  assign n16070 = ~n10269 & ~n10268;
  assign n10016 = ~n9113 & ~n9112;
  assign n13250 = ~n10378 & ~n10377;
  assign n9857 = n9853 ^ n17107;
  assign n9851 = ~n16534 | ~n17111;
  assign n9995 = n9991 ^ n17107;
  assign n15214 = n9601;
  assign n9183 = ~n10224 | ~n9034;
  assign n16006 = ~n15914 ^ n14506;
  assign n14147 = ~n16650;
  assign n10918 = ~n13265 ^ n11296;
  assign n10950 = n14261 ^ n11318;
  assign n10941 = n16188 ^ n11318;
  assign n15829 = ~n15945 | ~n15709;
  assign n9531 = ~n9530;
  assign n13204 = ~n10918 | ~n10919;
  assign n11267 = n16392 ^ n11296;
  assign n10245 = ~n11061;
  assign n15461 = ~n16382;
  assign n10587 = ~n10586 | ~n14424;
  assign n10393 = ~n13265 | ~n13017;
  assign n9750 = ~n16693 | ~n17111;
  assign n9994 = ~n9996;
  assign n9826 = n9822 ^ n17107;
  assign n9820 = ~n14605 | ~n17111;
  assign n9752 = ~n17107;
  assign n9601 = ~n9170 & ~n9034;
  assign n9774 = ~n9170 | ~n14627;
  assign n11245 = ~n11244;
  assign n10476 = ~n10245 & ~n10244;
  assign n10567 = ~n10586 | ~n14425;
  assign n10551 = ~n15258 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n10535 = ~n13535 | ~n10586;
  assign n10375 = ~n13032 | ~n12646;
  assign n12006 = n10720 | n10719;
  assign n9965 = ~n9967;
  assign n9859 = ~n9857;
  assign n12046 = ~n9656;
  assign n16079 = ~n16072 & ~n16071;
  assign n16273 = ~n16272;
  assign n16061 = ~n16308;
  assign n16729 = ~n16543;
  assign n16450 = ~n16449 | ~n16461;
  assign n15709 = ~n15546 & ~n15942;
  assign n11159 = ~n15928;
  assign n15104 = ~n11187 & ~n15926;
  assign n10628 = ~n10989 | ~n16067;
  assign n16143 = ~n12890 | ~n12687;
  assign n10276 = ~n15371 & ~n11487;
  assign n9174 = ~n12629 | ~n17111;
  assign n9770 = ~n12680;
  assign n9121 = ~n9092 | ~n9573;
  assign n9689 = ~n9684;
  assign n9515 = ~SI_9_;
  assign n9526 = ~P1_DATAO_REG_11__SCAN_IN;
  assign n9513 = ~n9440;
  assign n11298 = ~n16048 ^ n11296;
  assign n10904 = ~n12890 & ~n10888;
  assign n11239 = ~n15138;
  assign n11244 = n16366 ^ n11296;
  assign n10901 = ~n10899;
  assign n13556 = ~n13555 | ~n13554;
  assign n11213 = ~n14510 ^ n11296;
  assign n10555 = ~n11804 | ~P2_REG2_REG_15__SCAN_IN;
  assign n10539 = ~n9035 | ~n13997;
  assign n10540 = ~n11804 | ~P2_REG2_REG_14__SCAN_IN;
  assign n11804 = n10476;
  assign n13865 = ~n13874 ^ n13864;
  assign n10299 = ~n15371 & ~n10298;
  assign n10886 = ~n16472 & ~n16491;
  assign n15371 = ~n11632 | ~n9034;
  assign n15492 = ~n16392 ^ n15468;
  assign n15278 = ~n15479 ^ n16018;
  assign n11116 = ~n11115 ^ n11185;
  assign n10672 = ~n11111 ^ n11112;
  assign n10998 = n16067 ^ n10997;
  assign n12993 = ~n10358 & ~n10357;
  assign n10490 = ~n10487 | ~P2_IR_REG_12__SCAN_IN;
  assign n9661 = ~n16678 | ~n17111;
  assign n9967 = n9964 ^ n17107;
  assign n9962 = ~n15159 | ~n17111;
  assign n10081 = ~n16853 | ~n17104;
  assign n9878 = ~n15088 | ~n17111;
  assign n9881 = ~n15088 | ~n17104;
  assign n10032 = ~n10028 ^ n17107;
  assign n10027 = ~n16781 | ~n17111;
  assign n10030 = ~n16781 | ~n17104;
  assign n9786 = ~n16717 | ~n17111;
  assign n9993 = ~n15697 | ~n17104;
  assign n9931 = ~n15512 | ~n17111;
  assign n9553 = ~n13837 | ~n17111;
  assign n10058 = ~n10054 ^ n17107;
  assign n10053 = ~n16787 | ~n17111;
  assign n10056 = ~n16787 | ~n17104;
  assign n9314 = ~P1_REG3_REG_3__SCAN_IN;
  assign n9137 = ~n9136 & ~n9135;
  assign n11759 = ~n11974;
  assign n14591 = ~n14666;
  assign n12451 = ~n12763;
  assign n15635 = n15734 ^ n17021;
  assign n16531 = ~n16534;
  assign n14215 = ~n16680;
  assign n13587 = ~n13583 | ~n10774;
  assign n13583 = ~n16994 ^ n13952;
  assign n9237 = ~n9227 & ~n9226;
  assign n10014 = ~n10011 | ~n10010;
  assign n9896 = ~n9893 | ~n9892;
  assign n9763 = ~n9761;
  assign n9678 = ~SI_15_;
  assign n9563 = ~n9562;
  assign n9471 = n9514 ^ SI_9_;
  assign n10383 = ~n10382 | ~n10381;
  assign n11323 = ~n15777 ^ n11320;
  assign n11320 = ~n11319 ^ n11318;
  assign n10439 = ~n9035 | ~n10438;
  assign n10440 = ~n11803 | ~P2_REG0_REG_9__SCAN_IN;
  assign n11228 = ~n14893 | ~n14891;
  assign n15010 = n16337 ^ n11296;
  assign n11254 = ~n11251 & ~n15523;
  assign n11252 = ~n15524;
  assign n11264 = ~n11266;
  assign n11265 = ~n11267;
  assign n14433 = ~n11017;
  assign n16285 = ~n16277;
  assign n11193 = ~n11804 | ~P2_REG2_REG_25__SCAN_IN;
  assign n11166 = ~n11807 | ~P2_REG1_REG_24__SCAN_IN;
  assign n11153 = ~n11807 | ~P2_REG1_REG_23__SCAN_IN;
  assign n11118 = ~n11807 | ~P2_REG1_REG_22__SCAN_IN;
  assign n11100 = ~n11807 | ~P2_REG1_REG_21__SCAN_IN;
  assign n10677 = ~n11807 | ~P2_REG1_REG_20__SCAN_IN;
  assign n10251 = ~n11803 | ~P2_REG0_REG_19__SCAN_IN;
  assign n10242 = ~n11804 | ~P2_REG2_REG_19__SCAN_IN;
  assign n10622 = ~n9035 | ~n14505;
  assign n10621 = ~n11804 | ~P2_REG2_REG_18__SCAN_IN;
  assign n10619 = ~n11807 | ~P2_REG1_REG_18__SCAN_IN;
  assign n10597 = ~n9035 | ~n11007;
  assign n10596 = ~n11804 | ~P2_REG2_REG_17__SCAN_IN;
  assign n10592 = ~n11807 | ~P2_REG1_REG_17__SCAN_IN;
  assign n10573 = ~n11804 | ~P2_REG2_REG_16__SCAN_IN;
  assign n12307 = ~P2_REG2_REG_11__SCAN_IN ^ n12306;
  assign n13875 = ~n13874 ^ n13873;
  assign n14567 = ~n14875 ^ n14874;
  assign n14881 = n14880 ^ n14879;
  assign n15051 = ~n16337 ^ n15043;
  assign n14701 = ~n10729;
  assign n14102 = ~n14070 ^ n14063;
  assign n10473 = ~n12306 | ~n10586;
  assign n13696 = n15989 ^ n13695;
  assign n13740 = n15989 ^ n13690;
  assign n10362 = ~n10361 | ~n10360;
  assign n16038 = ~n16472;
  assign n10281 = ~n16070 | ~n16090;
  assign n14703 = ~n15914 | ~n16502;
  assign n14116 = n16001 ^ n14048;
  assign n14119 = ~n14117 | ~n16500;
  assign n14083 = ~n14081 | ~n16500;
  assign n14014 = ~n14012 | ~n16500;
  assign n13399 = n13173 ^ n13172;
  assign n10531 = ~P2_IR_REG_13__SCAN_IN;
  assign n10547 = ~P2_IR_REG_14__SCAN_IN;
  assign n9902 = ~n16739 | ~n17111;
  assign n9905 = ~n16739 | ~n17104;
  assign n14146 = ~n16666;
  assign n10000 = ~n9999;
  assign n9758 = ~n9757;
  assign n9810 = n9809 & n9808;
  assign n9808 = ~n15214 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n9848 = ~n9846 | ~n9845;
  assign n12041 = ~n9038;
  assign n11675 = ~n9612;
  assign n9614 = ~n9037 | ~P1_REG2_REG_13__SCAN_IN;
  assign n9071 = ~n14583;
  assign n9612 = ~n9656;
  assign n9215 = ~n9038 | ~n9314;
  assign n9214 = n9612 & P1_REG1_REG_3__SCAN_IN;
  assign n9144 = ~n9612 | ~P1_REG1_REG_1__SCAN_IN;
  assign n9143 = n9544 & P1_REG2_REG_1__SCAN_IN;
  assign n9074 = ~n9612 | ~P1_REG1_REG_0__SCAN_IN;
  assign n9075 = ~n9544 | ~P1_REG2_REG_0__SCAN_IN;
  assign n9069 = ~n12043 & ~n9068;
  assign n11691 = ~n11512 | ~n11511;
  assign n14834 = ~n14832 ^ n14831;
  assign n15198 = ~n15214 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n9605 = n9604 & n9603;
  assign n9603 = ~n9170 | ~n12983;
  assign n15743 = ~n15742 | ~n15741;
  assign n14277 = ~n14311 | ~n15791;
  assign n14371 = n14356 ^ n14355;
  assign n14294 = n17000 ^ n14280;
  assign n14391 = n16998 ^ n14216;
  assign n13657 = n16994 ^ n13960;
  assign n13407 = n13342 ^ n16991;
  assign n13342 = ~n13341 | ~n13590;
  assign n13166 = ~n13127 & ~n13126;
  assign n13425 = ~n13377 | ~n13376;
  assign n17073 = n9091 ^ P1_IR_REG_20__SCAN_IN;
  assign n9773 = ~n9772 | ~n9771;
  assign n14627 = n9805 ^ n9804;
  assign n9481 = ~P1_IR_REG_10__SCAN_IN;
  assign n9446 = ~n9445 | ~n9444;
  assign n10477 = ~n10476 | ~P2_REG2_REG_11__SCAN_IN;
  assign n14895 = P2_REG3_REG_21__SCAN_IN ^ n11119;
  assign n11025 = ~n11207 ^ n11024;
  assign n11024 = ~n11208 ^ n11205;
  assign n15439 = P2_REG3_REG_24__SCAN_IN ^ n11190;
  assign n10515 = ~n12919 | ~n10586;
  assign n13653 = ~n13651 | ~n13650;
  assign n13650 = ~n15527 | ~n13649;
  assign n13017 = ~n13288;
  assign n14425 = n10566 ^ n10565;
  assign n13886 = ~n13885 | ~n13884;
  assign n13734 = ~n13733 | ~n13894;
  assign n13715 = ~n13714 | ~n13713;
  assign n13496 = ~n13495 | ~n14993;
  assign n14850 = ~n15088;
  assign n14849 = ~n14848 ^ n14847;
  assign n14860 = ~n14859 | ~n14858;
  assign n14859 = ~n16548 | ~n15578;
  assign n13861 = ~n13852 | ~n13851;
  assign n14826 = n14824 ^ n14823;
  assign n14823 = ~n14822 | ~n14821;
  assign n14693 = n17010 ^ n14747;
  assign n14680 = ~n14688 | ~n15762;
  assign n14852 = ~P1_REG3_REG_19__SCAN_IN ^ n9870;
  assign n14502 = ~n14604 ^ n14484;
  assign n14318 = ~n14286 ^ n14481;
  assign n9082 = ~n9081;
  assign n16091 = ~n16099 | ~n16087;
  assign n16106 = ~n16105 | ~n16104;
  assign n16102 = ~n16101 | ~n16100;
  assign n16145 = ~n16114 & ~n16151;
  assign n16194 = ~n16174 & ~n16173;
  assign n16206 = ~n16194;
  assign n16219 = ~n16191 & ~n16190;
  assign n16217 = ~n16216 | ~n16215;
  assign n16238 = ~n16228 | ~n16227;
  assign n16627 = ~n16621 | ~n16620;
  assign n16259 = ~n16250 & ~n16249;
  assign n16275 = ~n16274 & ~n16273;
  assign n16656 = ~n16648 | ~n16647;
  assign n16648 = ~n16645 | ~n16644;
  assign n16673 = ~n16672 | ~n16671;
  assign n16684 = ~n16677 & ~n16676;
  assign n16698 = ~n16686 | ~n16685;
  assign n16312 = ~n16317 | ~n16311;
  assign n16709 = ~n16691 | ~n16690;
  assign n16708 = ~n16695 & ~n16694;
  assign n16705 = ~n16699 | ~n16698;
  assign n16707 = ~n16697 & ~n16696;
  assign n16696 = ~n16709 & ~n16708;
  assign n16697 = ~n16699 & ~n16698;
  assign n16329 = ~n16328;
  assign n16731 = ~n16727 | ~n16726;
  assign n16726 = ~n16725 | ~n16724;
  assign n16727 = ~n16721 | ~n16720;
  assign n16545 = ~n16729 | ~n16544;
  assign n15901 = ~n15897 | ~n15896;
  assign n15897 = ~n15893 | ~n15892;
  assign n15893 = ~n15891 | ~n15890;
  assign n16356 = ~n16355 | ~n16354;
  assign n16354 = ~n16353 | ~n16352;
  assign n16372 = ~n16369 | ~n16368;
  assign n16749 = ~n16748 | ~n16751;
  assign n16748 = ~n16747 & ~n16746;
  assign n16746 = ~n16745 | ~n16744;
  assign n16759 = ~n16752 | ~n16751;
  assign n16752 = ~n16750;
  assign n16758 = ~n16757 | ~n16756;
  assign n16757 = ~n16754 | ~n16753;
  assign n16756 = ~n16755 | ~n16866;
  assign n15915 = ~n16305 | ~n15912;
  assign n15912 = ~n15911 | ~n15910;
  assign n15910 = ~n15909 | ~n15908;
  assign n16387 = ~n16385;
  assign n16374 = ~n16373;
  assign n16399 = ~n16398;
  assign n16770 = ~n16767 | ~n16766;
  assign n16767 = ~n16765 | ~n17051;
  assign n16765 = ~n16764 & ~n16865;
  assign n16796 = ~n16794 | ~n16793;
  assign n16523 = ~n16861;
  assign n15931 = ~n15929 | ~n15928;
  assign n15925 = ~n15923 | ~n15922;
  assign n16415 = ~n16414 & ~n16461;
  assign n17046 = ~n16942 & ~n16941;
  assign n16813 = ~n16864 | ~n16947;
  assign n16429 = ~n16428 | ~n16427;
  assign n16442 = ~n16439;
  assign n16873 = ~n16872 | ~n16871;
  assign n16872 = ~n16868 | ~n16867;
  assign n16859 = ~n16856 & ~n16855;
  assign n16819 = ~n16818 | ~n16817;
  assign n16817 = ~n16816 | ~n16815;
  assign n16818 = ~n16813 | ~n16843;
  assign n16815 = ~n16814 & ~n16843;
  assign n16820 = ~n16812 & ~n16811;
  assign n16811 = ~n16810 | ~n16809;
  assign n16812 = ~n16808;
  assign n16785 = ~n16810 & ~n16809;
  assign n16803 = ~n16801 | ~n16688;
  assign n17013 = ~n17012 | ~n17011;
  assign n15941 = ~n15939 | ~n15938;
  assign n15918 = ~n14766;
  assign n15899 = ~n13717;
  assign n17055 = ~n17054 | ~n17053;
  assign n17053 = ~n17052 | ~n17051;
  assign n17052 = ~n17050 | ~n17049;
  assign n17049 = ~n17048 | ~n17047;
  assign n16829 = ~n17063 | ~n16843;
  assign n16949 = ~n17056 & ~n16948;
  assign n17005 = ~n16878;
  assign n9055 = ~P1_IR_REG_20__SCAN_IN;
  assign n9516 = ~n9514;
  assign n10935 = n16205 ^ n11296;
  assign n10395 = ~P1_DATAO_REG_8__SCAN_IN;
  assign n10923 = n16160 ^ n11296;
  assign n10947 = n16229 ^ n11318;
  assign n10928 = n16176 ^ n11296;
  assign n16026 = ~n16449 ^ n16452;
  assign n16028 = n15968 ^ n15967;
  assign n16453 = ~n16452 | ~n16461;
  assign n16251 = ~n13982;
  assign n10297 = ~n10310 | ~n11545;
  assign n16410 = ~n16427;
  assign n11188 = ~n15104 | ~n15928;
  assign n11084 = ~n15914;
  assign n10667 = ~n15907;
  assign n16062 = ~n15884;
  assign n16063 = ~n15883;
  assign n16243 = ~n16247;
  assign n13689 = ~n15892;
  assign n16165 = ~n16148;
  assign n16166 = ~n16135;
  assign n16150 = ~n16110;
  assign n10186 = ~P2_IR_REG_20__SCAN_IN;
  assign n10187 = ~P2_IR_REG_19__SCAN_IN;
  assign n17065 = ~n17063 | ~n17062;
  assign n16841 = ~n17036;
  assign n17029 = ~n17063 ^ n17062;
  assign n9571 = ~P2_DATAO_REG_12__SCAN_IN;
  assign n9533 = ~P2_DATAO_REG_11__SCAN_IN;
  assign n16628 = ~n13280;
  assign n9408 = ~P2_DATAO_REG_8__SCAN_IN;
  assign n9775 = ~n15214 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n14133 = ~n14216;
  assign n16892 = ~n13114 | ~n13371;
  assign n10787 = ~n12372;
  assign n12373 = ~n16979;
  assign n9094 = ~n9093;
  assign n9098 = ~n9092;
  assign n9725 = ~n9680 & ~SI_15_;
  assign n9404 = ~SI_8_;
  assign n10382 = ~n15258 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n10494 = ~P1_DATAO_REG_12__SCAN_IN;
  assign n11019 = ~n11014;
  assign n11218 = ~n15914 ^ n11296;
  assign n11229 = ~n14891;
  assign n10944 = ~n10941;
  assign n10897 = ~n16073 | ~n12806;
  assign n13021 = ~n10913 | ~n10914;
  assign n10521 = ~n9035 | ~n13924;
  assign n10522 = ~n11803 | ~P2_REG0_REG_13__SCAN_IN;
  assign n10523 = ~n11804 | ~P2_REG2_REG_13__SCAN_IN;
  assign n10504 = ~n9035 | ~n10503;
  assign n10505 = ~n9033 | ~P2_REG0_REG_12__SCAN_IN;
  assign n10506 = ~n11804 | ~P2_REG2_REG_12__SCAN_IN;
  assign n10461 = ~n9035 | ~n10460;
  assign n10462 = ~n11803 | ~P2_REG0_REG_10__SCAN_IN;
  assign n10464 = ~n11807 | ~P2_REG1_REG_10__SCAN_IN;
  assign n12064 = ~n11940 | ~n12060;
  assign n11934 = ~n12135;
  assign n12582 = P2_REG2_REG_12__SCAN_IN ^ n12311;
  assign n12586 = ~n12919;
  assign n12920 = P2_REG2_REG_13__SCAN_IN ^ n12586;
  assign n13536 = ~P2_REG2_REG_14__SCAN_IN ^ n13535;
  assign n10957 = ~P2_REG3_REG_14__SCAN_IN;
  assign n11327 = ~n15849;
  assign n15466 = ~n15940;
  assign n15467 = ~n15942;
  assign n14566 = ~n14876;
  assign n10534 = ~n15258 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n10472 = ~n15258 | ~P1_DATAO_REG_11__SCAN_IN;
  assign n10656 = ~n13184 | ~n16161;
  assign n10364 = ~P2_REG3_REG_6__SCAN_IN;
  assign n10355 = ~n10354 | ~n10353;
  assign n15833 = ~n15831 ^ n16024;
  assign n15708 = ~n15706 & ~n15705;
  assign n15777 = ~n11308 | ~n11307;
  assign n15712 = ~n15711 ^ n16022;
  assign n15710 = ~n15828;
  assign n15544 = ~n15945;
  assign n15550 = ~n16488;
  assign n15548 = n16030 ^ n15709;
  assign n15552 = ~n15868 | ~n15549;
  assign n15270 = ~n15936;
  assign n15271 = ~n15938;
  assign n11189 = n15275 ^ n16016;
  assign n15105 = ~n15104 ^ n16014;
  assign n15029 = n15028 ^ n16012;
  assign n11106 = ~n15920;
  assign n11107 = ~n15922;
  assign n14771 = n16008 ^ n14770;
  assign n14702 = n15914 ^ n11134;
  assign n10729 = n11111 ^ n11086;
  assign n10626 = ~n15881;
  assign n10625 = ~n16293;
  assign n10852 = ~n16003 ^ n10851;
  assign n14054 = n14053 ^ n16001;
  assign n14005 = ~n13994 ^ n13993;
  assign n13983 = ~n13985 | ~n13982;
  assign n13908 = ~n15994 ^ n13907;
  assign n13730 = ~n15992 ^ n13729;
  assign n10419 = ~n16164;
  assign n10652 = ~n12694 | ~n12695;
  assign n10649 = ~n12594 | ~n10647;
  assign n12900 = ~n16090 | ~n16071;
  assign n10218 = ~n10213 & ~n10608;
  assign n10447 = ~n10486;
  assign n10396 = ~P2_IR_REG_6__SCAN_IN;
  assign n17135 = ~n16853;
  assign n9430 = ~n9429 | ~n9428;
  assign n15690 = ~P1_REG3_REG_25__SCAN_IN;
  assign n9465 = ~n9461 ^ n17107;
  assign n9628 = n9591 ^ n9752;
  assign n12774 = ~n12819;
  assign n9356 = ~n12779;
  assign n11683 = ~n11521 | ~n11520;
  assign n11696 = ~n11691 | ~n11690;
  assign n11724 = ~P1_REG3_REG_9__SCAN_IN;
  assign n13462 = ~n13461 ^ n13759;
  assign n13761 = ~n13771 | ~n13759;
  assign n14336 = ~P1_REG3_REG_17__SCAN_IN;
  assign n14827 = ~P1_REG3_REG_19__SCAN_IN;
  assign n14236 = ~n14159 | ~n14158;
  assign n11981 = ~P1_REG3_REG_11__SCAN_IN;
  assign n9604 = ~n15214 | ~P2_DATAO_REG_13__SCAN_IN;
  assign n11524 = ~P1_REG3_REG_7__SCAN_IN;
  assign n9372 = ~n11626;
  assign n9315 = ~P1_REG3_REG_5__SCAN_IN | ~P1_REG3_REG_4__SCAN_IN;
  assign n15163 = n14655 & n17072;
  assign n15593 = n15633 ^ n17054;
  assign n15393 = ~n16864;
  assign n15300 = ~n15391 ^ n17024;
  assign n15170 = n17018 ^ n15305;
  assign n15155 = ~n15297 ^ n17018;
  assign n14969 = ~n17016 ^ n15153;
  assign n14909 = n17014 ^ n14967;
  assign n14732 = ~n17012 ^ n14907;
  assign n14670 = n17010 ^ n14730;
  assign n14593 = ~n14592 ^ n14608;
  assign n14471 = n14590 ^ n14484;
  assign n14349 = ~n14348 ^ n14354;
  assign n14150 = ~n14149 ^ n17000;
  assign n14229 = ~n14228 ^ n16998;
  assign n13965 = ~n16996;
  assign n13782 = n16989 ^ n13781;
  assign n13596 = ~n13595 | ~n13594;
  assign n13592 = n13591 & n13590;
  assign n13792 = ~n13837;
  assign n9293 = ~n11537;
  assign n9332 = ~n11474;
  assign n10021 = ~n10020;
  assign n9984 = ~n9981 | ~n9980;
  assign n9641 = ~n9640;
  assign n9673 = ~n9636 & ~n9635;
  assign n9636 = ~n9633 & ~n9632;
  assign n9567 = ~SI_12_;
  assign n9559 = ~n9525 | ~n9524;
  assign n9525 = ~n9522 | ~n9521;
  assign n9529 = ~SI_11_;
  assign n9445 = ~n9409;
  assign n9439 = ~n9401 | ~n9400;
  assign n9397 = n9399 ^ SI_7_;
  assign n9365 = n9367 ^ SI_6_;
  assign n9330 = n9288 ^ SI_5_;
  assign n9154 = ~P2_DATAO_REG_1__SCAN_IN;
  assign n9110 = ~n10810 | ~n9109;
  assign n15138 = ~n15115 ^ n11296;
  assign n10481 = ~n9035 | ~n13654;
  assign n10482 = ~n11807 | ~P2_REG1_REG_11__SCAN_IN;
  assign n10478 = ~n9033 | ~P2_REG0_REG_11__SCAN_IN;
  assign n12406 = n10899 ^ n10900;
  assign n14638 = n11218 ^ n11219;
  assign n11300 = ~n11297;
  assign n11299 = ~n11298;
  assign n13297 = ~n10922 | ~n13203;
  assign n12325 = n10890 ^ n10891;
  assign n16076 = ~n16073;
  assign n14891 = ~n14997 ^ n11296;
  assign n15524 = n16378 ^ n11296;
  assign n10514 = ~n15258 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n14256 = ~n14255 ^ n14254;
  assign n10479 = ~P2_REG3_REG_11__SCAN_IN;
  assign n12415 = n10897 ^ n10895;
  assign n11209 = ~n11208;
  assign n11215 = ~n11214;
  assign n11216 = ~n11213;
  assign n16392 = ~n11256 & ~n11255;
  assign n11314 = ~n11804 | ~P2_REG2_REG_28__SCAN_IN;
  assign n11274 = n11061 | n10244;
  assign n11276 = ~n11272 | ~n11271;
  assign n15564 = P2_REG3_REG_27__SCAN_IN ^ n11311;
  assign n11261 = ~n11804 | ~P2_REG2_REG_26__SCAN_IN;
  assign n11192 = ~n11807 | ~P2_REG1_REG_25__SCAN_IN;
  assign n10561 = ~n10556 | ~n10555;
  assign n10560 = ~n10559 | ~n10558;
  assign n10543 = ~n10542 | ~n10541;
  assign n10324 = ~n10323 | ~n10322;
  assign n10254 = ~n10412 | ~P2_REG3_REG_0__SCAN_IN;
  assign n11803 = ~n11274;
  assign n12129 = ~n12126 | ~n12127;
  assign n12123 = ~n12121 | ~n12120;
  assign n12913 = P2_REG1_REG_13__SCAN_IN ^ n12586;
  assign n13530 = ~P2_REG1_REG_14__SCAN_IN ^ n13535;
  assign n11662 = ~n14404;
  assign n16501 = ~n16503 ^ n15846;
  assign n15776 = n15777 ^ n15723;
  assign n15824 = ~n15777;
  assign n15659 = n15565 ^ n16048;
  assign n15473 = ~P2_REG3_REG_26__SCAN_IN ^ n11270;
  assign n15478 = ~n15560 ^ n16020;
  assign n15125 = n15114 ^ n15115;
  assign n16337 = ~n11145 & ~n11144;
  assign n14996 = n14997 ^ n11174;
  assign n14809 = n16302 ^ n14783;
  assign n10732 = ~n15847 | ~n14702;
  assign n14458 = n10992 ^ n14510;
  assign n10841 = ~n15720 | ~n10644;
  assign n14117 = n14447 ^ n14082;
  assign n14012 = ~n16247 ^ n14002;
  assign n14011 = ~n14005;
  assign n13932 = ~n15994 ^ n13902;
  assign n13890 = ~n15992 ^ n13719;
  assign n13438 = n15981 ^ n13250;
  assign n10641 = ~n16038 | ~n16491;
  assign n15547 = ~n16469 & ~n10671;
  assign n12008 = ~n10718 & ~n11611;
  assign n16500 = ~n14995;
  assign n15775 = ~n15823 ^ n16022;
  assign n15658 = ~n16030 ^ n15706;
  assign n15336 = n15462 ^ n16018;
  assign n15027 = ~n15024;
  assign n14808 = ~n16008 ^ n14768;
  assign n14459 = ~n14510 | ~n16502;
  assign n14457 = n16067 ^ n10989;
  assign n14204 = ~n16056 | ~n16502;
  assign n10846 = ~n10845 | ~n16500;
  assign n10845 = ~n16056 | ~n10844;
  assign n14203 = n16003 ^ n10840;
  assign n15657 = ~n15335;
  assign n14072 = n14071 ^ n14070;
  assign n13893 = ~n13722 | ~n13911;
  assign n13892 = n13890 & n14993;
  assign n13619 = ~n13618 | ~n13617;
  assign n13620 = ~n13616 | ~n13615;
  assign n13628 = ~n13624 | ~n13623;
  assign n13626 = ~n15988 ^ n13625;
  assign n13743 = ~n13742 | ~n13741;
  assign n13495 = n15986 ^ n13312;
  assign n13397 = ~n13396 | ~n13395;
  assign n14993 = ~n16498;
  assign n10883 = ~n16468 | ~n16472;
  assign n12021 = ~n12008 & ~n12007;
  assign n14961 = ~n10240 | ~n10238;
  assign n10238 = ~P2_IR_REG_29__SCAN_IN;
  assign n16487 = n10230 ^ P2_IR_REG_27__SCAN_IN;
  assign n10191 = ~P2_IR_REG_22__SCAN_IN;
  assign n10636 = ~n10635 | ~P2_IR_REG_31__SCAN_IN;
  assign n10493 = ~n10490 | ~n10489;
  assign n10271 = ~P2_IR_REG_1__SCAN_IN;
  assign n11487 = ~P1_DATAO_REG_1__SCAN_IN;
  assign n9361 = ~n9360 | ~n12779;
  assign n12749 = ~n9392 | ~n9393;
  assign n12748 = ~n9395 | ~n9394;
  assign n16524 = ~n10069 | ~n10068;
  assign n9243 = ~n9242 & ~n9241;
  assign n9856 = ~n9858;
  assign n17111 = ~n9934;
  assign n12822 = ~n12435;
  assign n16689 = ~n16693;
  assign n9793 = ~n9792;
  assign n9794 = ~n9791;
  assign n9997 = ~n9995;
  assign n12663 = n9277 ^ n9278;
  assign n13274 = n9465 ^ n9466;
  assign n9624 = ~n9623;
  assign n9625 = ~n9622;
  assign n13594 = ~n13783;
  assign n13961 = ~n13855;
  assign n9554 = ~n9556;
  assign n9557 = ~n9555;
  assign n10861 = n10751 & n10750;
  assign n10136 = ~n10147 | ~n13968;
  assign n12780 = ~n9357;
  assign n12781 = ~n9357 | ~n9356;
  assign n15809 = n10058 ^ n10057;
  assign n17079 = ~n17078;
  assign n10039 = ~n10036 | ~n10035;
  assign n10007 = ~n10004 | ~n10003;
  assign n9977 = ~n9974 | ~n9973;
  assign n9959 = ~n9956 | ~n9955;
  assign n9928 = ~n9925 | ~n9924;
  assign n9889 = ~n9886 | ~n9885;
  assign n9875 = ~n9872 | ~n9871;
  assign n9817 = ~n9814 | ~n9813;
  assign n9252 = ~n9248 | ~n9247;
  assign n9198 = n9612 & P1_REG1_REG_2__SCAN_IN;
  assign n11516 = ~n11557 | ~n11446;
  assign n11512 = ~n11510 | ~n11509;
  assign n14333 = ~n14833;
  assign n13452 = P1_REG2_REG_14__SCAN_IN ^ n12986;
  assign n13455 = ~n13770 ^ n13461;
  assign n13773 = ~n13771 | ~n13770;
  assign n14325 = ~n14825;
  assign n15764 = ~n16520;
  assign n17127 = ~n17110;
  assign n15621 = ~n16524 ^ n15609;
  assign n15610 = P1_REG3_REG_27__SCAN_IN ^ n10152;
  assign n15812 = P1_REG3_REG_26__SCAN_IN ^ n10070;
  assign n15323 = ~n16782 ^ n15312;
  assign n15691 = ~P1_REG3_REG_25__SCAN_IN ^ n10034;
  assign n15585 = P1_REG3_REG_24__SCAN_IN ^ n10002;
  assign n15510 = P1_REG3_REG_23__SCAN_IN ^ n9972;
  assign n14977 = ~n14926 & ~n14925;
  assign n14925 = ~n16741;
  assign n14930 = n14981 ^ n14980;
  assign n15231 = ~n14981;
  assign n15230 = P1_REG3_REG_22__SCAN_IN ^ n9954;
  assign n14753 = ~n16738 ^ n14916;
  assign n14688 = n14748 ^ n14739;
  assign n14495 = n14598 ^ n14797;
  assign n16728 = ~n14797;
  assign n14311 = ~n16716 ^ n14476;
  assign n16712 = ~n16716;
  assign n16687 = ~n16692;
  assign n14217 = ~n16657;
  assign n15671 = ~n15748 ^ n17021;
  assign n15639 = ~n15638 | ~n15637;
  assign n15620 = n15644 ^ n17054;
  assign n15421 = n15601 ^ n17026;
  assign n15322 = ~n17024 ^ n15401;
  assign n15068 = n17016 ^ n15158;
  assign n14931 = ~n14981 | ~n15793;
  assign n14754 = ~n16738 | ~n15793;
  assign n14689 = ~n14748 | ~n15793;
  assign n14656 = n14683 ^ n14608;
  assign n14478 = ~n14495 | ~n15791;
  assign n15185 = ~n12281 | ~n17073;
  assign n13601 = ~n13587 | ~n13586;
  assign n13358 = ~n13356 | ~n13355;
  assign n13160 = ~n16985 ^ n13222;
  assign n9116 = ~n9170 | ~P1_IR_REG_0__SCAN_IN;
  assign n12180 = ~n10122 | ~n11368;
  assign n12182 = n12158 & n12157;
  assign n15254 = n11066 ^ SI_30_;
  assign n14574 = n11049 ^ SI_29_;
  assign n11306 = ~n11044 | ~n11302;
  assign n11845 = n9108 ^ P1_IR_REG_27__SCAN_IN;
  assign n10065 = ~n10062 | ~n10061;
  assign n10119 = n9087 ^ P1_IR_REG_26__SCAN_IN;
  assign n14095 = n10062 ^ n10049;
  assign n10049 = ~n10061;
  assign n9084 = ~n9081 & ~n9733;
  assign n13943 = n10043 ^ n10042;
  assign n9078 = ~P1_IR_REG_24__SCAN_IN;
  assign n9081 = ~n10130 & ~P1_IR_REG_24__SCAN_IN;
  assign n13508 = ~n9944 ^ n9943;
  assign n17037 = ~n9104 & ~n9103;
  assign n9104 = ~n9118;
  assign n11096 = ~n9914 ^ n9913;
  assign n9865 = ~n9862 | ~n9861;
  assign n17072 = ~n9127 | ~n9126;
  assign n13065 = ~n9862 ^ n9837;
  assign n12842 = ~n9831 ^ n9803;
  assign n12680 = n9769 ^ n9796;
  assign n14328 = n9734 ^ P1_IR_REG_16__SCAN_IN;
  assign n12427 = ~n9761 ^ n9730;
  assign n12295 = n9724 ^ n9682;
  assign n12146 = n9673 ^ n9671;
  assign n12077 = ~n9633 ^ n9631;
  assign n9572 = ~P1_IR_REG_11__SCAN_IN;
  assign n11995 = ~n9595 ^ n9594;
  assign n11822 = n9559 ^ n9560;
  assign n11831 = ~n9476 ^ n9519;
  assign n11721 = n9479 ^ P1_IR_REG_9__SCAN_IN;
  assign n11778 = n9472 ^ n9471;
  assign n11693 = n9410 ^ P1_IR_REG_8__SCAN_IN;
  assign n9410 = ~n9409 | ~P1_IR_REG_31__SCAN_IN;
  assign n11739 = ~n9439 ^ n9438;
  assign n11626 = ~n9398 ^ n9397;
  assign n11537 = ~n9366 ^ n9365;
  assign n11474 = ~n9331 ^ n9330;
  assign n9281 = n9283 ^ SI_4_;
  assign n10417 = ~n10416 | ~n10415;
  assign n10418 = ~n10414 | ~n10413;
  assign n10952 = ~n10972 ^ n10973;
  assign n15142 = P2_REG3_REG_23__SCAN_IN ^ n11167;
  assign n15141 = ~n15140 ^ n15139;
  assign n15139 = n15138 ^ n15137;
  assign n13524 = ~n13523 | ~n13522;
  assign n14639 = ~n14638 ^ n14637;
  assign n14647 = ~n14646 | ~n14645;
  assign n10443 = ~n10442 | ~n10441;
  assign n14894 = ~n14893 ^ n14892;
  assign n14892 = n14891 ^ n14890;
  assign n14900 = ~n15867 | ~n16321;
  assign n15529 = P2_REG3_REG_25__SCAN_IN ^ n11259;
  assign n15528 = ~n15526 ^ n15525;
  assign n15525 = n15524 ^ n15523;
  assign n14444 = ~n14443 ^ n14442;
  assign n14442 = ~n14441 | ~n14440;
  assign n15438 = ~n15437 ^ n15436;
  assign n13561 = ~n13560 | ~n13559;
  assign n14780 = P2_REG3_REG_20__SCAN_IN ^ n11101;
  assign n14719 = ~n14718 ^ n14717;
  assign n14724 = ~n15867 | ~n16298;
  assign n10964 = ~n10963;
  assign n15040 = P2_REG3_REG_22__SCAN_IN ^ n11154;
  assign n15013 = ~n15012 ^ n15011;
  assign n15011 = ~n15010 ^ n15009;
  assign n10268 = ~n10267 | ~n10266;
  assign n14505 = n10620 ^ P2_REG3_REG_18__SCAN_IN;
  assign n14519 = ~n14518 ^ n14517;
  assign n14517 = ~n14516 | ~n14515;
  assign n15527 = ~n10963 & ~n10884;
  assign n10884 = ~n15451 | ~n16039;
  assign n11269 = n11291 ^ n11268;
  assign n15530 = ~n10882 & ~P2_U3152;
  assign n10881 = ~n10880 | ~n10879;
  assign n10981 = ~n10980 ^ n14433;
  assign n11263 = n11258 & n11257;
  assign n11257 = ~n11803 | ~P2_REG0_REG_26__SCAN_IN;
  assign n11194 = ~n9033 | ~P2_REG0_REG_25__SCAN_IN;
  assign n11171 = n11166 & n11165;
  assign n11165 = ~n11803 | ~P2_REG0_REG_24__SCAN_IN;
  assign n11158 = n11153 & n11152;
  assign n11152 = ~n11803 | ~P2_REG0_REG_23__SCAN_IN;
  assign n11117 = ~n9033 | ~P2_REG0_REG_22__SCAN_IN;
  assign n11099 = ~n11803 | ~P2_REG0_REG_21__SCAN_IN;
  assign n10674 = ~n9033 | ~P2_REG0_REG_20__SCAN_IN;
  assign n10243 = ~n11807 | ~P2_REG1_REG_19__SCAN_IN;
  assign n10624 = n10619 & n10618;
  assign n10618 = ~n9033 | ~P2_REG0_REG_18__SCAN_IN;
  assign n10599 = n10592 & n10591;
  assign n10591 = ~n9033 | ~P2_REG0_REG_17__SCAN_IN;
  assign n10575 = n10574 & n10573;
  assign n10576 = n10572 & n10571;
  assign n16230 = ~n16226;
  assign n16189 = ~n16192;
  assign n16195 = ~n13642;
  assign n16177 = ~n16209;
  assign n10390 = n10389 & n10388;
  assign n10391 = n10387 & n10386;
  assign n10373 = n10372 & n10371;
  assign n10374 = n10370 & n10369;
  assign n10344 = n10343 & n10342;
  assign n16116 = ~n12890;
  assign n10308 = ~n10307 | ~n10306;
  assign n10306 = ~n11803 | ~P2_REG0_REG_3__SCAN_IN;
  assign n12273 = ~n10359 ^ P2_IR_REG_6__SCAN_IN;
  assign n12070 = n10380 ^ P2_IR_REG_7__SCAN_IN;
  assign n13543 = ~n13542 | ~n13541;
  assign n14422 = ~n14421 | ~n14420;
  assign n14421 = ~n14419 | ~n11932;
  assign n14569 = ~n14561 | ~n11932;
  assign n14561 = ~n14868 ^ n14867;
  assign n14873 = n14872 ^ n14871;
  assign n15450 = n15961 ^ n15375;
  assign n15382 = n16449 ^ n15374;
  assign n11180 = ~n16362 | ~n15566;
  assign n11136 = ~n11133 | ~n11132;
  assign n14784 = ~n15847 | ~n14809;
  assign n14640 = P2_REG3_REG_19__SCAN_IN ^ n10675;
  assign n10850 = ~n14203 | ~n14047;
  assign n14091 = ~n14086 | ~n14085;
  assign n14086 = ~n14078 | ~n14102;
  assign n13931 = ~n13926 | ~n13925;
  assign n13702 = ~n13740 | ~n10644;
  assign n13176 = ~n13175 | ~n13174;
  assign n13147 = ~n13146 | ~n13145;
  assign n14708 = ~n14707;
  assign n14120 = ~n14119 | ~n14118;
  assign n14018 = ~n14010;
  assign n14015 = ~n14014 | ~n14013;
  assign n13915 = ~n13933 | ~n13914;
  assign n13011 = ~n13008 | ~n13007;
  assign n12020 = ~n10723 & ~n10722;
  assign n11612 = ~P2_U3152 & ~n10878;
  assign n13947 = n10195 ^ P2_IR_REG_25__SCAN_IN;
  assign n13806 = n10216 ^ P2_IR_REG_24__SCAN_IN;
  assign n12681 = ~n10585 | ~n10584;
  assign n13874 = ~n10550 ^ P2_IR_REG_15__SCAN_IN;
  assign n13535 = n10548 ^ n10547;
  assign n12919 = n10513 ^ P2_IR_REG_13__SCAN_IN;
  assign n12581 = ~n12311;
  assign n12306 = n10471 ^ P2_IR_REG_11__SCAN_IN;
  assign n11962 = ~n11944;
  assign n10133 = n17103 ^ n17102;
  assign n14186 = ~n14185 ^ n14184;
  assign n15508 = n15507 ^ n15506;
  assign n13486 = ~n13484 | ~n13483;
  assign n12731 = n9244 ^ n9243;
  assign n17146 = ~n17150 & ~n17121;
  assign n17150 = ~n17103 & ~n17102;
  assign n16629 = ~n13474;
  assign n15085 = ~P1_REG3_REG_21__SCAN_IN ^ n9923;
  assign n15084 = ~n15083 ^ n15082;
  assign n15082 = ~n15081 ^ n15080;
  assign n15688 = n15687 ^ n15686;
  assign n14526 = n14525 ^ n14524;
  assign n14543 = n14542 ^ n14541;
  assign n14541 = ~n14540 | ~n14539;
  assign n15577 = ~n15576 ^ n15575;
  assign n14947 = ~P1_REG3_REG_20__SCAN_IN ^ n9884;
  assign n14946 = ~n15077 ^ n15076;
  assign n15582 = ~n15159;
  assign n15229 = ~n15228 ^ n15227;
  assign n14795 = ~P1_REG3_REG_18__SCAN_IN ^ n9844;
  assign n14794 = ~n14793 ^ n14792;
  assign n14804 = ~n14803 | ~n14802;
  assign n16777 = ~n16781;
  assign n15811 = n15810 ^ n15809;
  assign n14136 = ~n9705 | ~n9740;
  assign n10866 = ~n10865 ^ n10864;
  assign n10864 = ~n10863 ^ n10862;
  assign n9850 = ~n14852 | ~n9038;
  assign n9615 = n9614 & n9613;
  assign n9323 = n9322 & n9321;
  assign n9346 = n9345 & n9344;
  assign n9347 = ~n9342 & ~n9341;
  assign n12495 = ~n12825;
  assign n9218 = ~n9214 & ~n9213;
  assign n9142 = ~n12043 & ~n9141;
  assign n9076 = ~n9070 & ~n9069;
  assign n14340 = ~n14339 | ~n14338;
  assign n14625 = ~n14624 | ~n14623;
  assign n14623 = ~n14622 | ~n14830;
  assign n15359 = n16836 ^ n15217;
  assign n15350 = ~n17063 ^ n15760;
  assign n14975 = ~n15218 | ~n14974;
  assign n14936 = n17014 ^ n14977;
  assign n14920 = ~n14930 | ~n15762;
  assign n14758 = ~n17012 ^ n14923;
  assign n14743 = ~n14753 | ~n15762;
  assign n14927 = ~n15758;
  assign n13971 = ~n13970 | ~n13969;
  assign n13834 = ~n13833 | ~n13832;
  assign n15218 = ~n15745;
  assign n10763 = ~n12180 | ~n10762;
  assign n15805 = ~n15799 | ~n15798;
  assign n14278 = ~n14277 | ~n14276;
  assign n14375 = ~n14374 | ~n14373;
  assign n14299 = ~n14298 | ~n14297;
  assign n14395 = ~n14394 | ~n14393;
  assign n13247 = ~n13244 | ~n13243;
  assign n13169 = ~n13166 | ~n13165;
  assign n13383 = ~n13380 | ~n13379;
  assign n12745 = ~n12742 | ~n12741;
  assign n11074 = n11073 ^ SI_31_;
  assign n11060 = ~n15254;
  assign n14409 = ~P2_DATAO_REG_28__SCAN_IN;
  assign n14385 = ~n11034 ^ n11033;
  assign n13938 = ~n9084 ^ P1_IR_REG_25__SCAN_IN;
  assign n13155 = n9893 ^ n9892;
  assign n14828 = ~n9807 ^ P1_IR_REG_18__SCAN_IN;
  assign n9807 = ~n9806 | ~P1_IR_REG_31__SCAN_IN;
  assign n13774 = ~n14328;
  assign n13458 = n9646 ^ P1_IR_REG_14__SCAN_IN;
  assign n12983 = n9644 ^ P1_IR_REG_13__SCAN_IN;
  assign n12477 = n9574 ^ n9686;
  assign n9574 = ~n9684 | ~P1_IR_REG_31__SCAN_IN;
  assign n12105 = n9534 ^ P1_IR_REG_11__SCAN_IN;
  assign n11974 = n9482 ^ n9481;
  assign n9480 = ~n9479 | ~n9478;
  assign n11614 = n9375 ^ P1_IR_REG_7__SCAN_IN;
  assign n11469 = ~n9335 ^ P1_IR_REG_5__SCAN_IN;
  assign n11480 = n9282 ^ n9281;
  assign n11486 = ~n9161 ^ SI_1_;
  assign n9161 = ~n9186 | ~n9184;
  assign n11361 = ~n10815 | ~n10814;
  assign n10820 = ~n11379 | ~n11378;
  assign n11345 = ~n11344;
  assign n11032 = ~n11009 | ~n11008;
  assign n13656 = ~n13653 & ~n13652;
  assign n13889 = ~n13887 & ~n13886;
  assign n14050 = ~n14046 | ~n14045;
  assign n14007 = ~n14004 | ~n14003;
  assign n13735 = ~n13734 | ~n15720;
  assign n13635 = ~n13634 | ~n13633;
  assign n13269 = ~n13268 | ~n13267;
  assign n13681 = ~n16514 | ~n13680;
  assign n13750 = ~n16514 | ~n13749;
  assign n13498 = ~n16514 | ~n13500;
  assign n13678 = ~n16510 | ~n13680;
  assign n13747 = ~n16510 | ~n13749;
  assign n13501 = ~n16510 | ~n13500;
  assign n14862 = ~n14861 & ~n14860;
  assign n13862 = n13861 & n13860;
  assign n14681 = ~n14680 | ~n14679;
  assign n14664 = ~n14663 | ~n14662;
  assign n14500 = ~n14499 | ~n14498;
  assign n14319 = ~n14318 | ~n14927;
  assign n14316 = ~n14315 | ~n14314;
  assign n14241 = ~n14224 & ~n14223;
  assign n13608 = ~n13607 | ~n13606;
  assign n13668 = ~n15804 | ~n13667;
  assign n13800 = ~n15804 | ~n13802;
  assign n13665 = ~n15800 | ~n13667;
  assign n13803 = ~n15800 | ~n13802;
  assign n13757 = ~n13752 | ~n14582;
  assign n9170 = n11846 & n11845;
  assign n10888 = ~n14995 & ~n16472;
  assign n9041 = n9072 | n14583;
  assign n16391 = ~n16471 | ~n16080;
  assign n16461 = ~n16391;
  assign n9042 = n9558 & n13566;
  assign n16071 = ~n10645;
  assign n9043 = n9075 & n9074;
  assign n16082 = ~n16080;
  assign n16147 = ~n16146;
  assign n16212 = ~n16198;
  assign n15889 = ~n15887;
  assign n16306 = ~n16305;
  assign n16375 = ~n16372;
  assign n16390 = ~n16402 | ~n16398;
  assign n16822 = ~n16821;
  assign n15954 = ~n15953;
  assign n10931 = ~n10928;
  assign n11926 = ~P2_REG1_REG_7__SCAN_IN;
  assign n10892 = ~n10891;
  assign n10397 = ~P2_IR_REG_7__SCAN_IN;
  assign n11093 = ~n16316;
  assign n11692 = ~P1_REG2_REG_8__SCAN_IN;
  assign n9443 = ~P2_DATAO_REG_9__SCAN_IN;
  assign n16660 = ~n14144;
  assign n16616 = ~n16609;
  assign n10503 = ~n14164;
  assign n11175 = ~n11174;
  assign n14104 = ~n16266;
  assign n9394 = ~n9393;
  assign n9912 = ~n9910 | ~n9909;
  assign n15751 = ~n15748 & ~n17110;
  assign n14151 = ~n16678;
  assign n9406 = ~n9405;
  assign n9254 = ~P1_IR_REG_4__SCAN_IN;
  assign n11243 = ~n11242 | ~n11241;
  assign n10248 = ~n10519;
  assign n16199 = ~n16176;
  assign n16701 = ~n14527;
  assign n13371 = ~n16595;
  assign n9827 = ~n9826;
  assign n9701 = ~n9704;
  assign n9779 = ~P1_REG0_REG_17__SCAN_IN;
  assign n9488 = ~P1_REG0_REG_10__SCAN_IN;
  assign n11494 = ~n14837;
  assign n15646 = ~n15644 | ~n15643;
  assign n14984 = ~n15171;
  assign n14924 = ~n16739;
  assign n9800 = ~n9797 | ~n9796;
  assign n9564 = ~n9561 | ~n9560;
  assign n11632 = ~n10586;
  assign n12418 = ~n12414;
  assign n10367 = ~n10385;
  assign n15103 = ~n15099;
  assign n10240 = ~n10237 & ~P2_IR_REG_28__SCAN_IN;
  assign n11562 = ~n11469;
  assign n12986 = ~n13458;
  assign n15205 = ~n15759;
  assign n9065 = ~n9105 | ~n9063;
  assign n9761 = ~n9727 | ~n9726;
  assign n9595 = ~n9564 | ~n9563;
  assign n10221 = ~n10725;
  assign n14096 = ~P1_DATAO_REG_26__SCAN_IN;
  assign n11475 = ~n11935;
  assign n13598 = ~n13818;
  assign n16161 = ~n13317;
  assign n12671 = ~n9218 | ~n9217;
  assign P2_U3966 = ~n13390;
  assign n9189 = ~n9044 | ~n9164;
  assign n9045 = ~P1_IR_REG_6__SCAN_IN & ~P1_IR_REG_7__SCAN_IN;
  assign n9224 = ~P1_IR_REG_3__SCAN_IN;
  assign n9302 = ~n9254 | ~n9224;
  assign n9047 = ~n9046 & ~n9302;
  assign n9409 = ~n9304 | ~n9047;
  assign n9049 = ~P1_IR_REG_12__SCAN_IN & ~P1_IR_REG_11__SCAN_IN;
  assign n9048 = ~P1_IR_REG_13__SCAN_IN & ~P1_IR_REG_14__SCAN_IN;
  assign n9051 = ~P1_IR_REG_15__SCAN_IN & ~P1_IR_REG_16__SCAN_IN;
  assign n9052 = ~n9051 | ~n9050;
  assign n9054 = ~P1_IR_REG_22__SCAN_IN & ~P1_IR_REG_21__SCAN_IN;
  assign n9095 = ~P1_IR_REG_19__SCAN_IN & ~P1_IR_REG_10__SCAN_IN;
  assign n9058 = ~n9057 & ~n9056;
  assign n9059 = ~n9092 | ~n9058;
  assign n9107 = ~n10124 | ~n9062;
  assign n9105 = ~n9107 & ~P1_IR_REG_27__SCAN_IN;
  assign n11079 = ~n9065 & ~P1_IR_REG_29__SCAN_IN;
  assign n9064 = ~n11079 & ~n9733;
  assign n9066 = ~n9065 | ~P1_IR_REG_31__SCAN_IN;
  assign n9067 = ~P1_REG3_REG_0__SCAN_IN;
  assign n9070 = ~n9041 & ~n9067;
  assign n9068 = ~P1_REG0_REG_0__SCAN_IN;
  assign n9544 = ~n9072 & ~n9071;
  assign n11054 = ~n9072;
  assign n9073 = ~n11054 & ~n14583;
  assign n9656 = ~n9073;
  assign n10130 = ~n10124 | ~n10127;
  assign n13753 = ~n9083 | ~n9082;
  assign n9088 = ~n13938 & ~n13753;
  assign n9087 = ~n9086 | ~n9085;
  assign n11416 = ~n9088 | ~n10119;
  assign n9573 = ~n9409 & ~n9089;
  assign n9126 = ~n9090 | ~n9123;
  assign n9091 = ~n9126 | ~P1_IR_REG_31__SCAN_IN;
  assign n9102 = ~n9100 | ~P1_IR_REG_31__SCAN_IN;
  assign n9118 = ~n9102 | ~n9101;
  assign n9133 = ~n12534 | ~n17111;
  assign n9108 = ~n9107 | ~P1_IR_REG_31__SCAN_IN;
  assign n9114 = ~SI_0_;
  assign n9115 = ~n11089 & ~n9114;
  assign n11357 = n9115 ^ P2_DATAO_REG_0__SCAN_IN;
  assign n9117 = ~n10224 | ~n11357;
  assign n12282 = ~n9117 | ~n9116;
  assign n13503 = n9120 ^ n9119;
  assign n16962 = ~n13503 | ~n17072;
  assign n10791 = ~n9128 | ~n16962;
  assign n9271 = ~n10791 | ~n11416;
  assign n9131 = ~n12934 & ~n9271;
  assign n9129 = ~P1_REG1_REG_0__SCAN_IN;
  assign n9130 = ~n11416 & ~n9129;
  assign n11844 = ~n9133 | ~n9132;
  assign n9134 = ~n11844;
  assign n17107 = ~n10796 | ~n16962;
  assign n9140 = ~n9134 | ~n9752;
  assign n12281 = ~n13503 & ~n17037;
  assign n14237 = ~n15185 & ~n14836;
  assign n9136 = ~n12934 & ~n9934;
  assign n9135 = ~n11416 & ~n9044;
  assign n11843 = ~n9138 | ~n9137;
  assign n9139 = ~n11843 | ~n11844;
  assign n9178 = ~n9140 | ~n9139;
  assign n9141 = ~P1_REG0_REG_1__SCAN_IN;
  assign n9145 = ~n9038 | ~P1_REG3_REG_1__SCAN_IN;
  assign n9146 = n9145 & n9144;
  assign n12629 = ~n9147 | ~n9146;
  assign n9148 = ~P1_DATAO_REG_0__SCAN_IN;
  assign n9149 = ~n9148 & ~n11487;
  assign n9150 = P2_DATAO_REG_1__SCAN_IN & P2_DATAO_REG_0__SCAN_IN;
  assign n9151 = ~n9034 | ~n9150;
  assign n9155 = ~P2_DATAO_REG_0__SCAN_IN | ~SI_0_;
  assign n9156 = ~n9155 | ~n9154;
  assign n9160 = ~n10016 & ~n9156;
  assign n9157 = ~P1_DATAO_REG_0__SCAN_IN | ~SI_0_;
  assign n9158 = ~n9157 | ~n11487;
  assign n9159 = ~n9034 & ~n9158;
  assign n9184 = ~n9160 & ~n9159;
  assign n9162 = ~n11486;
  assign n9166 = ~n9163 | ~P1_IR_REG_1__SCAN_IN;
  assign n9165 = ~n9164 | ~P1_IR_REG_31__SCAN_IN;
  assign n9167 = ~n9166 | ~n9165;
  assign n11424 = ~n9167 | ~n9189;
  assign n9168 = ~n10224 & ~n11424;
  assign n9171 = ~n9601 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n12542 = ~n9172 | ~n9171;
  assign n17109 = ~n9271;
  assign n9173 = ~n12542 | ~n17109;
  assign n9175 = ~n9174 | ~n9173;
  assign n12550 = ~n12629;
  assign n9935 = ~n17104;
  assign n9177 = ~n12550 & ~n9935;
  assign n9176 = ~n12522 & ~n9934;
  assign n9182 = ~n12537 | ~n12539;
  assign n9181 = ~n9178;
  assign n12538 = ~n9181 | ~n9180;
  assign n10746 = ~n9182 | ~n12538;
  assign n9229 = ~n9186 | ~n9185;
  assign n9187 = ~n9034 | ~P2_DATAO_REG_2__SCAN_IN;
  assign n11545 = n9229 ^ n9228;
  assign n9192 = ~n15212 | ~n11545;
  assign n9190 = ~n9189 | ~P1_IR_REG_31__SCAN_IN;
  assign n11859 = ~n9190 ^ P1_IR_REG_2__SCAN_IN;
  assign n9191 = ~n9170 | ~n11859;
  assign n9195 = ~n9192 | ~n9191;
  assign n9839 = ~n9601;
  assign n9193 = ~P2_DATAO_REG_2__SCAN_IN;
  assign n12559 = ~n9195 & ~n9194;
  assign n16561 = ~n12559;
  assign n9204 = ~n16561 | ~n17109;
  assign n9196 = ~P1_REG0_REG_2__SCAN_IN;
  assign n9197 = ~n12043 & ~n9196;
  assign n9200 = ~n9544 | ~P1_REG2_REG_2__SCAN_IN;
  assign n9199 = ~n9038 | ~P1_REG3_REG_2__SCAN_IN;
  assign n9201 = n9200 & n9199;
  assign n12721 = ~n9202 | ~n9201;
  assign n9203 = ~n12721 | ~n17111;
  assign n16562 = ~n12721;
  assign n9207 = ~n16562 & ~n9935;
  assign n9206 = ~n12559 & ~n9934;
  assign n10745 = n9209 ^ n9208;
  assign n9211 = ~n10746 | ~n10745;
  assign n9210 = ~n9209 | ~n9208;
  assign n12730 = ~n9211 | ~n9210;
  assign n9212 = ~P1_REG0_REG_3__SCAN_IN;
  assign n9213 = ~n12043 & ~n9212;
  assign n9216 = ~n9544 | ~P1_REG2_REG_3__SCAN_IN;
  assign n9239 = ~n12671 | ~n17111;
  assign n9219 = ~P2_DATAO_REG_3__SCAN_IN;
  assign n9227 = ~n9839 & ~n9219;
  assign n9220 = ~n9304;
  assign n9221 = ~n9220 | ~P1_IR_REG_31__SCAN_IN;
  assign n9223 = ~n9221 | ~P1_IR_REG_3__SCAN_IN;
  assign n9222 = ~n9224 | ~P1_IR_REG_31__SCAN_IN;
  assign n9225 = ~n9223 | ~n9222;
  assign n9257 = ~n9304 | ~n9224;
  assign n11428 = ~n9225 | ~n9257;
  assign n9226 = ~n10224 & ~n11428;
  assign n9263 = ~n9232 | ~n9231;
  assign n11386 = ~n9263 ^ n9262;
  assign n9235 = ~n11386;
  assign n9236 = ~n15212 | ~n9235;
  assign n12720 = ~n9237 | ~n9236;
  assign n9238 = ~n12720 | ~n17109;
  assign n9244 = n9240 ^ n17107;
  assign n9242 = ~n16568 & ~n9935;
  assign n16567 = ~n12720;
  assign n9241 = ~n16567 & ~n9934;
  assign n9246 = ~n12730 | ~n12731;
  assign n9245 = ~n9244 | ~n9243;
  assign n12664 = ~n9246 | ~n9245;
  assign n9248 = ~n11671 | ~P1_REG0_REG_4__SCAN_IN;
  assign n9957 = ~n9544;
  assign n9247 = ~n9037 | ~P1_REG2_REG_4__SCAN_IN;
  assign n12791 = P1_REG3_REG_3__SCAN_IN ^ P1_REG3_REG_4__SCAN_IN;
  assign n9250 = ~n9038 | ~n12791;
  assign n9249 = ~n9612 | ~P1_REG1_REG_4__SCAN_IN;
  assign n9251 = ~n9250 | ~n9249;
  assign n12825 = ~n9252 & ~n9251;
  assign n9273 = ~n12825 & ~n9934;
  assign n11395 = ~P2_DATAO_REG_4__SCAN_IN;
  assign n9261 = ~n9839 & ~n11395;
  assign n9253 = ~n9257 | ~P1_IR_REG_31__SCAN_IN;
  assign n9256 = ~n9253 | ~P1_IR_REG_4__SCAN_IN;
  assign n9255 = ~n9254 | ~P1_IR_REG_31__SCAN_IN;
  assign n9259 = ~n9256 | ~n9255;
  assign n9334 = ~n9257 & ~P1_IR_REG_4__SCAN_IN;
  assign n9258 = ~n9334;
  assign n11452 = ~n9259 | ~n9258;
  assign n9260 = ~n10224 & ~n11452;
  assign n9270 = ~n9261 & ~n9260;
  assign n9282 = ~n9266 | ~n9265;
  assign n9269 = ~n11480 | ~n15212;
  assign n9272 = ~n12794 & ~n9271;
  assign n9277 = n9274 ^ n17107;
  assign n9276 = ~n12825 & ~n9935;
  assign n9275 = ~n12794 & ~n9934;
  assign n9278 = ~n9276 & ~n9275;
  assign n9279 = ~n9277;
  assign n9280 = ~n9279 & ~n9278;
  assign n12776 = ~n12666 & ~n9280;
  assign n9331 = ~n9285 | ~n9284;
  assign n9366 = ~n9290 | ~n9289;
  assign n9294 = ~P2_DATAO_REG_6__SCAN_IN;
  assign n9307 = ~n9839 & ~n9294;
  assign n9295 = ~n9334 | ~n9300;
  assign n9296 = ~n9295 | ~P1_IR_REG_31__SCAN_IN;
  assign n9298 = ~n9296 | ~P1_IR_REG_6__SCAN_IN;
  assign n9299 = ~P1_IR_REG_6__SCAN_IN;
  assign n9297 = ~n9299 | ~P1_IR_REG_31__SCAN_IN;
  assign n9305 = ~n9298 | ~n9297;
  assign n9301 = ~n9300 | ~n9299;
  assign n9303 = ~n9302 & ~n9301;
  assign n9374 = ~n9304 | ~n9303;
  assign n9306 = ~n10224 & ~n11532;
  assign n9308 = ~n9307 & ~n9306;
  assign n13114 = ~n9309 | ~n9308;
  assign n9326 = ~n13114 | ~n17109;
  assign n9310 = ~P1_REG1_REG_6__SCAN_IN;
  assign n9313 = ~n11675 & ~n9310;
  assign n9311 = ~P1_REG0_REG_6__SCAN_IN;
  assign n9312 = ~n12043 & ~n9311;
  assign n9324 = ~n9313 & ~n9312;
  assign n9322 = ~n9037 | ~P1_REG2_REG_6__SCAN_IN;
  assign n9317 = ~n9318;
  assign n9316 = ~P1_REG3_REG_6__SCAN_IN;
  assign n9319 = ~n9317 | ~n9316;
  assign n12767 = ~n9319 | ~n9418;
  assign n9320 = ~n12767;
  assign n9321 = ~n9038 | ~n9320;
  assign n16595 = ~n9324 | ~n9323;
  assign n9325 = ~n16595 | ~n17111;
  assign n9357 = n9327 ^ n17107;
  assign n9329 = ~n13114 | ~n17111;
  assign n9328 = ~n16595 | ~n17104;
  assign n9333 = ~P2_DATAO_REG_5__SCAN_IN;
  assign n9337 = ~n9839 & ~n9333;
  assign n9335 = ~n9334 & ~n9733;
  assign n9336 = ~n10224 & ~n11469;
  assign n9338 = ~n9337 & ~n9336;
  assign n12435 = ~n9339 | ~n9338;
  assign n9349 = ~n12435 | ~n17109;
  assign n9340 = ~P1_REG0_REG_5__SCAN_IN;
  assign n9341 = ~n12043 & ~n9340;
  assign n9343 = ~P1_REG3_REG_3__SCAN_IN | ~P1_REG3_REG_4__SCAN_IN;
  assign n12818 = ~n9343 ^ P1_REG3_REG_5__SCAN_IN;
  assign n9345 = ~n9038 | ~n12818;
  assign n9344 = ~n9612 | ~P1_REG1_REG_5__SCAN_IN;
  assign n12763 = ~n9347 | ~n9346;
  assign n9348 = ~n12763 | ~n17111;
  assign n12775 = n9350 ^ n17107;
  assign n9352 = ~n12763 | ~n17104;
  assign n9351 = ~n12435 | ~n17111;
  assign n9353 = ~n12775 | ~n12774;
  assign n9364 = ~n12776 & ~n9354;
  assign n9355 = ~n12775;
  assign n9359 = ~n9355 | ~n12819;
  assign n9358 = ~n9359 | ~n9356;
  assign n12751 = ~n9364 & ~n9363;
  assign n9398 = ~n9369 | ~n9368;
  assign n9373 = ~P2_DATAO_REG_7__SCAN_IN;
  assign n9377 = ~n9839 & ~n9373;
  assign n9375 = ~n9374 | ~P1_IR_REG_31__SCAN_IN;
  assign n9376 = ~n10224 & ~n11614;
  assign n9378 = ~n9377 & ~n9376;
  assign n13364 = ~n9379 | ~n9378;
  assign n9388 = ~n13364 | ~n17109;
  assign n9382 = n9037 & P1_REG2_REG_7__SCAN_IN;
  assign n9380 = ~P1_REG0_REG_7__SCAN_IN;
  assign n9381 = ~n12043 & ~n9380;
  assign n9386 = ~n9382 & ~n9381;
  assign n13420 = ~n9418 ^ P1_REG3_REG_7__SCAN_IN;
  assign n9384 = ~n9038 | ~n13420;
  assign n9383 = ~n9612 | ~P1_REG1_REG_7__SCAN_IN;
  assign n9385 = n9384 & n9383;
  assign n9387 = ~n13104 | ~n17111;
  assign n9392 = ~n9389 ^ n17107;
  assign n9391 = ~n13364 | ~n17111;
  assign n9390 = ~n13104 | ~n17104;
  assign n9396 = ~n12751 | ~n12749;
  assign n9395 = ~n9392;
  assign n9433 = ~n9396 | ~n12748;
  assign n9401 = ~n9398 | ~n9397;
  assign n9414 = ~n11739 | ~n15212;
  assign n9412 = ~n9839 & ~n9408;
  assign n9411 = ~n10224 & ~n11693;
  assign n9413 = ~n9412 & ~n9411;
  assign n13223 = ~n9414 | ~n9413;
  assign n9429 = ~n13223 | ~n17109;
  assign n9417 = n9612 & P1_REG1_REG_8__SCAN_IN;
  assign n9415 = ~P1_REG0_REG_8__SCAN_IN;
  assign n9416 = ~n12043 & ~n9415;
  assign n9427 = ~n9417 & ~n9416;
  assign n9425 = ~n9037 | ~P1_REG2_REG_8__SCAN_IN;
  assign n9420 = ~n9421;
  assign n9419 = ~P1_REG3_REG_8__SCAN_IN;
  assign n9422 = ~n9420 | ~n9419;
  assign n13130 = ~n9422 | ~n9491;
  assign n9423 = ~n13130;
  assign n9424 = ~n9038 | ~n9423;
  assign n9426 = n9425 & n9424;
  assign n9428 = ~n13228 | ~n17111;
  assign n9434 = n9430 ^ n17107;
  assign n12955 = ~n9433 | ~n9434;
  assign n9432 = ~n13223 | ~n17111;
  assign n9431 = ~n13228 | ~n17104;
  assign n12957 = ~n9432 | ~n9431;
  assign n9437 = ~n12955 | ~n12957;
  assign n9436 = ~n9433;
  assign n9435 = ~n9434;
  assign n12956 = ~n9436 | ~n9435;
  assign n13273 = ~n9437 | ~n12956;
  assign n9464 = ~n13273;
  assign n9472 = ~n9511 & ~n9513;
  assign n9448 = ~n9839 & ~n9443;
  assign n9444 = ~P1_IR_REG_8__SCAN_IN;
  assign n9447 = ~n10224 & ~n11721;
  assign n13280 = ~n9450 | ~n9449;
  assign n9460 = ~n13280 | ~n17109;
  assign n13285 = ~n9491 ^ P1_REG3_REG_9__SCAN_IN;
  assign n9451 = ~n13285;
  assign n9454 = ~n12041 & ~n9451;
  assign n9452 = ~P1_REG0_REG_9__SCAN_IN;
  assign n9453 = ~n12043 & ~n9452;
  assign n9458 = ~n9454 & ~n9453;
  assign n9456 = ~n9037 | ~P1_REG2_REG_9__SCAN_IN;
  assign n9455 = ~n9612 | ~P1_REG1_REG_9__SCAN_IN;
  assign n9457 = n9456 & n9455;
  assign n9459 = ~n13474 | ~n17111;
  assign n9463 = ~n13280 | ~n17111;
  assign n9462 = ~n13474 | ~n17104;
  assign n9470 = ~n9464 | ~n13274;
  assign n9506 = ~n9470 | ~n9469;
  assign n9477 = ~P2_DATAO_REG_10__SCAN_IN;
  assign n9484 = ~n9839 & ~n9477;
  assign n9478 = ~P1_IR_REG_9__SCAN_IN;
  assign n9483 = ~n10224 & ~n11759;
  assign n13611 = ~n9486 | ~n9485;
  assign n9502 = ~n13611 | ~n17109;
  assign n9487 = ~P1_REG1_REG_10__SCAN_IN;
  assign n9490 = ~n11675 & ~n9487;
  assign n9489 = ~n12043 & ~n9488;
  assign n9500 = ~n9490 & ~n9489;
  assign n9498 = ~n9037 | ~P1_REG2_REG_10__SCAN_IN;
  assign n9493 = ~n9494;
  assign n9492 = ~P1_REG3_REG_10__SCAN_IN;
  assign n9495 = ~n9493 | ~n9492;
  assign n13473 = ~n9495 | ~n9584;
  assign n9496 = ~n13473;
  assign n9497 = ~n9038 | ~n9496;
  assign n9499 = n9498 & n9497;
  assign n9501 = ~n13783 | ~n17111;
  assign n13484 = ~n9506 | ~n9507;
  assign n9505 = ~n13611 | ~n17111;
  assign n9504 = ~n13783 | ~n17104;
  assign n9510 = ~n13484 | ~n13485;
  assign n9509 = ~n9506;
  assign n13483 = ~n9509 | ~n9508;
  assign n13568 = ~n9510 | ~n13483;
  assign n9522 = ~n9511 | ~n9512;
  assign n9537 = ~n9839 & ~n9533;
  assign n9535 = ~n12105;
  assign n9536 = ~n10224 & ~n9535;
  assign n9540 = ~P1_REG1_REG_11__SCAN_IN;
  assign n9543 = ~n11675 & ~n9540;
  assign n9541 = ~P1_REG0_REG_11__SCAN_IN;
  assign n9542 = ~n12043 & ~n9541;
  assign n9548 = ~n9543 & ~n9542;
  assign n9546 = ~n9037 | ~P1_REG2_REG_11__SCAN_IN;
  assign n13842 = ~n9584 ^ P1_REG3_REG_11__SCAN_IN;
  assign n9545 = ~n9038 | ~n13842;
  assign n9547 = n9546 & n9545;
  assign n9549 = ~n13818 | ~n17111;
  assign n9552 = ~n13818 | ~n17104;
  assign n9558 = ~n13568 | ~n13565;
  assign n9577 = ~n9839 & ~n9571;
  assign n9686 = ~P1_IR_REG_12__SCAN_IN;
  assign n9575 = ~n12477;
  assign n9576 = ~n10224 & ~n9575;
  assign n13973 = ~n9579 | ~n9578;
  assign n9590 = ~n13973 | ~n17109;
  assign n9580 = ~P1_REG1_REG_12__SCAN_IN;
  assign n9583 = ~n11675 & ~n9580;
  assign n9581 = ~P1_REG0_REG_12__SCAN_IN;
  assign n9582 = ~n12043 & ~n9581;
  assign n9586 = ~n9037 | ~P1_REG2_REG_12__SCAN_IN;
  assign n13811 = n9652 ^ P1_REG3_REG_12__SCAN_IN;
  assign n9585 = ~n9038 | ~n13811;
  assign n9587 = n9586 & n9585;
  assign n9589 = ~n13855 | ~n17111;
  assign n9593 = ~n13973 | ~n17111;
  assign n9592 = ~n13855 | ~n17104;
  assign n9598 = ~n9595 | ~n9594;
  assign n16668 = ~n9606 | ~n9605;
  assign n9607 = ~n9652 | ~P1_REG3_REG_12__SCAN_IN;
  assign n13979 = ~n9607 ^ P1_REG3_REG_13__SCAN_IN;
  assign n9608 = ~n13979;
  assign n9611 = ~n12041 & ~n9608;
  assign n9609 = ~P1_REG0_REG_13__SCAN_IN;
  assign n9610 = ~n12043 & ~n9609;
  assign n9613 = ~n9612 | ~P1_REG1_REG_13__SCAN_IN;
  assign n9617 = ~n16666 | ~n17111;
  assign n9621 = ~n16668 | ~n17111;
  assign n9620 = ~n16666 | ~n17104;
  assign n13852 = ~n13812 | ~n9629;
  assign n9674 = ~n9640 | ~n9639;
  assign n9648 = ~n9839 & ~n9643;
  assign n9645 = ~n9644 & ~P1_IR_REG_13__SCAN_IN;
  assign n9647 = ~n12986 & ~n10224;
  assign n16657 = ~n9650 | ~n9649;
  assign n14218 = n9704 ^ P1_REG3_REG_14__SCAN_IN;
  assign n9655 = ~n12041 & ~n14218;
  assign n9653 = ~P1_REG0_REG_14__SCAN_IN;
  assign n9654 = ~n12043 & ~n9653;
  assign n9658 = ~n9037 | ~P1_REG2_REG_14__SCAN_IN;
  assign n9657 = ~n12046 | ~P1_REG1_REG_14__SCAN_IN;
  assign n9659 = n9658 & n9657;
  assign n14182 = ~n9666 | ~n9667;
  assign n9665 = ~n16657 | ~n17111;
  assign n9664 = ~n16678 | ~n17104;
  assign n9670 = ~n14182 | ~n14184;
  assign n9669 = ~n9666;
  assign n14183 = ~n9669 | ~n9668;
  assign n10865 = ~n9670 | ~n14183;
  assign n9716 = ~n10865;
  assign n9675 = ~n9673 | ~n9672;
  assign n9679 = ~n9677 & ~n9676;
  assign n9723 = ~n9681 & ~n9725;
  assign n9698 = ~n9839 & ~n9683;
  assign n9685 = ~P1_IR_REG_13__SCAN_IN;
  assign n9687 = ~n9686 | ~n9685;
  assign n9688 = ~n9687 & ~P1_IR_REG_14__SCAN_IN;
  assign n9690 = ~n9694 | ~P1_IR_REG_31__SCAN_IN;
  assign n9693 = ~n9690 | ~P1_IR_REG_15__SCAN_IN;
  assign n9691 = ~P1_IR_REG_15__SCAN_IN;
  assign n9692 = ~n9691 | ~P1_IR_REG_31__SCAN_IN;
  assign n9696 = ~n9693 | ~n9692;
  assign n9695 = ~n9772;
  assign n9697 = ~n10224 & ~n13461;
  assign n14296 = ~n9700 | ~n9699;
  assign n9702 = ~n9701 | ~P1_REG3_REG_14__SCAN_IN;
  assign n10867 = ~P1_REG3_REG_15__SCAN_IN;
  assign n9705 = ~n9702 | ~n10867;
  assign n9740 = ~n9741;
  assign n9708 = ~n12041 & ~n14136;
  assign n9706 = ~P1_REG0_REG_15__SCAN_IN;
  assign n9707 = ~n12043 & ~n9706;
  assign n9710 = ~n9037 | ~P1_REG2_REG_15__SCAN_IN;
  assign n9709 = ~n12046 | ~P1_REG1_REG_15__SCAN_IN;
  assign n9711 = n9710 & n9709;
  assign n9713 = ~n14527 | ~n17111;
  assign n9719 = ~n9716 | ~n10863;
  assign n9717 = ~n14527 | ~n17104;
  assign n9722 = ~n9719 | ~n10862;
  assign n9721 = ~n10865 | ~n9720;
  assign n9732 = ~P2_DATAO_REG_16__SCAN_IN;
  assign n9736 = ~n9839 & ~n9732;
  assign n9734 = ~n9772 & ~n9733;
  assign n9735 = ~n13774 & ~n10224;
  assign n16692 = ~n9738 | ~n9737;
  assign n9739 = ~P1_REG3_REG_16__SCAN_IN;
  assign n9742 = ~n9740 | ~n9739;
  assign n14536 = ~n9742 | ~n9812;
  assign n9745 = ~n12041 & ~n14536;
  assign n9743 = ~P1_REG0_REG_16__SCAN_IN;
  assign n9744 = ~n12043 & ~n9743;
  assign n9747 = ~n9037 | ~P1_REG2_REG_16__SCAN_IN;
  assign n9746 = ~n12046 | ~P1_REG1_REG_16__SCAN_IN;
  assign n9748 = n9747 & n9746;
  assign n9754 = ~n16693 | ~n17104;
  assign n9760 = ~n14525 & ~n14522;
  assign n14542 = ~n9760 & ~n14523;
  assign n9766 = ~n9763 | ~n9762;
  assign n9765 = ~n9764 | ~SI_16_;
  assign n9769 = ~n9797;
  assign n9777 = ~n9770 | ~n15212;
  assign n9771 = ~P1_IR_REG_16__SCAN_IN;
  assign n9804 = ~P1_IR_REG_17__SCAN_IN;
  assign n16716 = ~n9777 | ~n9776;
  assign n9778 = ~P1_REG2_REG_17__SCAN_IN;
  assign n9781 = ~n9957 & ~n9778;
  assign n9780 = ~n12043 & ~n9779;
  assign n9785 = ~n9781 & ~n9780;
  assign n14544 = ~n9812 ^ P1_REG3_REG_17__SCAN_IN;
  assign n9783 = ~n9038 | ~n14544;
  assign n9782 = ~n12046 | ~P1_REG1_REG_17__SCAN_IN;
  assign n9784 = n9783 & n9782;
  assign n9789 = ~n16717 | ~n17104;
  assign n9795 = ~n14542 | ~n14540;
  assign n9825 = ~n9795 | ~n14539;
  assign n9799 = ~n9798 | ~SI_17_;
  assign n9811 = ~n12842 | ~n15212;
  assign n9806 = ~n9805 | ~n9804;
  assign n9809 = ~n14828 | ~n9170;
  assign n14797 = ~n9811 | ~n9810;
  assign n9819 = n14795 | n12041;
  assign n9814 = ~n11671 | ~P1_REG0_REG_18__SCAN_IN;
  assign n9813 = ~n9037 | ~P1_REG2_REG_18__SCAN_IN;
  assign n9815 = ~P1_REG1_REG_18__SCAN_IN;
  assign n9816 = ~n11675 & ~n9815;
  assign n14790 = ~n9825 | ~n9826;
  assign n9823 = ~n14605 | ~n17104;
  assign n9829 = ~n14790 | ~n14792;
  assign n9828 = ~n9825;
  assign n14791 = ~n9828 | ~n9827;
  assign n14848 = ~n9829 | ~n14791;
  assign n9833 = ~n9832 | ~SI_18_;
  assign n9862 = ~n9834 | ~n9833;
  assign n9843 = ~n13065 | ~n15212;
  assign n9838 = ~P2_DATAO_REG_19__SCAN_IN;
  assign n9841 = ~n9839 & ~n9838;
  assign n9840 = ~n10224 & ~n17072;
  assign n16548 = ~n9843 | ~n9842;
  assign n9846 = ~n11671 | ~P1_REG0_REG_19__SCAN_IN;
  assign n9845 = ~n12046 | ~P1_REG1_REG_19__SCAN_IN;
  assign n14659 = ~P1_REG2_REG_19__SCAN_IN;
  assign n9847 = ~n9957 & ~n14659;
  assign n9854 = ~n16534 | ~n17104;
  assign n9860 = ~n14848 | ~n14845;
  assign n15077 = ~n9860 | ~n14846;
  assign n9869 = ~n13155 | ~n15212;
  assign n9877 = n14947 | n12041;
  assign n9872 = ~n11671 | ~P1_REG0_REG_20__SCAN_IN;
  assign n9871 = ~n9037 | ~P1_REG2_REG_20__SCAN_IN;
  assign n9873 = ~P1_REG1_REG_20__SCAN_IN;
  assign n9874 = ~n11675 & ~n9873;
  assign n9891 = n15085 | n12041;
  assign n9886 = ~n11671 | ~P1_REG0_REG_21__SCAN_IN;
  assign n9885 = ~n9037 | ~P1_REG2_REG_21__SCAN_IN;
  assign n9887 = ~P1_REG1_REG_21__SCAN_IN;
  assign n9888 = ~n11675 & ~n9887;
  assign n9895 = ~n9894 | ~SI_20_;
  assign n9914 = ~n9896 | ~n9895;
  assign n9900 = ~n13334 | ~n15212;
  assign n9917 = ~n9914 | ~n9913;
  assign n9916 = ~n9915 | ~SI_21_;
  assign n9944 = ~n9917 | ~n9916;
  assign n9922 = ~n9920 | ~n15212;
  assign n9930 = ~n15230 | ~n9038;
  assign n9925 = ~n11671 | ~P1_REG0_REG_22__SCAN_IN;
  assign n9924 = ~n12046 | ~P1_REG1_REG_22__SCAN_IN;
  assign n9926 = ~P1_REG2_REG_22__SCAN_IN;
  assign n9927 = ~n9957 & ~n9926;
  assign n15225 = ~n9938 & ~n9939;
  assign n9936 = ~n14906 & ~n9935;
  assign n9942 = ~n15225 & ~n15227;
  assign n9941 = ~n9938;
  assign n15226 = ~n9941 & ~n9940;
  assign n9966 = ~n9968;
  assign n9946 = ~n9945 | ~SI_22_;
  assign n9981 = ~n9947 | ~n9946;
  assign n9982 = ~n9949 | ~n9948;
  assign n9953 = ~n9951 | ~n15212;
  assign n9961 = ~n15510 | ~n9038;
  assign n9956 = ~n11671 | ~P1_REG0_REG_23__SCAN_IN;
  assign n9955 = ~n12046 | ~P1_REG1_REG_23__SCAN_IN;
  assign n14974 = ~P1_REG2_REG_23__SCAN_IN;
  assign n9958 = ~n9957 & ~n14974;
  assign n15159 = ~n9961 | ~n9960;
  assign n15504 = ~n9966 & ~n9965;
  assign n9969 = ~n15159 | ~n17104;
  assign n9971 = ~n15505 & ~n15506;
  assign n15576 = ~n15504 & ~n9971;
  assign n9979 = ~n15585 | ~n9038;
  assign n9974 = ~n11671 | ~P1_REG0_REG_24__SCAN_IN;
  assign n9973 = ~n9037 | ~P1_REG2_REG_24__SCAN_IN;
  assign n9975 = ~P1_REG1_REG_24__SCAN_IN;
  assign n9976 = ~n11675 & ~n9975;
  assign n15697 = ~n9979 | ~n9978;
  assign n9983 = ~n9982 | ~SI_23_;
  assign n10012 = ~n9986 | ~n9985;
  assign n9988 = ~n13752 | ~n15212;
  assign n10001 = ~n15576 & ~n15575;
  assign n15687 = ~n10001 & ~n10000;
  assign n10009 = ~n15691 | ~n9038;
  assign n10004 = ~n9037 | ~P1_REG2_REG_25__SCAN_IN;
  assign n10003 = ~n12046 | ~P1_REG1_REG_25__SCAN_IN;
  assign n10005 = ~P1_REG0_REG_25__SCAN_IN;
  assign n10006 = ~n12043 & ~n10005;
  assign n10013 = ~n10012 | ~SI_24_;
  assign n10043 = ~n10014 | ~n10013;
  assign n10020 = ~n10018 & ~n10017;
  assign n10044 = ~n10020 | ~n10019;
  assign n10025 = ~n10023 | ~n15212;
  assign n15810 = ~n10033 & ~n15684;
  assign n10041 = ~n15812 | ~n9038;
  assign n10036 = ~n9037 | ~P1_REG2_REG_26__SCAN_IN;
  assign n10035 = ~n12046 | ~P1_REG1_REG_26__SCAN_IN;
  assign n10037 = ~P1_REG0_REG_26__SCAN_IN;
  assign n10038 = ~n12043 & ~n10037;
  assign n10046 = ~n10043 & ~n10042;
  assign n10063 = ~n10048 | ~n10047;
  assign n10051 = ~n14037 | ~n15212;
  assign n10060 = ~n15810 | ~n15809;
  assign n17103 = n10060 & n10059;
  assign n11035 = ~n10067 | ~n10066;
  assign n10069 = ~n14197 | ~n15212;
  assign n10068 = ~n15214 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n10071 = ~P1_REG0_REG_27__SCAN_IN;
  assign n10072 = ~n12043 & ~n10071;
  assign n10075 = ~n9037 | ~P1_REG2_REG_27__SCAN_IN;
  assign n10074 = ~n12046 | ~P1_REG1_REG_27__SCAN_IN;
  assign n10076 = n10075 & n10074;
  assign n10084 = ~P1_D_REG_12__SCAN_IN & ~P1_D_REG_13__SCAN_IN;
  assign n10083 = ~P1_D_REG_10__SCAN_IN & ~P1_D_REG_11__SCAN_IN;
  assign n10088 = ~n10084 | ~n10083;
  assign n10086 = ~P1_D_REG_8__SCAN_IN & ~P1_D_REG_9__SCAN_IN;
  assign n10085 = ~P1_D_REG_6__SCAN_IN & ~P1_D_REG_7__SCAN_IN;
  assign n10087 = ~n10086 | ~n10085;
  assign n10110 = n10088 | n10087;
  assign n10090 = ~P1_D_REG_4__SCAN_IN & ~P1_D_REG_5__SCAN_IN;
  assign n10089 = ~P1_D_REG_2__SCAN_IN & ~P1_D_REG_3__SCAN_IN;
  assign n10091 = ~n10090 | ~n10089;
  assign n10108 = ~n10091 & ~P1_D_REG_29__SCAN_IN;
  assign n10093 = ~P1_D_REG_28__SCAN_IN & ~P1_D_REG_31__SCAN_IN;
  assign n10092 = ~P1_D_REG_26__SCAN_IN & ~P1_D_REG_27__SCAN_IN;
  assign n10097 = ~n10093 | ~n10092;
  assign n10095 = ~P1_D_REG_15__SCAN_IN & ~P1_D_REG_17__SCAN_IN;
  assign n10094 = ~P1_D_REG_16__SCAN_IN & ~P1_D_REG_14__SCAN_IN;
  assign n10096 = ~n10095 | ~n10094;
  assign n10105 = ~n10097 & ~n10096;
  assign n10099 = ~P1_D_REG_24__SCAN_IN & ~P1_D_REG_25__SCAN_IN;
  assign n10098 = ~P1_D_REG_22__SCAN_IN & ~P1_D_REG_23__SCAN_IN;
  assign n10103 = ~n10099 | ~n10098;
  assign n10101 = ~P1_D_REG_20__SCAN_IN & ~P1_D_REG_21__SCAN_IN;
  assign n10100 = ~P1_D_REG_18__SCAN_IN & ~P1_D_REG_19__SCAN_IN;
  assign n10102 = ~n10101 | ~n10100;
  assign n10104 = ~n10103 & ~n10102;
  assign n10106 = ~n10105 | ~n10104;
  assign n10107 = ~n10106 & ~P1_D_REG_30__SCAN_IN;
  assign n10109 = ~n10108 | ~n10107;
  assign n10116 = ~n10110 & ~n10109;
  assign n10112 = ~P1_B_REG_SCAN_IN;
  assign n10117 = ~n10115 | ~n10119;
  assign n12154 = ~n10116 & ~n10117;
  assign n10118 = ~P1_D_REG_1__SCAN_IN;
  assign n12158 = ~n10120 | ~n11365;
  assign n10121 = ~P1_D_REG_0__SCAN_IN;
  assign n10125 = ~n10124;
  assign n17086 = ~n10131 | ~n10130;
  assign n10174 = ~n17092 & ~P1_U3084;
  assign n17089 = ~n17073 | ~n17072;
  assign n15422 = ~n12281 | ~n17089;
  assign n10222 = ~n13503 | ~n17037;
  assign n10132 = n10147 & n10137;
  assign n10173 = ~n10133 | ~n10132;
  assign n10134 = ~n15594 & ~n17089;
  assign n17136 = ~n10147 | ~n10134;
  assign n10171 = ~n16816 & ~n17136;
  assign n10135 = ~n12281;
  assign n12156 = ~n15619 & ~n17037;
  assign n10140 = n10749 & n10137;
  assign n10138 = ~n10175 & ~n17092;
  assign n10139 = ~n10138 | ~n10760;
  assign n10146 = ~n10751 & ~P1_U3084;
  assign n10144 = ~n10749;
  assign n10142 = ~n11369 & ~n10222;
  assign n13152 = ~n17073 & ~P1_U3084;
  assign n10143 = ~n10142 & ~n13152;
  assign n10145 = ~n10144 & ~n10143;
  assign n17130 = n10146 | n10145;
  assign n15086 = ~n17130;
  assign n10167 = ~n15086 & ~n15610;
  assign n10150 = ~n10147;
  assign n15636 = ~n10222 & ~n11423;
  assign n10148 = ~n17089;
  assign n10149 = ~n15636 | ~n10148;
  assign n17132 = ~n10150 & ~n10149;
  assign n10154 = ~P1_REG3_REG_28__SCAN_IN;
  assign n10151 = ~P1_REG3_REG_27__SCAN_IN;
  assign n10157 = ~P1_REG0_REG_28__SCAN_IN;
  assign n10158 = ~n12043 & ~n10157;
  assign n10161 = ~n9037 | ~P1_REG2_REG_28__SCAN_IN;
  assign n10160 = ~n12046 | ~P1_REG1_REG_28__SCAN_IN;
  assign n10162 = n10161 & n10160;
  assign n17112 = ~n10163 | ~n10162;
  assign n10165 = ~n17132 | ~n17112;
  assign n10164 = ~P1_U3084 | ~P1_REG3_REG_27__SCAN_IN;
  assign n10166 = ~n10165 | ~n10164;
  assign n10168 = ~n10167 & ~n10166;
  assign P1_U3212 = ~n10173 | ~n10172;
  assign n10177 = ~P2_IR_REG_14__SCAN_IN & ~P2_IR_REG_11__SCAN_IN;
  assign n10176 = ~P2_IR_REG_12__SCAN_IN & ~P2_IR_REG_10__SCAN_IN;
  assign n10178 = ~P2_IR_REG_15__SCAN_IN & ~P2_IR_REG_13__SCAN_IN;
  assign n10349 = ~P2_IR_REG_5__SCAN_IN;
  assign n10184 = n10180 | n10179;
  assign n10185 = ~n10184 & ~n10183;
  assign n10311 = ~n10289 & ~P2_IR_REG_2__SCAN_IN;
  assign n10326 = ~n10311 | ~n10312;
  assign n10350 = ~n10326 & ~P2_IR_REG_4__SCAN_IN;
  assign n10196 = ~n10185 | ~n10350;
  assign n10199 = ~P2_IR_REG_17__SCAN_IN & ~P2_IR_REG_16__SCAN_IN;
  assign n10194 = ~n10639 & ~n10193;
  assign n10195 = ~n10194 & ~n10608;
  assign n10232 = ~n10196;
  assign n10205 = ~n10204 & ~n10203;
  assign n10206 = ~n10209 | ~P2_IR_REG_31__SCAN_IN;
  assign n10229 = ~n10211 | ~n10210;
  assign n10716 = ~n10229 | ~n10212;
  assign n10213 = ~n10639 & ~P2_IR_REG_22__SCAN_IN;
  assign n10219 = ~n10215 | ~n10214;
  assign n10216 = ~n10219 | ~P2_IR_REG_31__SCAN_IN;
  assign n10725 = ~n10217 | ~n10721;
  assign n13709 = ~n10220 | ~n10219;
  assign n10228 = ~n10237 | ~P2_IR_REG_31__SCAN_IN;
  assign n14404 = n10228 ^ P2_IR_REG_28__SCAN_IN;
  assign n10230 = ~n10229 | ~P2_IR_REG_31__SCAN_IN;
  assign n10231 = ~P1_DATAO_REG_19__SCAN_IN;
  assign n10579 = ~n10232 | ~n10565;
  assign n10605 = ~n10579 & ~P2_IR_REG_17__SCAN_IN;
  assign n10611 = ~n10605 | ~n10606;
  assign n16472 = ~n10630 ^ P2_IR_REG_19__SCAN_IN;
  assign n10241 = ~n10240 & ~n10608;
  assign n10244 = n10241 ^ P2_IR_REG_29__SCAN_IN;
  assign n14576 = ~n10244;
  assign n10412 = ~n10245 & ~n14576;
  assign n10246 = P2_REG3_REG_3__SCAN_IN & P2_REG3_REG_5__SCAN_IN;
  assign n10255 = ~n9033 | ~P2_REG0_REG_0__SCAN_IN;
  assign n10259 = n10255 & n10254;
  assign n10257 = ~n11807 | ~P2_REG1_REG_0__SCAN_IN;
  assign n10258 = n10257 & n10256;
  assign n12383 = ~n10259 | ~n10258;
  assign n16081 = ~n12383;
  assign n10260 = ~n11089 | ~SI_0_;
  assign n10742 = n10260 ^ P1_DATAO_REG_0__SCAN_IN;
  assign n10263 = ~n10586 & ~n10742;
  assign n10262 = ~n11632 & ~n10261;
  assign n10645 = n10263 | n10262;
  assign n12345 = ~n16081 & ~n16071;
  assign n10280 = ~n12345;
  assign n10265 = ~n11803 | ~P2_REG0_REG_1__SCAN_IN;
  assign n10264 = ~n10412 | ~P2_REG3_REG_1__SCAN_IN;
  assign n10269 = ~n10265 | ~n10264;
  assign n10267 = ~n11807 | ~P2_REG1_REG_1__SCAN_IN;
  assign n10266 = ~n10476 | ~P2_REG2_REG_1__SCAN_IN;
  assign n10273 = ~n10270 | ~P2_IR_REG_1__SCAN_IN;
  assign n10272 = ~n10271 | ~P2_IR_REG_31__SCAN_IN;
  assign n10274 = ~n10273 | ~n10272;
  assign n11653 = ~n10274 | ~n10289;
  assign n10275 = ~n11632 & ~n11653;
  assign n10277 = ~n10310 | ~n11486;
  assign n12351 = ~n10278 | ~n10277;
  assign n10279 = ~n12388 | ~n12351;
  assign n10282 = ~n10280 | ~n10279;
  assign n16090 = ~n12351;
  assign n12596 = ~n10282 | ~n10281;
  assign n10284 = ~n11803 | ~P2_REG0_REG_2__SCAN_IN;
  assign n10283 = ~n10412 | ~P2_REG3_REG_2__SCAN_IN;
  assign n10286 = ~n11807 | ~P2_REG1_REG_2__SCAN_IN;
  assign n10285 = ~n10476 | ~P2_REG2_REG_2__SCAN_IN;
  assign n16073 = ~n10288 | ~n10287;
  assign n10290 = ~n10289 | ~P2_IR_REG_31__SCAN_IN;
  assign n10293 = ~n10290 | ~P2_IR_REG_2__SCAN_IN;
  assign n10291 = ~P2_IR_REG_2__SCAN_IN;
  assign n10292 = ~n10291 | ~P2_IR_REG_31__SCAN_IN;
  assign n10295 = ~n10293 | ~n10292;
  assign n10294 = ~n10311;
  assign n11655 = ~n10295 | ~n10294;
  assign n12236 = ~n11655;
  assign n10296 = ~n10586 | ~n12236;
  assign n10298 = ~P1_DATAO_REG_2__SCAN_IN;
  assign n13050 = ~n10300 & ~n10299;
  assign n16093 = ~n13050;
  assign n10301 = ~n16073 | ~n16093;
  assign n10302 = ~n12596 | ~n10301;
  assign n16104 = ~n16076 | ~n13050;
  assign n12888 = ~n10302 | ~n16104;
  assign n10305 = ~n10476 | ~P2_REG2_REG_3__SCAN_IN;
  assign n10303 = ~P2_REG3_REG_3__SCAN_IN;
  assign n10304 = ~n9035 | ~n10303;
  assign n10307 = ~n11807 | ~P2_REG1_REG_3__SCAN_IN;
  assign n10313 = ~n10311 & ~n10608;
  assign n11657 = n10313 ^ n10312;
  assign n10314 = ~n11632 & ~n11657;
  assign n10317 = ~n10315 & ~n10314;
  assign n10316 = ~n15258 | ~P1_DATAO_REG_3__SCAN_IN;
  assign n13144 = ~n10317 | ~n10316;
  assign n12889 = n16124 ^ n13144;
  assign n10319 = ~n12888 | ~n15971;
  assign n16125 = ~n13144;
  assign n10318 = ~n16124 | ~n16125;
  assign n12691 = ~n10319 | ~n10318;
  assign n10321 = ~n11807 | ~P2_REG1_REG_4__SCAN_IN;
  assign n10320 = ~n10476 | ~P2_REG2_REG_4__SCAN_IN;
  assign n10325 = ~n10321 | ~n10320;
  assign n10323 = ~n11803 | ~P2_REG0_REG_4__SCAN_IN;
  assign n12848 = P2_REG3_REG_4__SCAN_IN ^ P2_REG3_REG_3__SCAN_IN;
  assign n10322 = ~n9035 | ~n12848;
  assign n12890 = ~n10325 & ~n10324;
  assign n11481 = ~P1_DATAO_REG_4__SCAN_IN;
  assign n10334 = ~n15371 & ~n11481;
  assign n10327 = ~n10326 | ~P2_IR_REG_31__SCAN_IN;
  assign n10330 = ~n10327 | ~P2_IR_REG_4__SCAN_IN;
  assign n10328 = ~P2_IR_REG_4__SCAN_IN;
  assign n10329 = ~n10328 | ~P2_IR_REG_31__SCAN_IN;
  assign n10332 = ~n10330 | ~n10329;
  assign n10331 = ~n10350;
  assign n11659 = ~n10332 | ~n10331;
  assign n10333 = ~n11632 & ~n11659;
  assign n10336 = ~n10334 & ~n10333;
  assign n10335 = ~n10310 | ~n11480;
  assign n12695 = n12890 ^ n12687;
  assign n10338 = ~n12691 | ~n15976;
  assign n10337 = ~n12890 | ~n16115;
  assign n12865 = ~n10338 | ~n10337;
  assign n10341 = ~n11803 | ~P2_REG0_REG_5__SCAN_IN;
  assign n10339 = ~P2_REG3_REG_4__SCAN_IN | ~P2_REG3_REG_3__SCAN_IN;
  assign n13075 = ~n10339 ^ P2_REG3_REG_5__SCAN_IN;
  assign n10340 = ~n9035 | ~n13075;
  assign n10343 = ~n11807 | ~P2_REG1_REG_5__SCAN_IN;
  assign n10342 = ~n10476 | ~P2_REG2_REG_5__SCAN_IN;
  assign n13014 = ~n10345 | ~n10344;
  assign n10356 = ~n11474 & ~n9036;
  assign n10354 = ~n15258 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n10346 = ~n10350 & ~n10608;
  assign n10348 = ~n10346 & ~n10349;
  assign n10347 = ~n10608 & ~P2_IR_REG_5__SCAN_IN;
  assign n10352 = ~n10348 & ~n10347;
  assign n10399 = ~n10350 | ~n10349;
  assign n10351 = ~n10399;
  assign n10353 = ~n10586 | ~n11935;
  assign n13078 = ~n10356 & ~n10355;
  assign n16111 = ~n12994 & ~n12876;
  assign n16136 = ~n16111;
  assign n15969 = ~n16136 | ~n16150;
  assign n12866 = ~n15969;
  assign n10358 = ~n12865 & ~n12866;
  assign n10357 = ~n12994 & ~n13078;
  assign n10363 = ~n11537 & ~n9036;
  assign n10361 = ~n15258 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n10359 = ~n10399 | ~P2_IR_REG_31__SCAN_IN;
  assign n10360 = ~n10586 | ~n12273;
  assign n13032 = ~n10363 & ~n10362;
  assign n10370 = ~n9033 | ~P2_REG0_REG_6__SCAN_IN;
  assign n10366 = ~n10365 | ~n10364;
  assign n13033 = ~n10367 | ~n10366;
  assign n10368 = ~n13033;
  assign n10369 = ~n9035 | ~n10368;
  assign n10372 = ~n11807 | ~P2_REG1_REG_6__SCAN_IN;
  assign n10371 = ~n11804 | ~P2_REG2_REG_6__SCAN_IN;
  assign n13251 = ~n10374 | ~n10373;
  assign n10378 = ~n12993 & ~n15977;
  assign n10377 = ~n10376;
  assign n10384 = ~n11626 & ~n9036;
  assign n10379 = ~n10399 & ~P2_IR_REG_6__SCAN_IN;
  assign n10380 = ~n10379 & ~n10608;
  assign n10381 = ~n10586 | ~n12070;
  assign n13265 = ~n10384 & ~n10383;
  assign n10387 = ~n11807 | ~P2_REG1_REG_7__SCAN_IN;
  assign n13260 = n10385 ^ P2_REG3_REG_7__SCAN_IN;
  assign n10386 = ~n9035 | ~n13260;
  assign n10389 = ~n11803 | ~P2_REG0_REG_7__SCAN_IN;
  assign n10388 = ~n11804 | ~P2_REG2_REG_7__SCAN_IN;
  assign n15981 = ~n16165 & ~n16166;
  assign n13172 = ~n10394 | ~n10393;
  assign n10408 = ~n15371 & ~n10395;
  assign n10400 = ~n10404 & ~n10608;
  assign n10402 = ~n10400 & ~n10403;
  assign n10401 = ~n10608 & ~P2_IR_REG_8__SCAN_IN;
  assign n10406 = ~n10402 & ~n10401;
  assign n10405 = ~n10426;
  assign n10407 = ~n11632 & ~n11934;
  assign n10414 = ~n11803 | ~P2_REG0_REG_8__SCAN_IN;
  assign n13293 = n10432 ^ P2_REG3_REG_8__SCAN_IN;
  assign n10411 = ~n13293;
  assign n10413 = ~n10412 | ~n10411;
  assign n10416 = ~n11807 | ~P2_REG1_REG_8__SCAN_IN;
  assign n10415 = ~n10476 | ~P2_REG2_REG_8__SCAN_IN;
  assign n16181 = ~n16160 | ~n16161;
  assign n10420 = ~n13172 | ~n16181;
  assign n13312 = ~n10420 | ~n10419;
  assign n10421 = ~P1_DATAO_REG_9__SCAN_IN;
  assign n10429 = ~n15371 & ~n10421;
  assign n10422 = ~n10426 | ~P2_IR_REG_31__SCAN_IN;
  assign n10425 = ~n10422 | ~P2_IR_REG_9__SCAN_IN;
  assign n10423 = ~P2_IR_REG_9__SCAN_IN;
  assign n10424 = ~n10423 | ~P2_IR_REG_31__SCAN_IN;
  assign n10427 = ~n10425 | ~n10424;
  assign n10428 = ~n11632 & ~n11944;
  assign n16176 = ~n10431 | ~n10430;
  assign n10433 = ~n10432;
  assign n10435 = ~n10433 | ~P2_REG3_REG_8__SCAN_IN;
  assign n10434 = ~P2_REG3_REG_9__SCAN_IN;
  assign n10437 = ~n10435 | ~n10434;
  assign n10458 = ~n10436;
  assign n13549 = ~n10437 | ~n10458;
  assign n10438 = ~n13549;
  assign n10442 = ~n11807 | ~P2_REG1_REG_9__SCAN_IN;
  assign n10441 = ~n10476 | ~P2_REG2_REG_9__SCAN_IN;
  assign n16180 = ~n16176 | ~n16177;
  assign n10446 = ~n13312 | ~n16180;
  assign n10448 = ~P2_IR_REG_10__SCAN_IN;
  assign n10451 = ~n10449 & ~n10448;
  assign n10454 = ~n11967 & ~n11632;
  assign n10452 = ~P1_DATAO_REG_10__SCAN_IN;
  assign n10453 = ~n15371 & ~n10452;
  assign n16205 = ~n10456 | ~n10455;
  assign n10457 = ~P2_REG3_REG_10__SCAN_IN;
  assign n10459 = ~n10458 | ~n10457;
  assign n13683 = ~n10459 | ~n10480;
  assign n10460 = ~n13683;
  assign n10463 = ~n10476 | ~P2_REG2_REG_10__SCAN_IN;
  assign n10467 = ~n16205 | ~n16195;
  assign n10469 = ~n13690 | ~n10467;
  assign n13618 = ~n10469 | ~n10468;
  assign n16188 = ~n10475 | ~n10474;
  assign n13654 = n10480 ^ n10479;
  assign n10487 = ~n10491 | ~P2_IR_REG_31__SCAN_IN;
  assign n10488 = ~P2_IR_REG_12__SCAN_IN;
  assign n10489 = ~n10488 | ~P2_IR_REG_31__SCAN_IN;
  assign n10492 = ~n10532;
  assign n10496 = ~n12311 & ~n11632;
  assign n10495 = ~n15371 & ~n10494;
  assign n16229 = ~n10498 | ~n10497;
  assign n10501 = ~n10499;
  assign n10500 = ~P2_REG3_REG_12__SCAN_IN;
  assign n10502 = ~n10501 | ~n10500;
  assign n14164 = ~n10502 | ~n10519;
  assign n10507 = ~n11807 | ~P2_REG1_REG_12__SCAN_IN;
  assign n10510 = ~n16229 | ~n16230;
  assign n10512 = ~n13719 | ~n10510;
  assign n13902 = ~n10512 | ~n10511;
  assign n14261 = ~n10517 | ~n10516;
  assign n10518 = ~P2_REG3_REG_13__SCAN_IN;
  assign n10520 = ~n10519 | ~n10518;
  assign n14242 = ~n10520 | ~n10538;
  assign n13924 = ~n14242;
  assign n10524 = ~n11807 | ~P2_REG1_REG_13__SCAN_IN;
  assign n10527 = ~n14261 | ~n13988;
  assign n10530 = ~n13902 | ~n10527;
  assign n10528 = ~n14261;
  assign n13993 = ~n10530 | ~n10529;
  assign n16247 = ~n10537 | ~n10536;
  assign n13997 = ~n10538 ^ P2_REG3_REG_14__SCAN_IN;
  assign n10542 = ~n11807 | ~P2_REG1_REG_14__SCAN_IN;
  assign n10541 = ~n9033 | ~P2_REG0_REG_14__SCAN_IN;
  assign n10546 = ~n13993 | ~n13994;
  assign n14063 = ~n10546 | ~n10545;
  assign n16266 = ~n10554 | ~n10553;
  assign n10556 = ~n11803 | ~P2_REG0_REG_15__SCAN_IN;
  assign n10559 = ~n11807 | ~P2_REG1_REG_15__SCAN_IN;
  assign n14087 = n10557 ^ P2_REG3_REG_15__SCAN_IN;
  assign n10558 = ~n9035 | ~n14087;
  assign n10563 = ~n14063 | ~n14070;
  assign n10566 = ~n10564 | ~P2_IR_REG_31__SCAN_IN;
  assign n10572 = ~n11807 | ~P2_REG1_REG_16__SCAN_IN;
  assign n14432 = ~n10593 ^ P2_REG3_REG_16__SCAN_IN;
  assign n10571 = ~n9035 | ~n14432;
  assign n10574 = ~n11803 | ~P2_REG0_REG_16__SCAN_IN;
  assign n10840 = ~n10578 | ~n10577;
  assign n10601 = ~n10840;
  assign n10580 = ~n10579 | ~P2_IR_REG_31__SCAN_IN;
  assign n10583 = ~n10580 | ~P2_IR_REG_17__SCAN_IN;
  assign n10581 = ~P2_IR_REG_17__SCAN_IN;
  assign n10582 = ~n10581 | ~P2_IR_REG_31__SCAN_IN;
  assign n10585 = ~n10583 | ~n10582;
  assign n10584 = ~n10605;
  assign n16053 = ~n10590 & ~n10589;
  assign n13882 = ~P2_REG3_REG_16__SCAN_IN;
  assign n10594 = ~n10593 & ~n13882;
  assign n10595 = ~n10594 & ~P2_REG3_REG_17__SCAN_IN;
  assign n10603 = ~n10601 | ~n10600;
  assign n15884 = ~n16056 | ~n16054;
  assign n16003 = ~n16062 & ~n16063;
  assign n10989 = ~n10603 | ~n10602;
  assign n10617 = ~n12842 | ~n10310;
  assign n10604 = ~P1_DATAO_REG_18__SCAN_IN;
  assign n10607 = ~n10605 & ~n10608;
  assign n10610 = ~n10607 & ~n10606;
  assign n10609 = ~n10608 & ~P2_IR_REG_18__SCAN_IN;
  assign n10613 = ~n10610 & ~n10609;
  assign n10612 = ~n10611;
  assign n16293 = ~n10731 & ~n11788;
  assign n16067 = ~n10626 | ~n10625;
  assign n11086 = ~n10628 | ~n10627;
  assign n10631 = ~n10630 | ~n10629;
  assign n10633 = ~n10632;
  assign n16031 = ~n10638 | ~n10639;
  assign n10885 = ~n9039 | ~n16471;
  assign n10640 = ~n10639 | ~P2_IR_REG_31__SCAN_IN;
  assign n10643 = n10885 & n10886;
  assign n14769 = ~n10643 & ~n10642;
  assign n16084 = ~n12383 & ~n16071;
  assign n12338 = ~n12346 | ~n16084;
  assign n10646 = ~n16070 | ~n12351;
  assign n12594 = ~n12338 | ~n10646;
  assign n10647 = ~n16073 | ~n13050;
  assign n10648 = ~n16076 | ~n16093;
  assign n12895 = ~n10649 | ~n10648;
  assign n10651 = ~n12895 | ~n12889;
  assign n10650 = ~n16124 | ~n13144;
  assign n12999 = ~n10653 & ~n16111;
  assign n10654 = ~n12999 | ~n16132;
  assign n13256 = ~n10654 | ~n16146;
  assign n10655 = ~n13256 | ~n16135;
  assign n13180 = ~n10655 | ~n16148;
  assign n10658 = ~n13180 | ~n13173;
  assign n15887 = ~n10658 | ~n10657;
  assign n10659 = ~n15887 | ~n15890;
  assign n13695 = ~n10659 | ~n15888;
  assign n15892 = ~n16205 | ~n13642;
  assign n10660 = ~n13695 & ~n13689;
  assign n13625 = ~n10660 & ~n15895;
  assign n13729 = ~n10661 & ~n15894;
  assign n13907 = ~n10662 & ~n15902;
  assign n13985 = ~n13907 | ~n10663;
  assign n14052 = ~n13985 | ~n15905;
  assign n10668 = ~n14052 | ~n10667;
  assign n10851 = ~n10668 | ~n16279;
  assign n10669 = ~n10851 | ~n15883;
  assign n10997 = ~n10669 | ~n15884;
  assign n10670 = ~n10997 & ~n16293;
  assign n11112 = ~n10670 & ~n15881;
  assign n16469 = ~n16038 & ~n16491;
  assign n10671 = ~n9039 & ~n16031;
  assign n16299 = ~n10679 | ~n10678;
  assign n11631 = ~n16031 & ~n16491;
  assign n10681 = ~n16299 | ~n15549;
  assign n16488 = ~n11631 | ~n11662;
  assign n10680 = ~n11788 | ~n15550;
  assign n10682 = ~n10681 | ~n10680;
  assign n10687 = ~P2_D_REG_12__SCAN_IN & ~P2_D_REG_13__SCAN_IN;
  assign n10686 = ~P2_D_REG_10__SCAN_IN & ~P2_D_REG_11__SCAN_IN;
  assign n10691 = ~n10687 | ~n10686;
  assign n10689 = ~P2_D_REG_8__SCAN_IN & ~P2_D_REG_9__SCAN_IN;
  assign n10688 = ~P2_D_REG_6__SCAN_IN & ~P2_D_REG_7__SCAN_IN;
  assign n10690 = ~n10689 | ~n10688;
  assign n10713 = n10691 | n10690;
  assign n10693 = ~P2_D_REG_4__SCAN_IN & ~P2_D_REG_5__SCAN_IN;
  assign n10692 = ~P2_D_REG_2__SCAN_IN & ~P2_D_REG_3__SCAN_IN;
  assign n10694 = ~n10693 | ~n10692;
  assign n10711 = ~n10694 & ~P2_D_REG_29__SCAN_IN;
  assign n10696 = ~P2_D_REG_28__SCAN_IN & ~P2_D_REG_31__SCAN_IN;
  assign n10695 = ~P2_D_REG_26__SCAN_IN & ~P2_D_REG_27__SCAN_IN;
  assign n10700 = ~n10696 | ~n10695;
  assign n10698 = ~P2_D_REG_15__SCAN_IN & ~P2_D_REG_17__SCAN_IN;
  assign n10697 = ~P2_D_REG_16__SCAN_IN & ~P2_D_REG_14__SCAN_IN;
  assign n10699 = ~n10698 | ~n10697;
  assign n10708 = ~n10700 & ~n10699;
  assign n10702 = ~P2_D_REG_24__SCAN_IN & ~P2_D_REG_25__SCAN_IN;
  assign n10701 = ~P2_D_REG_22__SCAN_IN & ~P2_D_REG_23__SCAN_IN;
  assign n10706 = ~n10702 | ~n10701;
  assign n10704 = ~P2_D_REG_20__SCAN_IN & ~P2_D_REG_21__SCAN_IN;
  assign n10703 = ~P2_D_REG_18__SCAN_IN & ~P2_D_REG_19__SCAN_IN;
  assign n10705 = ~n10704 | ~n10703;
  assign n10707 = ~n10706 & ~n10705;
  assign n10709 = ~n10708 | ~n10707;
  assign n10710 = ~n10709 & ~P2_D_REG_30__SCAN_IN;
  assign n10712 = ~n10711 | ~n10710;
  assign n10878 = ~n13709 | ~n10725;
  assign n16486 = ~n10880 | ~n11612;
  assign n16468 = ~n12014;
  assign n14995 = ~n16468 | ~n9039;
  assign n12004 = ~n14995 & ~n16038;
  assign n15272 = ~n10885 & ~n16038;
  assign n15285 = ~n9039 & ~n12014;
  assign n10733 = ~n15566 | ~n15914;
  assign n13071 = n15488 | n12806;
  assign n10730 = ~n16125 | ~n13050;
  assign n12899 = ~n12900 & ~n10730;
  assign n10739 = ~n15725 | ~n14640;
  assign n10738 = ~n15488 | ~P2_REG2_REG_19__SCAN_IN;
  assign n10740 = ~n10739 | ~n10738;
  assign P2_U3277 = n10741 | n10740;
  assign n10744 = n10742 | P2_STATE_REG_SCAN_IN;
  assign n10743 = ~P2_IR_REG_0__SCAN_IN | ~P2_STATE_REG_SCAN_IN;
  assign P2_U3358 = ~n10744 | ~n10743;
  assign n10747 = ~n10746 ^ n10745;
  assign n10753 = ~n10747 | ~n10132;
  assign n12521 = ~n13968;
  assign n10748 = ~n12521 | ~n10222;
  assign n10750 = ~n10749 | ~n10748;
  assign n12628 = ~P1_STATE_REG_SCAN_IN | ~n10861;
  assign n10752 = ~P1_REG3_REG_2__SCAN_IN | ~n12628;
  assign n10759 = ~n10753 | ~n10752;
  assign n10755 = ~n15689 & ~n16568;
  assign n10754 = ~n17136 & ~n12550;
  assign n10757 = ~n10755 & ~n10754;
  assign n10756 = ~n15578 | ~n16561;
  assign n10758 = ~n10757 | ~n10756;
  assign P1_U3235 = n10759 | n10758;
  assign n10800 = ~n15766 & ~n12767;
  assign n10762 = ~n12153;
  assign n16981 = ~n13114 ^ n16595;
  assign n16554 = ~n12534 & ~n12934;
  assign n16553 = ~n12629 & ~n12522;
  assign n16563 = ~n16554 & ~n16553;
  assign n16974 = ~n12629 | ~n12522;
  assign n12553 = ~n16976 | ~n16974;
  assign n10767 = ~n16562 & ~n12559;
  assign n10781 = ~n12721 & ~n16561;
  assign n16574 = ~n12721 & ~n12559;
  assign n16896 = ~n10768 & ~n16574;
  assign n16581 = ~n12671 | ~n16567;
  assign n17043 = ~n16581;
  assign n16579 = ~n16568 | ~n12720;
  assign n16971 = ~n17043 & ~n17041;
  assign n10770 = ~n10769 | ~n16971;
  assign n12449 = ~n10770 | ~n16579;
  assign n16888 = ~n12495 | ~n12794;
  assign n16901 = ~n12825 | ~n12668;
  assign n12362 = ~n10771 | ~n16901;
  assign n16890 = ~n12822 | ~n12763;
  assign n16598 = ~n12451 | ~n12435;
  assign n13113 = ~n10772 | ~n16598;
  assign n10775 = n16981 ^ n13113;
  assign n10773 = ~n16847;
  assign n13329 = ~n17037;
  assign n15738 = ~n10773 & ~n16967;
  assign n10777 = ~n10775 & ~n15738;
  assign n10776 = ~n13121 & ~n15595;
  assign n10795 = ~n10777 & ~n10776;
  assign n12167 = ~n12534 | ~n12282;
  assign n10778 = ~n12629 & ~n12542;
  assign n10780 = ~n12167 & ~n10778;
  assign n10779 = ~n12550 & ~n12522;
  assign n12549 = ~n10780 & ~n10779;
  assign n10783 = ~n12549 | ~n16969;
  assign n10782 = ~n10781;
  assign n12500 = ~n12501 | ~n12502;
  assign n16569 = ~n12671 & ~n12720;
  assign n10784 = ~n16569;
  assign n12456 = ~n12500 | ~n10784;
  assign n16972 = ~n16888 | ~n16901;
  assign n10786 = ~n12456 | ~n16972;
  assign n10785 = ~n12825 | ~n12794;
  assign n16590 = ~n12822 | ~n12451;
  assign n10788 = ~n10787 | ~n16590;
  assign n16589 = ~n12435 | ~n12763;
  assign n13100 = ~n10788 | ~n16589;
  assign n12738 = n16981 ^ n13100;
  assign n10789 = ~n16962;
  assign n10790 = ~n10789 | ~n10796;
  assign n10793 = ~n12738 & ~n15404;
  assign n10792 = ~n12451 & ~n15594;
  assign n10794 = ~n10793 & ~n10792;
  assign n12739 = ~n10795 | ~n10794;
  assign n12789 = ~n10796 & ~n17072;
  assign n13107 = ~n12789;
  assign n10797 = ~n12738 & ~n13107;
  assign n10798 = ~n12739 & ~n10797;
  assign n10799 = ~n15218 & ~n10798;
  assign n10802 = ~n10800 & ~n10799;
  assign n10801 = ~n15218 | ~P1_REG2_REG_6__SCAN_IN;
  assign n10809 = ~n10802 | ~n10801;
  assign n15174 = ~n15745 | ~n14237;
  assign n12560 = ~n12542 & ~n12282;
  assign n12506 = ~n12560 | ~n12559;
  assign n12505 = ~n12506 & ~n12720;
  assign n10803 = ~n12435 & ~n12668;
  assign n10804 = ~n12505 | ~n10803;
  assign n13365 = ~n10804 & ~n13114;
  assign n12370 = ~n10804;
  assign n16596 = ~n13114;
  assign n10805 = ~n12370 & ~n16596;
  assign n12735 = ~n13365 & ~n10805;
  assign n10807 = ~n15762 | ~n12735;
  assign n10806 = ~n15313 | ~n13114;
  assign n10808 = ~n10807 | ~n10806;
  assign P1_U3285 = n10809 | n10808;
  assign n10839 = ~n10810 ^ P2_ADDR_REG_19__SCAN_IN;
  assign n10837 = ~P1_ADDR_REG_18__SCAN_IN & ~P2_ADDR_REG_18__SCAN_IN;
  assign n13386 = P1_ADDR_REG_17__SCAN_IN & P2_ADDR_REG_17__SCAN_IN;
  assign n13195 = P1_ADDR_REG_16__SCAN_IN & P2_ADDR_REG_16__SCAN_IN;
  assign n12834 = P1_ADDR_REG_15__SCAN_IN & P2_ADDR_REG_15__SCAN_IN;
  assign n12571 = P2_ADDR_REG_14__SCAN_IN & P1_ADDR_REG_14__SCAN_IN;
  assign n12319 = P2_ADDR_REG_13__SCAN_IN & P1_ADDR_REG_13__SCAN_IN;
  assign n12138 = P2_ADDR_REG_12__SCAN_IN & P1_ADDR_REG_12__SCAN_IN;
  assign n12000 = P2_ADDR_REG_11__SCAN_IN & P1_ADDR_REG_11__SCAN_IN;
  assign n11812 = P2_ADDR_REG_10__SCAN_IN & P1_ADDR_REG_10__SCAN_IN;
  assign n10827 = ~P2_ADDR_REG_9__SCAN_IN & ~P1_ADDR_REG_9__SCAN_IN;
  assign n10825 = ~P2_ADDR_REG_8__SCAN_IN & ~P1_ADDR_REG_8__SCAN_IN;
  assign n10823 = ~P2_ADDR_REG_7__SCAN_IN & ~P1_ADDR_REG_7__SCAN_IN;
  assign n10821 = ~P1_ADDR_REG_6__SCAN_IN | ~P2_ADDR_REG_6__SCAN_IN;
  assign n11379 = P1_ADDR_REG_6__SCAN_IN ^ P2_ADDR_REG_6__SCAN_IN;
  assign n10819 = ~P2_ADDR_REG_5__SCAN_IN & ~P1_ADDR_REG_5__SCAN_IN;
  assign n10817 = ~P2_ADDR_REG_4__SCAN_IN & ~P1_ADDR_REG_4__SCAN_IN;
  assign n10815 = ~P1_ADDR_REG_3__SCAN_IN | ~P2_ADDR_REG_3__SCAN_IN;
  assign n11356 = P1_ADDR_REG_3__SCAN_IN ^ P2_ADDR_REG_3__SCAN_IN;
  assign n10813 = ~P1_ADDR_REG_2__SCAN_IN | ~P2_ADDR_REG_2__SCAN_IN;
  assign n11348 = P1_ADDR_REG_0__SCAN_IN & P2_ADDR_REG_0__SCAN_IN;
  assign n11351 = ~P1_ADDR_REG_1__SCAN_IN & ~n11348;
  assign n11350 = P1_ADDR_REG_1__SCAN_IN & n11348;
  assign n10811 = ~P2_ADDR_REG_1__SCAN_IN & ~n11350;
  assign n11354 = ~n11351 & ~n10811;
  assign n11353 = P1_ADDR_REG_2__SCAN_IN ^ P2_ADDR_REG_2__SCAN_IN;
  assign n10812 = ~n11354 | ~n11353;
  assign n11355 = ~n10813 | ~n10812;
  assign n10814 = ~n11356 | ~n11355;
  assign n11360 = ~P2_ADDR_REG_4__SCAN_IN ^ P1_ADDR_REG_4__SCAN_IN;
  assign n10816 = ~n11361 & ~n11360;
  assign n11362 = ~P2_ADDR_REG_5__SCAN_IN ^ P1_ADDR_REG_5__SCAN_IN;
  assign n10818 = ~n11363 & ~n11362;
  assign n11435 = ~P2_ADDR_REG_7__SCAN_IN ^ P1_ADDR_REG_7__SCAN_IN;
  assign n11543 = ~P2_ADDR_REG_8__SCAN_IN ^ P1_ADDR_REG_8__SCAN_IN;
  assign n11732 = ~P2_ADDR_REG_9__SCAN_IN ^ P1_ADDR_REG_9__SCAN_IN;
  assign n11813 = ~P2_ADDR_REG_10__SCAN_IN & ~P1_ADDR_REG_10__SCAN_IN;
  assign n12001 = ~P2_ADDR_REG_11__SCAN_IN & ~P1_ADDR_REG_11__SCAN_IN;
  assign n12139 = ~P2_ADDR_REG_12__SCAN_IN & ~P1_ADDR_REG_12__SCAN_IN;
  assign n12320 = ~P2_ADDR_REG_13__SCAN_IN & ~P1_ADDR_REG_13__SCAN_IN;
  assign n12572 = ~P2_ADDR_REG_14__SCAN_IN & ~P1_ADDR_REG_14__SCAN_IN;
  assign n12835 = ~P1_ADDR_REG_15__SCAN_IN & ~P2_ADDR_REG_15__SCAN_IN;
  assign n13196 = ~P1_ADDR_REG_16__SCAN_IN & ~P2_ADDR_REG_16__SCAN_IN;
  assign n13387 = ~P1_ADDR_REG_17__SCAN_IN & ~P2_ADDR_REG_17__SCAN_IN;
  assign n13547 = ~P1_ADDR_REG_18__SCAN_IN ^ P2_ADDR_REG_18__SCAN_IN;
  assign n10836 = ~n13548 & ~n13547;
  assign n10838 = ~n10837 & ~n10836;
  assign ADD_1071_U4 = n10839 ^ n10838;
  assign n10843 = ~n15566 | ~n16056;
  assign n10842 = ~n15725 | ~n11007;
  assign n10848 = ~n10843 | ~n10842;
  assign n14205 = n10846 | n10992;
  assign n10847 = ~n14079 & ~n14205;
  assign n10854 = ~n14642 & ~n15713;
  assign n10853 = ~n16285 & ~n16488;
  assign n10855 = ~n10854 & ~n10853;
  assign n10857 = ~n15720 & ~P2_REG2_REG_17__SCAN_IN;
  assign P2_U3279 = n10860 | n10859;
  assign n14853 = ~n10861 & ~P1_U3084;
  assign n10876 = ~n14796 & ~n14136;
  assign n10872 = ~n16700 & ~n17126;
  assign n10868 = ~n17136 & ~n14151;
  assign n13465 = ~n10867 & ~P1_STATE_REG_SCAN_IN;
  assign n10870 = ~n10868 & ~n13465;
  assign n10869 = ~n17132 | ~n16693;
  assign n10871 = ~n10870 | ~n10869;
  assign n10873 = ~n10872 & ~n10871;
  assign P1_U3239 = n10876 | n10875;
  assign n10960 = ~n12008 & ~n10877;
  assign n10879 = ~n10878;
  assign n10954 = ~n13997 | ~n15530;
  assign n16039 = ~n11631;
  assign n10975 = ~n16244 & ~n10888;
  assign n10890 = ~n16070 & ~n10888;
  assign n12386 = ~n12345 | ~n12806;
  assign n10889 = ~n16071 | ~n11296;
  assign n12326 = n12386 & n10889;
  assign n12327 = ~n12325 | ~n12326;
  assign n10893 = ~n10890;
  assign n12416 = ~n12327 | ~n10894;
  assign n10895 = n13050 ^ n11318;
  assign n12414 = ~n12416 & ~n12415;
  assign n10896 = ~n10895;
  assign n10898 = ~n10897 & ~n10896;
  assign n12405 = ~n12414 & ~n10898;
  assign n10899 = ~n16124 & ~n10888;
  assign n10900 = n13144 ^ n11318;
  assign n10903 = ~n12405 & ~n12406;
  assign n10902 = ~n10901 & ~n10900;
  assign n10905 = n12687 ^ n11296;
  assign n12617 = n10904 ^ n10905;
  assign n12619 = ~n12618 | ~n12617;
  assign n10907 = ~n10904;
  assign n10906 = ~n10905;
  assign n10908 = ~n10907 | ~n10906;
  assign n10909 = ~n13078 ^ n11296;
  assign n10910 = ~n13014 | ~n12806;
  assign n12650 = n10909 ^ n10910;
  assign n12649 = ~n12651 & ~n12650;
  assign n10911 = ~n10909;
  assign n10912 = ~n10911 & ~n10910;
  assign n10913 = n13032 ^ n11318;
  assign n10914 = ~n12646 & ~n10888;
  assign n10917 = ~n13024 | ~n13021;
  assign n10916 = ~n10913;
  assign n10915 = ~n10914;
  assign n10919 = ~n13017 & ~n10888;
  assign n10921 = ~n10918;
  assign n10920 = ~n10919;
  assign n10924 = ~n13317 & ~n10888;
  assign n10927 = ~n13297 | ~n13294;
  assign n10926 = ~n10923;
  assign n10925 = ~n10924;
  assign n10929 = ~n16209 & ~n10888;
  assign n10930 = ~n10929;
  assign n13520 = ~n13556 | ~n10934;
  assign n10936 = ~n13642 & ~n10888;
  assign n10939 = ~n13520 | ~n13517;
  assign n10937 = ~n10936;
  assign n13648 = ~n10939 | ~n13518;
  assign n10942 = ~n16189 | ~n12806;
  assign n10945 = ~n10940 | ~n13646;
  assign n10943 = ~n10942;
  assign n10946 = ~n16230 | ~n12806;
  assign n14170 = ~n14248 | ~n14171;
  assign n10949 = ~n13988 | ~n12806;
  assign n10951 = ~n14170 | ~n10948;
  assign n10955 = ~n16486 & ~n15713;
  assign n15535 = ~n10960 | ~n10955;
  assign n10958 = ~n15535 & ~n10956;
  assign n12926 = ~P2_STATE_REG_SCAN_IN & ~n10957;
  assign n10962 = n10958 | n12926;
  assign n10959 = ~n16486 & ~n16488;
  assign n15872 = ~n10960 | ~n10959;
  assign n10961 = ~n15872 & ~n14167;
  assign n10967 = ~n10962 & ~n10961;
  assign n10966 = ~n15867 | ~n16247;
  assign n10968 = ~n10967 | ~n10966;
  assign P2_U3217 = n10969 | n10968;
  assign n10971 = ~n15530 | ~n14087;
  assign n10970 = ~n15867 | ~n16266;
  assign n10988 = ~n10971 | ~n10970;
  assign n10979 = ~n10973 | ~n10972;
  assign n10976 = ~n10975;
  assign n14436 = n11012 | n11014;
  assign n14434 = ~n11012 | ~n11014;
  assign n11017 = ~n16265 | ~n12806;
  assign n10982 = ~n15532 | ~n16248;
  assign n13529 = ~P2_REG3_REG_15__SCAN_IN | ~P2_U3152;
  assign n10984 = ~n10982 | ~n13529;
  assign n10983 = ~n15535 & ~n16285;
  assign n10985 = ~n10984 & ~n10983;
  assign P2_U3243 = n10988 | n10987;
  assign n10991 = ~n15566 | ~n14510;
  assign n10990 = ~n15725 | ~n14505;
  assign n10994 = ~n10991 | ~n10990;
  assign n10993 = ~n13071 & ~n14458;
  assign n11000 = ~n15913 & ~n15713;
  assign n10999 = ~n16054 & ~n16488;
  assign n11001 = ~n11000 & ~n10999;
  assign n11003 = ~n15720 & ~P2_REG2_REG_18__SCAN_IN;
  assign P2_U3278 = n11006 | n11005;
  assign n11009 = ~n15530 | ~n11007;
  assign n11008 = ~n15867 | ~n16056;
  assign n14437 = ~n16277 | ~n12806;
  assign n11023 = ~n11012 & ~n11011;
  assign n11018 = ~n11017 & ~n14437;
  assign n11205 = ~n16054 & ~n10888;
  assign n11026 = ~n15869 | ~n11788;
  assign n14415 = ~P2_REG3_REG_17__SCAN_IN | ~P2_U3152;
  assign n11028 = ~n11026 | ~n14415;
  assign n11027 = ~n15872 & ~n16285;
  assign n11029 = ~n11028 & ~n11027;
  assign P2_U3230 = n11032 | n11031;
  assign n11039 = n11089 & P1_DATAO_REG_28__SCAN_IN;
  assign n11041 = ~n11039 & ~n11038;
  assign n11040 = ~SI_28_;
  assign n11045 = ~n11042 & ~SI_28_;
  assign n11302 = ~n11043 & ~n11045;
  assign n11048 = ~n9034 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n11047 = ~n11089 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n11051 = ~n14575 | ~n14574;
  assign n11050 = ~n11049 | ~SI_29_;
  assign n11053 = ~n9034 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n11052 = ~n11089 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n14384 = ~n9034 | ~P1_U3084;
  assign n11056 = ~n11054 | ~P1_STATE_REG_SCAN_IN;
  assign n14585 = ~n11089 | ~P1_U3084;
  assign n11055 = ~n14388 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n11057 = ~n11056 | ~n11055;
  assign P1_U3323 = n11058 | n11057;
  assign n11063 = ~n11061 | ~P2_STATE_REG_SCAN_IN;
  assign n11062 = ~n14577 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n11064 = ~n11063 | ~n11062;
  assign P2_U3328 = n11065 | n11064;
  assign n11070 = ~n11066 | ~SI_30_;
  assign n11069 = ~n11068 | ~n11067;
  assign n11072 = ~n9034 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n11071 = ~n11089 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n11073 = ~n11072 | ~n11071;
  assign n11076 = ~P1_IR_REG_30__SCAN_IN;
  assign n11077 = ~n11076 | ~P1_IR_REG_31__SCAN_IN;
  assign n11078 = ~n11077 & ~P1_U3084;
  assign n11081 = ~n11079 | ~n11078;
  assign n11080 = ~n14388 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n11082 = ~n11081 | ~n11080;
  assign P1_U3322 = n11083 | n11082;
  assign n11088 = ~n11086 | ~n11085;
  assign n14768 = ~n11088 | ~n11087;
  assign n11095 = ~n14768 | ~n11093;
  assign n11109 = ~n11095 | ~n11094;
  assign n11108 = ~n11109;
  assign n13335 = ~P1_DATAO_REG_21__SCAN_IN;
  assign n16322 = ~n11105 | ~n11104;
  assign n11142 = ~n11108 | ~n11115;
  assign n11110 = ~n11109 | ~n16010;
  assign n14994 = ~n11142 | ~n11110;
  assign n16294 = ~n15914 & ~n15913;
  assign n14770 = ~n11113 & ~n16294;
  assign n15916 = ~n16302 & ~n16299;
  assign n11114 = ~n14770 & ~n15916;
  assign n11185 = ~n11114 & ~n15918;
  assign n11125 = ~n16299 | ~n15550;
  assign n16334 = ~n11123 | ~n11122;
  assign n11124 = ~n16334 | ~n15549;
  assign n11126 = ~n11125 | ~n11124;
  assign n11133 = ~n15566 | ~n16321;
  assign n11132 = ~n15725 | ~n14895;
  assign P2_U3275 = n11140 | n11139;
  assign n15025 = ~n11142 | ~n11141;
  assign n11143 = ~P1_DATAO_REG_22__SCAN_IN;
  assign n15926 = ~n16333 & ~n16338;
  assign n16012 = ~n11147 | ~n11146;
  assign n15024 = ~n15025 | ~n16012;
  assign n15101 = ~n15024 | ~n11148;
  assign n11151 = ~n13708 & ~n9036;
  assign n11149 = ~P1_DATAO_REG_23__SCAN_IN;
  assign n16014 = ~n11160 & ~n11159;
  assign n15099 = ~n15101 | ~n15100;
  assign n11172 = ~n15099 | ~n11161;
  assign n11162 = ~P1_DATAO_REG_24__SCAN_IN;
  assign n16363 = ~n11171 | ~n11170;
  assign n16016 = ~n15274 | ~n15276;
  assign n11173 = n11172 | n16016;
  assign n15242 = ~n11173 | ~n15269;
  assign n11178 = ~n11176 | ~n16500;
  assign n15244 = n11178 | n15283;
  assign n11179 = ~n15725 | ~n15439;
  assign n11186 = ~n11185 | ~n15920;
  assign n15028 = ~n11186 | ~n15922;
  assign n11187 = ~n15028 & ~n15924;
  assign n15275 = ~n11188 | ~n15930;
  assign n11198 = ~n15030 & ~n16488;
  assign n15463 = ~n11196 | ~n11195;
  assign n11197 = ~n16379 & ~n15713;
  assign n11199 = ~n11198 & ~n11197;
  assign P2_U3272 = n11204 | n11203;
  assign n11206 = ~n11207 & ~n11208;
  assign n11210 = ~n11207;
  assign n11211 = ~n11210 & ~n11209;
  assign n14518 = ~n11212 & ~n11211;
  assign n11214 = ~n11788 | ~n12806;
  assign n14637 = ~n11217 | ~n14515;
  assign n11219 = ~n15913 & ~n10888;
  assign n14718 = ~n11222 & ~n11221;
  assign n11224 = ~n16299 | ~n12806;
  assign n14893 = ~n11227 | ~n14716;
  assign n14890 = ~n16322 | ~n12806;
  assign n11230 = ~n14893;
  assign n11231 = ~n11230 | ~n11229;
  assign n15012 = ~n11232 | ~n11231;
  assign n11233 = ~n15012 & ~n15010;
  assign n15009 = ~n16338 & ~n10888;
  assign n11237 = ~n11233 & ~n15009;
  assign n11235 = ~n15012;
  assign n15140 = ~n11237 & ~n11236;
  assign n15137 = ~n16347 | ~n12806;
  assign n11242 = ~n11238 | ~n15137;
  assign n11240 = ~n15140;
  assign n11241 = ~n11240 | ~n11239;
  assign n15436 = ~n16367 & ~n10888;
  assign n11247 = ~n15434 | ~n15436;
  assign n11246 = ~n11243;
  assign n15435 = ~n11246 | ~n11245;
  assign n15526 = ~n11247 | ~n15435;
  assign n11249 = ~n13943 & ~n9036;
  assign n13944 = ~P1_DATAO_REG_25__SCAN_IN;
  assign n15523 = ~n16379 & ~n10888;
  assign n11253 = ~n15526 & ~n11252;
  assign n11291 = ~n11254 & ~n11253;
  assign n11256 = ~n14095 & ~n9036;
  assign n11258 = ~n11807 | ~P2_REG1_REG_26__SCAN_IN;
  assign n11266 = ~n15557 | ~n12806;
  assign n11289 = ~n11269 & ~n15861;
  assign n11279 = ~P2_REG3_REG_26__SCAN_IN;
  assign n11272 = ~n11807 | ~P2_REG1_REG_27__SCAN_IN;
  assign n11271 = ~n11804 | ~P2_REG2_REG_27__SCAN_IN;
  assign n11273 = ~P2_REG0_REG_27__SCAN_IN;
  assign n11275 = ~n11274 & ~n11273;
  assign n15704 = ~n11278 | ~n11277;
  assign n11287 = ~n15704 | ~n15869;
  assign n11283 = ~n15530 | ~n15473;
  assign n11281 = ~n15872 & ~n16379;
  assign n11280 = ~n11279 & ~P2_STATE_REG_SCAN_IN;
  assign n11282 = ~n11281 & ~n11280;
  assign n11284 = ~n11283 | ~n11282;
  assign P2_U3242 = n11289 | n11288;
  assign n11293 = ~n11291 | ~n11290;
  assign n15860 = ~n11293 | ~n11292;
  assign n11297 = ~n16405 & ~n10888;
  assign n11295 = ~n14385 & ~n9036;
  assign n14198 = ~P1_DATAO_REG_27__SCAN_IN;
  assign n15863 = ~n15860 | ~n15859;
  assign n15202 = ~n11306 | ~n11305;
  assign n11310 = ~n11807 | ~P2_REG1_REG_28__SCAN_IN;
  assign n11309 = ~n9033 | ~P2_REG0_REG_28__SCAN_IN;
  assign n11317 = n11310 & n11309;
  assign n15868 = ~n11317 | ~n11316;
  assign n11319 = ~n15868 | ~n12806;
  assign n11343 = ~n15863 | ~n11322;
  assign n11339 = ~n16405 & ~n15872;
  assign n11337 = ~n15777 | ~n15867;
  assign n11335 = n15530 & n15724;
  assign n11326 = ~n11807 | ~P2_REG1_REG_29__SCAN_IN;
  assign n11325 = ~n11803 | ~P2_REG0_REG_29__SCAN_IN;
  assign n11331 = n11326 & n11325;
  assign n11328 = ~n11804 | ~P2_REG2_REG_29__SCAN_IN;
  assign n11333 = ~n15869 | ~n16427;
  assign n11332 = ~P2_REG3_REG_28__SCAN_IN | ~P2_U3152;
  assign n11334 = ~n11333 | ~n11332;
  assign n11336 = ~n11335 & ~n11334;
  assign n11347 = ~n11343 | ~n11342;
  assign n11346 = ~n15863 & ~n11345;
  assign P2_U3222 = n11347 | n11346;
  assign U126 = ~P1_RD_REG_SCAN_IN ^ P2_RD_REG_SCAN_IN;
  assign U123 = ~P1_WR_REG_SCAN_IN ^ P2_WR_REG_SCAN_IN;
  assign n11349 = ~P1_ADDR_REG_0__SCAN_IN & ~P2_ADDR_REG_0__SCAN_IN;
  assign ADD_1071_U46 = ~n11349 & ~n11348;
  assign n11352 = ~n11351 & ~n11350;
  assign ADD_1071_U5 = n11352 ^ P2_ADDR_REG_1__SCAN_IN;
  assign ADD_1071_U54 = n11354 ^ n11353;
  assign ADD_1071_U53 = n11356 ^ n11355;
  assign n11359 = ~n11357 | ~P1_U3084;
  assign n11358 = ~P1_IR_REG_0__SCAN_IN | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3353 = ~n11359 | ~n11358;
  assign ADD_1071_U52 = ~n11361 ^ n11360;
  assign ADD_1071_U51 = ~n11363 ^ n11362;
  assign n11367 = ~P1_D_REG_1__SCAN_IN & ~n11372;
  assign n11366 = ~n11369 & ~n11365;
  assign P1_U3441 = ~n11367 & ~n11366;
  assign n11371 = ~P1_D_REG_0__SCAN_IN & ~n11372;
  assign n11370 = ~n11369 & ~n11368;
  assign P1_U3440 = ~n11371 & ~n11370;
  assign P1_U3320 = P1_D_REG_3__SCAN_IN & n11373;
  assign P1_U3293 = P1_D_REG_30__SCAN_IN & n11373;
  assign P1_U3298 = P1_D_REG_25__SCAN_IN & n11373;
  assign P1_U3319 = P1_D_REG_4__SCAN_IN & n11373;
  assign P1_U3300 = P1_D_REG_23__SCAN_IN & n11373;
  assign P1_U3301 = P1_D_REG_22__SCAN_IN & n11373;
  assign P1_U3302 = P1_D_REG_21__SCAN_IN & n11373;
  assign P1_U3311 = P1_D_REG_12__SCAN_IN & n11373;
  assign P1_U3310 = P1_D_REG_13__SCAN_IN & n11373;
  assign P1_U3292 = P1_D_REG_31__SCAN_IN & n11373;
  assign P1_U3303 = P1_D_REG_20__SCAN_IN & n11373;
  assign P1_U3294 = P1_D_REG_29__SCAN_IN & n11373;
  assign P1_U3295 = P1_D_REG_28__SCAN_IN & n11373;
  assign P1_U3306 = P1_D_REG_17__SCAN_IN & n11373;
  assign P1_U3299 = P1_D_REG_24__SCAN_IN & n11373;
  assign P1_U3321 = P1_D_REG_2__SCAN_IN & n11373;
  assign P1_U3317 = P1_D_REG_6__SCAN_IN & n11373;
  assign P1_U3305 = P1_D_REG_18__SCAN_IN & n11373;
  assign P1_U3296 = P1_D_REG_27__SCAN_IN & n11373;
  assign P1_U3297 = P1_D_REG_26__SCAN_IN & n11373;
  assign P1_U3318 = P1_D_REG_5__SCAN_IN & n11373;
  assign P1_U3312 = P1_D_REG_11__SCAN_IN & n11373;
  assign P1_U3316 = P1_D_REG_7__SCAN_IN & n11373;
  assign P1_U3315 = P1_D_REG_8__SCAN_IN & n11373;
  assign P1_U3314 = P1_D_REG_9__SCAN_IN & n11373;
  assign P1_U3313 = P1_D_REG_10__SCAN_IN & n11373;
  assign P1_U3308 = P1_D_REG_15__SCAN_IN & n11373;
  assign P1_U3307 = P1_D_REG_16__SCAN_IN & n11373;
  assign P1_U3309 = P1_D_REG_14__SCAN_IN & n11373;
  assign P1_U3304 = P1_D_REG_19__SCAN_IN & n11373;
  assign n11375 = ~n11386 & ~n14384;
  assign n11374 = ~n11428 & ~P1_U3084;
  assign n11377 = ~n11375 & ~n11374;
  assign n11376 = ~n14388 | ~P2_DATAO_REG_3__SCAN_IN;
  assign P1_U3350 = ~n11377 | ~n11376;
  assign ADD_1071_U50 = n11379 ^ n11378;
  assign n11381 = ~n12534 | ~P1_U4006;
  assign n11380 = ~n12117 | ~P1_DATAO_REG_0__SCAN_IN;
  assign P1_U3555 = ~n11381 | ~n11380;
  assign n11383 = ~n13818 | ~P1_U4006;
  assign n11382 = ~n12117 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P1_U3566 = ~n11383 | ~n11382;
  assign n11385 = ~n13783 | ~P1_U4006;
  assign n11384 = ~n12117 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P1_U3565 = ~n11385 | ~n11384;
  assign n11388 = ~n11386 & ~n14094;
  assign n11387 = ~n11657 & ~P2_U3152;
  assign n11390 = ~n11388 & ~n11387;
  assign n11389 = ~n14577 | ~P1_DATAO_REG_3__SCAN_IN;
  assign P2_U3355 = ~n11390 | ~n11389;
  assign n11392 = ~n12671 | ~P1_U4006;
  assign n11391 = ~n12117 | ~P1_DATAO_REG_3__SCAN_IN;
  assign P1_U3558 = ~n11392 | ~n11391;
  assign n11394 = ~n12721 | ~P1_U4006;
  assign n11393 = ~n12117 | ~P1_DATAO_REG_2__SCAN_IN;
  assign P1_U3557 = ~n11394 | ~n11393;
  assign n11399 = ~n11480 | ~n14582;
  assign n11397 = ~n11452 & ~P1_U3084;
  assign n11396 = ~n14585 & ~n11395;
  assign n11398 = ~n11397 & ~n11396;
  assign P1_U3349 = ~n11399 | ~n11398;
  assign n11403 = ~n11486 | ~n14582;
  assign n11401 = ~n14388 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n11584 = ~n11424;
  assign n11400 = ~n11584 | ~P1_STATE_REG_SCAN_IN;
  assign n11402 = n11401 & n11400;
  assign P1_U3352 = ~n11403 | ~n11402;
  assign n11405 = ~n16717 | ~P1_U4006;
  assign n11404 = ~n12117 | ~P1_DATAO_REG_17__SCAN_IN;
  assign P1_U3572 = ~n11405 | ~n11404;
  assign n11407 = ~n12629 | ~P1_U4006;
  assign n11406 = ~n12117 | ~P1_DATAO_REG_1__SCAN_IN;
  assign P1_U3556 = ~n11407 | ~n11406;
  assign n12726 = ~P1_REG3_REG_3__SCAN_IN | ~P1_U3084;
  assign n11570 = ~n11424 ^ P1_REG1_REG_1__SCAN_IN;
  assign n11569 = P1_IR_REG_0__SCAN_IN & P1_REG1_REG_0__SCAN_IN;
  assign n11572 = ~n11570 | ~n11569;
  assign n11408 = ~n11584 | ~P1_REG1_REG_1__SCAN_IN;
  assign n11852 = ~n11572 | ~n11408;
  assign n11851 = n11859 ^ P1_REG1_REG_2__SCAN_IN;
  assign n11853 = ~n11852 | ~n11851;
  assign n11409 = ~n11859 | ~P1_REG1_REG_2__SCAN_IN;
  assign n11413 = ~n11853 | ~n11409;
  assign n11412 = ~n11428 ^ P1_REG1_REG_3__SCAN_IN;
  assign n11411 = ~n11413 & ~n11412;
  assign n14411 = ~n11846 & ~P1_U3084;
  assign n11410 = n14411 & n11845;
  assign n11414 = ~n11411 & ~n14833;
  assign n11444 = ~n11413 | ~n11412;
  assign n11415 = ~n11414 | ~n11444;
  assign n11421 = ~n12726 | ~n11415;
  assign n17096 = ~n11416 & ~n17092;
  assign n14842 = ~P1_U3083 & ~n17096;
  assign n11419 = ~n14842 | ~P1_ADDR_REG_3__SCAN_IN;
  assign n14386 = ~n11845 & ~P1_U3084;
  assign n11422 = ~n11417 | ~n14386;
  assign n14837 = ~n11422 & ~n11423;
  assign n11449 = ~n11428;
  assign n11418 = ~n14837 | ~n11449;
  assign n11420 = ~n11419 | ~n11418;
  assign n11434 = ~n11421 & ~n11420;
  assign n11492 = ~n11422;
  assign n11836 = ~P1_REG2_REG_0__SCAN_IN;
  assign n11838 = ~n9044 & ~n11836;
  assign n11576 = ~n11424 ^ P1_REG2_REG_1__SCAN_IN;
  assign n11578 = ~n11838 | ~n11576;
  assign n11425 = ~n11584 | ~P1_REG2_REG_1__SCAN_IN;
  assign n11857 = ~n11578 | ~n11425;
  assign n11856 = n11859 ^ P1_REG2_REG_2__SCAN_IN;
  assign n11427 = ~n11857 | ~n11856;
  assign n11426 = ~n11859 | ~P1_REG2_REG_2__SCAN_IN;
  assign n11431 = ~n11427 | ~n11426;
  assign n11430 = ~n11428 ^ P1_REG2_REG_3__SCAN_IN;
  assign n11429 = ~n11431 & ~n11430;
  assign n11432 = ~n14825 & ~n11429;
  assign n11451 = ~n11431 | ~n11430;
  assign n11433 = ~n11432 | ~n11451;
  assign P1_U3244 = ~n11434 | ~n11433;
  assign ADD_1071_U49 = ~n11436 ^ n11435;
  assign n11463 = ~n11612;
  assign n11438 = ~P2_D_REG_0__SCAN_IN | ~n11463;
  assign n11437 = ~n11612 | ~n12020;
  assign P2_U3437 = ~n11438 | ~n11437;
  assign n11440 = ~n11545 | ~n14582;
  assign n11439 = ~n11859 | ~P1_STATE_REG_SCAN_IN;
  assign n11442 = n11440 & n11439;
  assign n11441 = ~n14388 | ~P2_DATAO_REG_2__SCAN_IN;
  assign P1_U3351 = ~n11442 | ~n11441;
  assign n12766 = ~P1_REG3_REG_6__SCAN_IN | ~P1_U3084;
  assign n11443 = ~n11449 | ~P1_REG1_REG_3__SCAN_IN;
  assign n11911 = ~n11444 | ~n11443;
  assign n11910 = ~n11452 ^ P1_REG1_REG_4__SCAN_IN;
  assign n11912 = ~n11911 | ~n11910;
  assign n11907 = ~n11452;
  assign n11445 = ~n11907 | ~P1_REG1_REG_4__SCAN_IN;
  assign n11556 = ~n11912 | ~n11445;
  assign n11555 = ~n11469 ^ P1_REG1_REG_5__SCAN_IN;
  assign n11557 = ~n11556 | ~n11555;
  assign n11446 = ~n11562 | ~P1_REG1_REG_5__SCAN_IN;
  assign n11515 = n11532 ^ P1_REG1_REG_6__SCAN_IN;
  assign n11447 = ~n11516 ^ n11515;
  assign n11448 = ~n11447 | ~n14333;
  assign n11460 = ~n12766 | ~n11448;
  assign n11450 = ~n11449 | ~P1_REG2_REG_3__SCAN_IN;
  assign n11905 = ~n11451 | ~n11450;
  assign n11904 = ~n11452 ^ P1_REG2_REG_4__SCAN_IN;
  assign n11454 = ~n11905 | ~n11904;
  assign n11453 = ~n11907 | ~P1_REG2_REG_4__SCAN_IN;
  assign n11551 = ~n11454 | ~n11453;
  assign n11550 = ~n11469 ^ P1_REG2_REG_5__SCAN_IN;
  assign n11552 = ~n11551 | ~n11550;
  assign n11455 = ~n11562 | ~P1_REG2_REG_5__SCAN_IN;
  assign n11508 = ~n11552 | ~n11455;
  assign n11507 = ~n11532 ^ P1_REG2_REG_6__SCAN_IN;
  assign n11456 = n11508 ^ n11507;
  assign n11458 = ~n11456 | ~n14325;
  assign n11517 = ~n11532;
  assign n11457 = ~n14837 | ~n11517;
  assign n11459 = ~n11458 | ~n11457;
  assign n11462 = ~n11460 & ~n11459;
  assign n11461 = ~n14842 | ~P1_ADDR_REG_6__SCAN_IN;
  assign P1_U3247 = ~n11462 | ~n11461;
  assign n11466 = ~P2_D_REG_1__SCAN_IN | ~n11463;
  assign n11465 = ~n11612 | ~n11464;
  assign P2_U3438 = ~n11466 | ~n11465;
  assign n11468 = ~P1_DATAO_REG_19__SCAN_IN | ~n12117;
  assign n11467 = ~P1_U4006 | ~n16534;
  assign P1_U3574 = ~n11468 | ~n11467;
  assign n11471 = ~n11474 & ~n14384;
  assign n11470 = ~n11469 & ~P1_U3084;
  assign n11473 = ~n11471 & ~n11470;
  assign n11472 = ~n14388 | ~P2_DATAO_REG_5__SCAN_IN;
  assign P1_U3348 = ~n11473 | ~n11472;
  assign n11477 = ~n11474 & ~n14094;
  assign n11476 = ~n11475 & ~P2_U3152;
  assign n11479 = ~n11477 & ~n11476;
  assign n11478 = ~n14577 | ~P1_DATAO_REG_5__SCAN_IN;
  assign P2_U3353 = ~n11479 | ~n11478;
  assign n11485 = ~n11480 | ~n11059;
  assign n11483 = ~n11659 & ~P2_U3152;
  assign n11482 = ~n14962 & ~n11481;
  assign n11484 = ~n11483 & ~n11482;
  assign P2_U3354 = ~n11485 | ~n11484;
  assign n11491 = ~n11486 | ~n11059;
  assign n11489 = ~n14962 & ~n11487;
  assign n11488 = ~n11653 & ~P2_U3152;
  assign n11490 = ~n11489 & ~n11488;
  assign P2_U3357 = ~n11491 | ~n11490;
  assign n11496 = ~n14833 & ~P1_REG1_REG_0__SCAN_IN;
  assign n11493 = ~n11492 | ~n11836;
  assign n11495 = ~n11494 | ~n11493;
  assign n11497 = ~n11496 & ~n11495;
  assign n11501 = ~n11497 & ~n9044;
  assign n11499 = ~P1_ADDR_REG_0__SCAN_IN | ~n14842;
  assign n11498 = ~P1_REG3_REG_0__SCAN_IN | ~P1_U3084;
  assign n11500 = ~n11499 | ~n11498;
  assign n11506 = ~n11501 & ~n11500;
  assign n11503 = ~n14325 | ~P1_REG2_REG_0__SCAN_IN;
  assign n11502 = ~n14333 | ~P1_REG1_REG_0__SCAN_IN;
  assign n11504 = ~n11503 | ~n11502;
  assign n11505 = ~n11504 | ~n9044;
  assign P1_U3241 = ~n11506 | ~n11505;
  assign n11510 = ~n11508 | ~n11507;
  assign n11509 = ~n11517 | ~P1_REG2_REG_6__SCAN_IN;
  assign n11511 = ~n11614 ^ P1_REG2_REG_7__SCAN_IN;
  assign n11514 = ~n11512 & ~n11511;
  assign n11513 = ~n11691 | ~n14325;
  assign n11529 = ~n11514 & ~n11513;
  assign n11519 = ~n11516 & ~n11515;
  assign n11518 = ~n11517 & ~P1_REG1_REG_6__SCAN_IN;
  assign n11521 = ~n11519 & ~n11518;
  assign n11520 = ~n11614 ^ P1_REG1_REG_7__SCAN_IN;
  assign n11523 = ~n11521 & ~n11520;
  assign n11522 = ~n14333 | ~n11683;
  assign n11525 = ~n11523 & ~n11522;
  assign n12755 = ~P1_STATE_REG_SCAN_IN & ~n11524;
  assign n11527 = ~n11525 & ~n12755;
  assign n11689 = ~n11614;
  assign n11526 = ~n14837 | ~n11689;
  assign n11528 = ~n11527 | ~n11526;
  assign n11531 = ~n11529 & ~n11528;
  assign n11530 = ~P1_ADDR_REG_7__SCAN_IN | ~n14842;
  assign P1_U3248 = ~n11531 | ~n11530;
  assign n11534 = ~n11537 & ~n14384;
  assign n11533 = ~n11532 & ~P1_U3084;
  assign n11536 = ~n11534 & ~n11533;
  assign n11535 = ~n14388 | ~P2_DATAO_REG_6__SCAN_IN;
  assign P1_U3347 = ~n11536 | ~n11535;
  assign n11540 = ~n11537 & ~n14094;
  assign n11538 = ~n12273;
  assign n11539 = ~n11538 & ~P2_U3152;
  assign n11542 = ~n11540 & ~n11539;
  assign n11541 = ~n14577 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P2_U3352 = ~n11542 | ~n11541;
  assign ADD_1071_U48 = ~n11544 ^ n11543;
  assign n11547 = ~n11545 | ~n11059;
  assign n11546 = ~n12236 | ~P2_STATE_REG_SCAN_IN;
  assign n11549 = n11547 & n11546;
  assign n11548 = ~n14577 | ~P1_DATAO_REG_2__SCAN_IN;
  assign P2_U3356 = ~n11549 | ~n11548;
  assign n11554 = ~n11551 & ~n11550;
  assign n11553 = ~n11552 | ~n14325;
  assign n11566 = ~n11554 & ~n11553;
  assign n11559 = ~n11556 & ~n11555;
  assign n11558 = ~n14333 | ~n11557;
  assign n11561 = ~n11559 & ~n11558;
  assign n11560 = ~P1_REG3_REG_5__SCAN_IN;
  assign n12826 = ~P1_STATE_REG_SCAN_IN & ~n11560;
  assign n11564 = ~n11561 & ~n12826;
  assign n11563 = ~n14837 | ~n11562;
  assign n11565 = ~n11564 | ~n11563;
  assign n11568 = ~n11566 & ~n11565;
  assign n11567 = ~P1_ADDR_REG_5__SCAN_IN | ~n14842;
  assign P1_U3246 = ~n11568 | ~n11567;
  assign n11571 = ~n11570 & ~n11569;
  assign n11573 = ~n11571 & ~n14833;
  assign n11575 = ~n11573 | ~n11572;
  assign n11574 = ~P1_REG3_REG_1__SCAN_IN | ~P1_U3084;
  assign n11583 = ~n11575 | ~n11574;
  assign n11581 = ~P1_ADDR_REG_1__SCAN_IN | ~n14842;
  assign n11577 = ~n11838 & ~n11576;
  assign n11579 = ~n14825 & ~n11577;
  assign n11580 = ~n11579 | ~n11578;
  assign n11582 = ~n11581 | ~n11580;
  assign n11586 = ~n11583 & ~n11582;
  assign n11585 = ~n14837 | ~n11584;
  assign P1_U3242 = ~n11586 | ~n11585;
  assign n11588 = ~n12763 | ~P1_U4006;
  assign n11587 = ~n12117 | ~P1_DATAO_REG_5__SCAN_IN;
  assign P1_U3560 = ~n11588 | ~n11587;
  assign n11590 = ~n13474 | ~P1_U4006;
  assign n11589 = ~n12117 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P1_U3564 = ~n11590 | ~n11589;
  assign n11592 = ~n13228 | ~P1_U4006;
  assign n11591 = ~n12117 | ~P1_DATAO_REG_8__SCAN_IN;
  assign P1_U3563 = ~n11592 | ~n11591;
  assign n11594 = ~n13104 | ~P1_U4006;
  assign n11593 = ~n12117 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P1_U3562 = ~n11594 | ~n11593;
  assign n11596 = ~P1_DATAO_REG_22__SCAN_IN | ~n12117;
  assign n11595 = ~P1_U4006 | ~n15512;
  assign P1_U3577 = ~n11596 | ~n11595;
  assign n11598 = ~n16693 | ~P1_U4006;
  assign n11597 = ~n12117 | ~P1_DATAO_REG_16__SCAN_IN;
  assign P1_U3571 = ~n11598 | ~n11597;
  assign n11600 = ~n16666 | ~P1_U4006;
  assign n11599 = ~n12117 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P1_U3568 = ~n11600 | ~n11599;
  assign n11602 = ~n13855 | ~P1_U4006;
  assign n11601 = ~n12117 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P1_U3567 = ~n11602 | ~n11601;
  assign n11604 = ~n16678 | ~P1_U4006;
  assign n11603 = ~n12117 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P1_U3569 = ~n11604 | ~n11603;
  assign n11606 = ~n14527 | ~P1_U4006;
  assign n11605 = ~n12117 | ~P1_DATAO_REG_15__SCAN_IN;
  assign P1_U3570 = ~n11606 | ~n11605;
  assign n11608 = ~n12495 | ~P1_U4006;
  assign n11607 = ~n12117 | ~P1_DATAO_REG_4__SCAN_IN;
  assign P1_U3559 = ~n11608 | ~n11607;
  assign n11610 = ~n16595 | ~P1_U4006;
  assign n11609 = ~n12117 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P1_U3561 = ~n11610 | ~n11609;
  assign P2_U3302 = P2_D_REG_26__SCAN_IN & n11613;
  assign P2_U3326 = P2_D_REG_2__SCAN_IN & n11613;
  assign P2_U3324 = P2_D_REG_4__SCAN_IN & n11613;
  assign P2_U3300 = P2_D_REG_28__SCAN_IN & n11613;
  assign P2_U3303 = P2_D_REG_25__SCAN_IN & n11613;
  assign P2_U3321 = P2_D_REG_7__SCAN_IN & n11613;
  assign P2_U3301 = P2_D_REG_27__SCAN_IN & n11613;
  assign P2_U3297 = P2_D_REG_31__SCAN_IN & n11613;
  assign P2_U3304 = P2_D_REG_24__SCAN_IN & n11613;
  assign P2_U3305 = P2_D_REG_23__SCAN_IN & n11613;
  assign P2_U3308 = P2_D_REG_20__SCAN_IN & n11613;
  assign P2_U3307 = P2_D_REG_21__SCAN_IN & n11613;
  assign P2_U3306 = P2_D_REG_22__SCAN_IN & n11613;
  assign P2_U3309 = P2_D_REG_19__SCAN_IN & n11613;
  assign P2_U3319 = P2_D_REG_9__SCAN_IN & n11613;
  assign P2_U3325 = P2_D_REG_3__SCAN_IN & n11613;
  assign P2_U3317 = P2_D_REG_11__SCAN_IN & n11613;
  assign P2_U3316 = P2_D_REG_12__SCAN_IN & n11613;
  assign P2_U3315 = P2_D_REG_13__SCAN_IN & n11613;
  assign P2_U3299 = P2_D_REG_29__SCAN_IN & n11613;
  assign P2_U3298 = P2_D_REG_30__SCAN_IN & n11613;
  assign P2_U3312 = P2_D_REG_16__SCAN_IN & n11613;
  assign P2_U3320 = P2_D_REG_8__SCAN_IN & n11613;
  assign P2_U3311 = P2_D_REG_17__SCAN_IN & n11613;
  assign P2_U3318 = P2_D_REG_10__SCAN_IN & n11613;
  assign P2_U3313 = P2_D_REG_15__SCAN_IN & n11613;
  assign P2_U3323 = P2_D_REG_5__SCAN_IN & n11613;
  assign P2_U3314 = P2_D_REG_14__SCAN_IN & n11613;
  assign P2_U3310 = P2_D_REG_18__SCAN_IN & n11613;
  assign P2_U3322 = P2_D_REG_6__SCAN_IN & n11613;
  assign n11616 = ~n11626 & ~n14384;
  assign n11615 = ~n11614 & ~P1_U3084;
  assign n11618 = ~n11616 & ~n11615;
  assign n11617 = ~n14388 | ~P2_DATAO_REG_7__SCAN_IN;
  assign P1_U3346 = ~n11618 | ~n11617;
  assign n11625 = ~P1_DATAO_REG_31__SCAN_IN | ~n12117;
  assign n11620 = ~n11671 | ~P1_REG0_REG_31__SCAN_IN;
  assign n11619 = ~n9544 | ~P1_REG2_REG_31__SCAN_IN;
  assign n11623 = ~n11620 | ~n11619;
  assign n11621 = ~P1_REG1_REG_31__SCAN_IN;
  assign n11622 = ~n11675 & ~n11621;
  assign n11624 = n12117 | n16837;
  assign P1_U3586 = ~n11625 | ~n11624;
  assign n11628 = ~n11626 & ~n14094;
  assign n11927 = ~n12070;
  assign n11627 = ~n11927 & ~P2_U3152;
  assign n11630 = ~n11628 & ~n11627;
  assign n11629 = ~n14577 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P2_U3351 = ~n11630 | ~n11629;
  assign n12644 = ~P2_REG3_REG_5__SCAN_IN | ~P2_U3152;
  assign n11633 = ~n11631 | ~n13709;
  assign n11634 = ~n11633 | ~n11632;
  assign n14864 = ~P2_U3152 & ~n11646;
  assign n11636 = ~n14864 | ~P2_ADDR_REG_5__SCAN_IN;
  assign n11652 = ~n12644 | ~n11636;
  assign n12187 = ~P2_REG1_REG_0__SCAN_IN;
  assign n12247 = ~n10261 & ~n12187;
  assign n12246 = ~n11653 ^ P2_REG1_REG_1__SCAN_IN;
  assign n12249 = ~n12247 | ~n12246;
  assign n12255 = ~n11653;
  assign n11637 = ~n12255 | ~P2_REG1_REG_1__SCAN_IN;
  assign n12223 = ~n12249 | ~n11637;
  assign n12222 = ~n11655 ^ P2_REG1_REG_2__SCAN_IN;
  assign n12225 = ~n12223 | ~n12222;
  assign n11638 = ~n12236 | ~P2_REG1_REG_2__SCAN_IN;
  assign n12204 = ~n12225 | ~n11638;
  assign n12203 = ~n11657 ^ P2_REG1_REG_3__SCAN_IN;
  assign n12206 = ~n12204 | ~n12203;
  assign n12217 = ~n11657;
  assign n11639 = ~n12217 | ~P2_REG1_REG_3__SCAN_IN;
  assign n12032 = ~n12206 | ~n11639;
  assign n12031 = n11659 ^ P2_REG1_REG_4__SCAN_IN;
  assign n11641 = ~n12032 & ~n12031;
  assign n12038 = ~n11659;
  assign n11640 = ~n12038 & ~P2_REG1_REG_4__SCAN_IN;
  assign n11643 = ~n11641 & ~n11640;
  assign n11642 = n11935 ^ P2_REG1_REG_5__SCAN_IN;
  assign n11924 = ~n11643 | ~n11642;
  assign n11645 = ~n11924;
  assign n11644 = ~n11643 & ~n11642;
  assign n11648 = ~n11645 & ~n11644;
  assign n11647 = ~n11662 | ~n16487;
  assign n11932 = ~n11664 & ~n11647;
  assign n11650 = ~n11648 | ~n11932;
  assign n14887 = ~n11664 & ~n11662;
  assign n11649 = ~n14887 | ~n11935;
  assign n11651 = ~n11650 | ~n11649;
  assign n11670 = ~n11652 & ~n11651;
  assign n12186 = ~P2_REG2_REG_0__SCAN_IN;
  assign n12240 = ~n10261 & ~n12186;
  assign n12239 = ~n11653 ^ P2_REG2_REG_1__SCAN_IN;
  assign n12242 = ~n12240 | ~n12239;
  assign n11654 = ~n12255 | ~P2_REG2_REG_1__SCAN_IN;
  assign n12228 = ~n12242 | ~n11654;
  assign n12227 = ~n11655 ^ P2_REG2_REG_2__SCAN_IN;
  assign n12230 = ~n12228 | ~n12227;
  assign n11656 = ~n12236 | ~P2_REG2_REG_2__SCAN_IN;
  assign n12209 = ~n12230 | ~n11656;
  assign n12208 = ~n11657 ^ P2_REG2_REG_3__SCAN_IN;
  assign n12211 = ~n12209 | ~n12208;
  assign n11658 = ~n12217 | ~P2_REG2_REG_3__SCAN_IN;
  assign n12029 = ~n12211 | ~n11658;
  assign n12028 = n11659 ^ P2_REG2_REG_4__SCAN_IN;
  assign n11661 = ~n12029 & ~n12028;
  assign n11660 = ~n12038 & ~P2_REG2_REG_4__SCAN_IN;
  assign n11667 = ~n11661 & ~n11660;
  assign n11666 = n11935 ^ P2_REG2_REG_5__SCAN_IN;
  assign n11665 = ~n11667 & ~n11666;
  assign n15261 = ~n16487;
  assign n11663 = ~n11662 | ~n15261;
  assign n14882 = ~n11664 & ~n11663;
  assign n12924 = ~n14882;
  assign n11668 = ~n11665 & ~n12924;
  assign n11937 = ~n11667 | ~n11666;
  assign n11669 = ~n11668 | ~n11937;
  assign P2_U3250 = ~n11670 | ~n11669;
  assign n11679 = ~P1_DATAO_REG_30__SCAN_IN | ~n12117;
  assign n11673 = ~n11671 | ~P1_REG0_REG_30__SCAN_IN;
  assign n11672 = ~n9544 | ~P1_REG2_REG_30__SCAN_IN;
  assign n11677 = ~n11673 | ~n11672;
  assign n11674 = ~P1_REG1_REG_30__SCAN_IN;
  assign n11676 = ~n11675 & ~n11674;
  assign n11678 = n12117 | n17062;
  assign P1_U3585 = ~n11679 | ~n11678;
  assign n11681 = ~P1_DATAO_REG_18__SCAN_IN | ~n12117;
  assign n11680 = ~P1_U4006 | ~n14605;
  assign P1_U3573 = ~n11681 | ~n11680;
  assign n12951 = ~P1_REG3_REG_8__SCAN_IN | ~P1_U3084;
  assign n11682 = ~n11689 | ~P1_REG1_REG_7__SCAN_IN;
  assign n11685 = ~n11693 ^ P1_REG1_REG_8__SCAN_IN;
  assign n11684 = ~n11686 & ~n11685;
  assign n11687 = ~n11684 & ~n14833;
  assign n11688 = ~n11687 | ~n11719;
  assign n11703 = ~n12951 | ~n11688;
  assign n11701 = ~n14842 | ~P1_ADDR_REG_8__SCAN_IN;
  assign n11690 = ~n11689 | ~P1_REG2_REG_7__SCAN_IN;
  assign n11734 = ~n11693;
  assign n11694 = ~n11734 | ~P1_REG2_REG_8__SCAN_IN;
  assign n11712 = ~n11693 | ~n11692;
  assign n11695 = ~n11694 | ~n11712;
  assign n11698 = ~n11714;
  assign n11697 = ~n11696 | ~n11695;
  assign n11699 = ~n11698 | ~n11697;
  assign n11700 = ~n11699 | ~n14325;
  assign n11702 = ~n11701 | ~n11700;
  assign n11705 = ~n11703 & ~n11702;
  assign n11704 = ~n14837 | ~n11734;
  assign P1_U3249 = ~n11705 | ~n11704;
  assign n11707 = ~P1_DATAO_REG_20__SCAN_IN | ~n12117;
  assign n11706 = ~P1_U4006 | ~n15088;
  assign P1_U3575 = ~n11707 | ~n11706;
  assign n11709 = ~P1_DATAO_REG_21__SCAN_IN | ~n12117;
  assign n11708 = ~P1_U4006 | ~n16739;
  assign P1_U3576 = ~n11709 | ~n11708;
  assign n11711 = ~P1_DATAO_REG_23__SCAN_IN | ~n12117;
  assign n11710 = ~P1_U4006 | ~n15159;
  assign P1_U3578 = ~n11711 | ~n11710;
  assign n11713 = ~n11712;
  assign n11779 = ~n11721;
  assign n11716 = ~n11779 | ~P1_REG2_REG_9__SCAN_IN;
  assign n11715 = ~P1_REG2_REG_9__SCAN_IN;
  assign n11756 = ~n11721 | ~n11715;
  assign n11754 = ~n11716 | ~n11756;
  assign n11717 = n11755 ^ n11754;
  assign n11729 = ~n11717 & ~n14825;
  assign n11718 = ~n11734 | ~P1_REG1_REG_8__SCAN_IN;
  assign n11722 = ~n11779 | ~P1_REG1_REG_9__SCAN_IN;
  assign n11720 = ~P1_REG1_REG_9__SCAN_IN;
  assign n11746 = ~n11721 | ~n11720;
  assign n11744 = ~n11722 | ~n11746;
  assign n11723 = n11745 ^ n11744;
  assign n11725 = ~n11723 & ~n14833;
  assign n13276 = ~P1_STATE_REG_SCAN_IN & ~n11724;
  assign n11727 = ~n11725 & ~n13276;
  assign n11726 = ~n14837 | ~n11779;
  assign n11728 = ~n11727 | ~n11726;
  assign n11731 = ~n11729 & ~n11728;
  assign n11730 = ~P1_ADDR_REG_9__SCAN_IN | ~n14842;
  assign P1_U3250 = ~n11731 | ~n11730;
  assign ADD_1071_U47 = ~n11733 ^ n11732;
  assign n11736 = ~n11739 | ~n14582;
  assign n11735 = ~n11734 | ~P1_STATE_REG_SCAN_IN;
  assign n11738 = n11736 & n11735;
  assign n11737 = ~n14388 | ~P2_DATAO_REG_8__SCAN_IN;
  assign P1_U3345 = ~n11738 | ~n11737;
  assign n11741 = ~n11739 | ~n11059;
  assign n11740 = ~n12135 | ~P2_STATE_REG_SCAN_IN;
  assign n11743 = n11741 & n11740;
  assign n11742 = ~n14577 | ~P1_DATAO_REG_8__SCAN_IN;
  assign P2_U3350 = ~n11743 | ~n11742;
  assign n13479 = ~P1_REG3_REG_10__SCAN_IN | ~P1_U3084;
  assign n11747 = ~n11746;
  assign n11750 = ~P1_REG1_REG_10__SCAN_IN ^ n11759;
  assign n11749 = ~n11751 & ~n11750;
  assign n11752 = ~n11749 & ~n14833;
  assign n11753 = ~n11752 | ~n11975;
  assign n11767 = ~n13479 | ~n11753;
  assign n11765 = ~n14837 | ~n11974;
  assign n11757 = ~n11756;
  assign n11761 = ~P1_REG2_REG_10__SCAN_IN ^ n11759;
  assign n11760 = ~n11762 & ~n11761;
  assign n11763 = ~n11760 & ~n14825;
  assign n11764 = ~n11763 | ~n11971;
  assign n11766 = ~n11765 | ~n11764;
  assign n11769 = ~n11767 & ~n11766;
  assign n11768 = ~n14842 | ~P1_ADDR_REG_10__SCAN_IN;
  assign P1_U3251 = ~n11769 | ~n11768;
  assign n11771 = ~P1_DATAO_REG_24__SCAN_IN | ~n12117;
  assign n11770 = ~P1_U4006 | ~n15697;
  assign P1_U3579 = ~n11771 | ~n11770;
  assign P2_U3151 = ~n14864 & ~P2_U3966;
  assign n11773 = ~P1_DATAO_REG_26__SCAN_IN | ~n12117;
  assign n11772 = ~P1_U4006 | ~n16787;
  assign P1_U3581 = ~n11773 | ~n11772;
  assign n11775 = ~n11778 | ~n11059;
  assign n11774 = ~n11962 | ~P2_STATE_REG_SCAN_IN;
  assign n11777 = n11775 & n11774;
  assign n11776 = ~n14577 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P2_U3349 = ~n11777 | ~n11776;
  assign n11781 = ~n11778 | ~n14582;
  assign n11780 = ~n11779 | ~P1_STATE_REG_SCAN_IN;
  assign n11783 = n11781 & n11780;
  assign n11782 = ~n14388 | ~P2_DATAO_REG_9__SCAN_IN;
  assign P1_U3344 = ~n11783 | ~n11782;
  assign n11785 = ~P1_DATAO_REG_25__SCAN_IN | ~n12117;
  assign n11784 = ~P1_U4006 | ~n16781;
  assign P1_U3580 = ~n11785 | ~n11784;
  assign n11787 = ~P2_DATAO_REG_22__SCAN_IN | ~n13390;
  assign n11786 = ~P2_U3966 | ~n16334;
  assign P2_U3574 = ~n11787 | ~n11786;
  assign n11790 = ~P2_DATAO_REG_18__SCAN_IN | ~n13390;
  assign n11789 = ~P2_U3966 | ~n11788;
  assign P2_U3570 = ~n11790 | ~n11789;
  assign n11796 = ~P2_DATAO_REG_30__SCAN_IN | ~n13390;
  assign n11792 = ~n11807 | ~P2_REG1_REG_30__SCAN_IN;
  assign n11791 = ~n11804 | ~P2_REG2_REG_30__SCAN_IN;
  assign n11794 = n11792 & n11791;
  assign n11793 = ~n11803 | ~P2_REG0_REG_30__SCAN_IN;
  assign n11795 = ~P2_U3966 | ~n16452;
  assign P2_U3582 = ~n11796 | ~n11795;
  assign n11798 = ~P2_DATAO_REG_21__SCAN_IN | ~n13390;
  assign n11797 = ~P2_U3966 | ~n16322;
  assign P2_U3573 = ~n11798 | ~n11797;
  assign n11800 = ~P2_DATAO_REG_19__SCAN_IN | ~n13390;
  assign n11799 = ~P2_U3966 | ~n14506;
  assign P2_U3571 = ~n11800 | ~n11799;
  assign n11802 = ~P2_DATAO_REG_20__SCAN_IN | ~n13390;
  assign n11801 = ~P2_U3966 | ~n16299;
  assign P2_U3572 = ~n11802 | ~n11801;
  assign n11811 = ~P2_DATAO_REG_31__SCAN_IN | ~n13390;
  assign n11806 = ~n9033 | ~P2_REG0_REG_31__SCAN_IN;
  assign n11805 = ~n11804 | ~P2_REG2_REG_31__SCAN_IN;
  assign n11809 = n11806 & n11805;
  assign n11808 = ~n11807 | ~P2_REG1_REG_31__SCAN_IN;
  assign n11810 = ~P2_U3966 | ~n15967;
  assign P2_U3583 = ~n11811 | ~n11810;
  assign n11815 = ~n11813 & ~n11812;
  assign ADD_1071_U63 = n11815 ^ n11814;
  assign n11817 = ~n16248 | ~P2_U3966;
  assign n11816 = ~P2_DATAO_REG_14__SCAN_IN | ~n13390;
  assign P2_U3566 = ~n11817 | ~n11816;
  assign n11819 = ~n11822 | ~n14582;
  assign n11818 = ~n12105 | ~P1_STATE_REG_SCAN_IN;
  assign n11821 = n11819 & n11818;
  assign n11820 = ~n14388 | ~P2_DATAO_REG_11__SCAN_IN;
  assign P1_U3342 = ~n11821 | ~n11820;
  assign n11824 = ~n11822 | ~n11059;
  assign n11823 = ~n12306 | ~P2_STATE_REG_SCAN_IN;
  assign n11826 = n11824 & n11823;
  assign n11825 = ~n14577 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P2_U3347 = ~n11826 | ~n11825;
  assign n11828 = ~n11831 | ~n11059;
  assign n11827 = ~n12088 | ~P2_STATE_REG_SCAN_IN;
  assign n11830 = n11828 & n11827;
  assign n11829 = ~n14577 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P2_U3348 = ~n11830 | ~n11829;
  assign n11833 = ~n11831 | ~n14582;
  assign n11832 = ~n11974 | ~P1_STATE_REG_SCAN_IN;
  assign n11835 = n11833 & n11832;
  assign n11834 = ~n14388 | ~P2_DATAO_REG_10__SCAN_IN;
  assign P1_U3343 = ~n11835 | ~n11834;
  assign n11837 = n11846 | n11836;
  assign n11840 = ~n9044 | ~n11837;
  assign n11839 = ~n11838 & ~n11845;
  assign n11842 = ~n11840 | ~n11839;
  assign n11841 = ~n11846 | ~P1_IR_REG_0__SCAN_IN;
  assign n11849 = ~n11842 | ~n11841;
  assign n12630 = n11844 ^ n11843;
  assign n17087 = ~n11845;
  assign n11847 = ~n11846 & ~n17087;
  assign n11848 = n12630 & n11847;
  assign n11850 = ~n11849 & ~n11848;
  assign n11918 = ~n12117 & ~n11850;
  assign n11855 = ~n11852 & ~n11851;
  assign n11854 = ~n14333 | ~n11853;
  assign n11863 = ~n11855 & ~n11854;
  assign n11858 = n11857 ^ n11856;
  assign n11861 = ~n14325 | ~n11858;
  assign n11860 = ~n14837 | ~n11859;
  assign n11862 = ~n11861 | ~n11860;
  assign n11865 = ~n11863 & ~n11862;
  assign n11864 = ~P1_REG3_REG_2__SCAN_IN | ~P1_U3084;
  assign n11866 = ~n11865 | ~n11864;
  assign n11868 = ~n11918 & ~n11866;
  assign n11867 = ~P1_ADDR_REG_2__SCAN_IN | ~n14842;
  assign P1_U3243 = ~n11868 | ~n11867;
  assign n11870 = ~n12383 | ~P2_U3966;
  assign n11869 = ~P2_DATAO_REG_0__SCAN_IN | ~n13390;
  assign P2_U3552 = ~n11870 | ~n11869;
  assign n11872 = ~n13988 | ~P2_U3966;
  assign n11871 = ~P2_DATAO_REG_13__SCAN_IN | ~n13390;
  assign P2_U3565 = ~n11872 | ~n11871;
  assign n11874 = ~n16230 | ~P2_U3966;
  assign n11873 = ~P2_DATAO_REG_12__SCAN_IN | ~n13390;
  assign P2_U3564 = ~n11874 | ~n11873;
  assign n11876 = ~n16189 | ~P2_U3966;
  assign n11875 = ~P2_DATAO_REG_11__SCAN_IN | ~n13390;
  assign P2_U3563 = ~n11876 | ~n11875;
  assign n11878 = ~n16195 | ~P2_U3966;
  assign n11877 = ~P2_DATAO_REG_10__SCAN_IN | ~n13390;
  assign P2_U3562 = ~n11878 | ~n11877;
  assign n11880 = ~n16177 | ~P2_U3966;
  assign n11879 = ~P2_DATAO_REG_9__SCAN_IN | ~n13390;
  assign P2_U3561 = ~n11880 | ~n11879;
  assign n11882 = ~n16161 | ~P2_U3966;
  assign n11881 = ~P2_DATAO_REG_8__SCAN_IN | ~n13390;
  assign P2_U3560 = ~n11882 | ~n11881;
  assign n11884 = ~n13288 | ~P2_U3966;
  assign n11883 = ~P2_DATAO_REG_7__SCAN_IN | ~n13390;
  assign P2_U3559 = ~n11884 | ~n11883;
  assign n11886 = ~n16073 | ~P2_U3966;
  assign n11885 = ~P2_DATAO_REG_2__SCAN_IN | ~n13390;
  assign P2_U3554 = ~n11886 | ~n11885;
  assign n11887 = ~n16124;
  assign n11889 = ~n11887 | ~P2_U3966;
  assign n11888 = ~P2_DATAO_REG_3__SCAN_IN | ~n13390;
  assign P2_U3555 = ~n11889 | ~n11888;
  assign n11891 = ~n12388 | ~P2_U3966;
  assign n11890 = ~P2_DATAO_REG_1__SCAN_IN | ~n13390;
  assign P2_U3553 = ~n11891 | ~n11890;
  assign n11893 = ~n16277 | ~P2_U3966;
  assign n11892 = ~P2_DATAO_REG_16__SCAN_IN | ~n13390;
  assign P2_U3568 = ~n11893 | ~n11892;
  assign n11895 = ~n13251 | ~P2_U3966;
  assign n11894 = ~P2_DATAO_REG_6__SCAN_IN | ~n13390;
  assign P2_U3558 = ~n11895 | ~n11894;
  assign n11897 = ~n16116 | ~P2_U3966;
  assign n11896 = ~P2_DATAO_REG_4__SCAN_IN | ~n13390;
  assign P2_U3556 = ~n11897 | ~n11896;
  assign n11899 = ~n13014 | ~P2_U3966;
  assign n11898 = ~P2_DATAO_REG_5__SCAN_IN | ~n13390;
  assign P2_U3557 = ~n11899 | ~n11898;
  assign n11901 = ~n16051 | ~P2_U3966;
  assign n11900 = ~P2_DATAO_REG_17__SCAN_IN | ~n13390;
  assign P2_U3569 = ~n11901 | ~n11900;
  assign n11903 = ~n16265 | ~P2_U3966;
  assign n11902 = ~P2_DATAO_REG_15__SCAN_IN | ~n13390;
  assign P2_U3567 = ~n11903 | ~n11902;
  assign n11906 = n11905 ^ n11904;
  assign n11909 = ~n11906 | ~n14325;
  assign n11908 = ~n14837 | ~n11907;
  assign n11916 = ~n11909 | ~n11908;
  assign n11914 = ~n11911 & ~n11910;
  assign n11913 = ~n14333 | ~n11912;
  assign n11915 = ~n11914 & ~n11913;
  assign n11917 = ~n11916 & ~n11915;
  assign n12672 = ~P1_REG3_REG_4__SCAN_IN | ~P1_U3084;
  assign n11919 = ~n11917 | ~n12672;
  assign n11921 = ~n11919 & ~n11918;
  assign n11920 = ~n14842 | ~P1_ADDR_REG_4__SCAN_IN;
  assign P1_U3245 = ~n11921 | ~n11920;
  assign n13550 = ~P2_REG3_REG_9__SCAN_IN | ~P2_U3152;
  assign n11922 = ~n14864 | ~P2_ADDR_REG_9__SCAN_IN;
  assign n11949 = ~n13550 | ~n11922;
  assign n11931 = ~P2_REG1_REG_8__SCAN_IN | ~n12135;
  assign n12126 = ~P2_REG1_REG_8__SCAN_IN ^ n11934;
  assign n11923 = ~n11935 | ~P2_REG1_REG_5__SCAN_IN;
  assign n12260 = ~n11924 | ~n11923;
  assign n12259 = n12273 ^ P2_REG1_REG_6__SCAN_IN;
  assign n12262 = ~n12260 | ~n12259;
  assign n11925 = ~n12273 | ~P2_REG1_REG_6__SCAN_IN;
  assign n12056 = ~n12262 | ~n11925;
  assign n11929 = ~n11927 | ~n11926;
  assign n11928 = ~n12070 | ~P2_REG1_REG_7__SCAN_IN;
  assign n12055 = ~n11929 | ~n11928;
  assign n12054 = ~n12056 & ~n12055;
  assign n11930 = ~n11929;
  assign n12127 = ~n12054 & ~n11930;
  assign n11953 = P2_REG1_REG_9__SCAN_IN ^ n11944;
  assign n11933 = ~n11954 ^ n11953;
  assign n11947 = ~n11933 | ~n11932;
  assign n11943 = ~P2_REG2_REG_8__SCAN_IN | ~n12135;
  assign n12121 = ~P2_REG2_REG_8__SCAN_IN ^ n11934;
  assign n11936 = ~n11935 | ~P2_REG2_REG_5__SCAN_IN;
  assign n12265 = ~n11937 | ~n11936;
  assign n12264 = n12273 ^ P2_REG2_REG_6__SCAN_IN;
  assign n12267 = ~n12265 | ~n12264;
  assign n11938 = ~n12273 | ~P2_REG2_REG_6__SCAN_IN;
  assign n12062 = ~n12267 | ~n11938;
  assign n11940 = ~n12062;
  assign n11939 = n12070 & P2_REG2_REG_7__SCAN_IN;
  assign n11941 = ~n12070 & ~P2_REG2_REG_7__SCAN_IN;
  assign n12060 = ~n11939 & ~n11941;
  assign n11942 = ~n12064;
  assign n11963 = P2_REG2_REG_9__SCAN_IN ^ n11944;
  assign n11945 = ~n11964 ^ n11963;
  assign n11946 = ~n11945 | ~n14882;
  assign n11948 = ~n11947 | ~n11946;
  assign n11951 = ~n11949 & ~n11948;
  assign n11950 = ~n14887 | ~n11962;
  assign P2_U3254 = ~n11951 | ~n11950;
  assign n13513 = ~P2_REG3_REG_10__SCAN_IN | ~P2_U3152;
  assign n11952 = ~n14864 | ~P2_ADDR_REG_10__SCAN_IN;
  assign n11961 = ~n13513 | ~n11952;
  assign n11959 = ~n14887 | ~n12088;
  assign n11956 = ~P2_REG1_REG_9__SCAN_IN & ~n11962;
  assign n11955 = ~n11954 & ~n11953;
  assign n12089 = P2_REG1_REG_10__SCAN_IN ^ n11967;
  assign n11957 = ~n12090 ^ n12089;
  assign n11958 = ~n11957 | ~n11932;
  assign n11960 = ~n11959 | ~n11958;
  assign n11970 = ~n11961 & ~n11960;
  assign n11966 = ~P2_REG2_REG_9__SCAN_IN & ~n11962;
  assign n12082 = P2_REG2_REG_10__SCAN_IN ^ n11967;
  assign n11968 = ~n12083 ^ n12082;
  assign n11969 = ~n14882 | ~n11968;
  assign P2_U3255 = ~n11970 | ~n11969;
  assign n12107 = ~n12105 ^ P1_REG2_REG_11__SCAN_IN;
  assign n11972 = ~n11974 | ~P1_REG2_REG_10__SCAN_IN;
  assign n11973 = n12107 ^ n12106;
  assign n11986 = ~n11973 & ~n14825;
  assign n11978 = n12105 ^ P1_REG1_REG_11__SCAN_IN;
  assign n11976 = ~n11974 | ~P1_REG1_REG_10__SCAN_IN;
  assign n11980 = ~n11978 & ~n11977;
  assign n11979 = ~n14333 | ~n12101;
  assign n11982 = ~n11980 & ~n11979;
  assign n13570 = ~P1_STATE_REG_SCAN_IN & ~n11981;
  assign n11984 = ~n11982 & ~n13570;
  assign n11983 = ~n14837 | ~n12105;
  assign n11985 = ~n11984 | ~n11983;
  assign n11988 = ~n11986 & ~n11985;
  assign n11987 = ~P1_ADDR_REG_11__SCAN_IN | ~n14842;
  assign P1_U3252 = ~n11988 | ~n11987;
  assign n11990 = ~P1_DATAO_REG_27__SCAN_IN | ~n12117;
  assign n11989 = ~P1_U4006 | ~n16853;
  assign P1_U3582 = ~n11990 | ~n11989;
  assign n11992 = ~n11995 | ~n14582;
  assign n11991 = ~n12477 | ~P1_STATE_REG_SCAN_IN;
  assign n11994 = n11992 & n11991;
  assign n11993 = ~n14388 | ~P2_DATAO_REG_12__SCAN_IN;
  assign P1_U3341 = ~n11994 | ~n11993;
  assign n11997 = ~n11995 | ~n11059;
  assign n11996 = ~n12581 | ~P2_STATE_REG_SCAN_IN;
  assign n11999 = n11997 & n11996;
  assign n11998 = ~n14577 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P2_U3346 = ~n11999 | ~n11998;
  assign n12003 = ~n12001 & ~n12000;
  assign ADD_1071_U62 = n12003 ^ n12002;
  assign n12019 = ~P2_REG0_REG_0__SCAN_IN | ~n16511;
  assign n12010 = ~n12383 & ~n10645;
  assign n15970 = ~n12010 & ~n12345;
  assign n12011 = ~n14769 | ~n15547;
  assign n12013 = ~n15970 | ~n12011;
  assign n12012 = ~n12388 | ~n15549;
  assign n13093 = n12013 & n12012;
  assign n13094 = ~n15970;
  assign n16498 = ~n16080 | ~n9039;
  assign n12016 = ~n13094 & ~n16498;
  assign n12015 = ~n16071 & ~n12014;
  assign n12017 = ~n12016 & ~n12015;
  assign n12022 = ~n13093 | ~n12017;
  assign n12018 = ~n16510 | ~n12022;
  assign P2_U3451 = ~n12019 | ~n12018;
  assign n12024 = ~P2_REG1_REG_0__SCAN_IN | ~n16516;
  assign n12023 = ~n16514 | ~n12022;
  assign P2_U3520 = ~n12024 | ~n12023;
  assign n12026 = ~P2_DATAO_REG_23__SCAN_IN | ~n13390;
  assign n12025 = ~P2_U3966 | ~n16347;
  assign P2_U3575 = ~n12026 | ~n12025;
  assign n12613 = ~P2_REG3_REG_4__SCAN_IN | ~P2_U3152;
  assign n12027 = ~n14864 | ~P2_ADDR_REG_4__SCAN_IN;
  assign n12037 = ~n12613 | ~n12027;
  assign n12030 = ~n12029 ^ n12028;
  assign n12035 = ~n12030 | ~n14882;
  assign n12033 = ~n12032 ^ n12031;
  assign n12034 = ~n11932 | ~n12033;
  assign n12036 = ~n12035 | ~n12034;
  assign n12040 = ~n12037 & ~n12036;
  assign n12039 = ~n14887 | ~n12038;
  assign P2_U3249 = ~n12040 | ~n12039;
  assign n12052 = ~P1_DATAO_REG_29__SCAN_IN | ~n12117;
  assign n12045 = ~n12041 & ~n15765;
  assign n12042 = ~P1_REG0_REG_29__SCAN_IN;
  assign n12044 = ~n12043 & ~n12042;
  assign n12050 = ~n12045 & ~n12044;
  assign n12048 = ~n9037 | ~P1_REG2_REG_29__SCAN_IN;
  assign n12047 = ~n12046 | ~P1_REG1_REG_29__SCAN_IN;
  assign n12049 = n12048 & n12047;
  assign n12051 = ~P1_U4006 | ~n17131;
  assign P1_U3584 = ~n12052 | ~n12051;
  assign n13199 = ~P2_REG3_REG_7__SCAN_IN | ~P2_U3152;
  assign n12053 = ~n14864 | ~P2_ADDR_REG_7__SCAN_IN;
  assign n12069 = ~n13199 | ~n12053;
  assign n12058 = ~n12054;
  assign n12057 = ~n12056 | ~n12055;
  assign n12059 = ~n12058 | ~n12057;
  assign n12067 = ~n12059 | ~n11932;
  assign n12061 = ~n12060;
  assign n12063 = ~n12062 | ~n12061;
  assign n12065 = ~n12064 | ~n12063;
  assign n12066 = ~n12065 | ~n14882;
  assign n12068 = ~n12067 | ~n12066;
  assign n12072 = ~n12069 & ~n12068;
  assign n12071 = ~n14887 | ~n12070;
  assign P2_U3252 = ~n12072 | ~n12071;
  assign n12074 = ~n12077 | ~n14582;
  assign n12073 = ~n12983 | ~P1_STATE_REG_SCAN_IN;
  assign n12076 = n12074 & n12073;
  assign n12075 = ~n14388 | ~P2_DATAO_REG_13__SCAN_IN;
  assign P1_U3340 = ~n12076 | ~n12075;
  assign n12079 = ~n12077 | ~n11059;
  assign n12078 = ~n12919 | ~P2_STATE_REG_SCAN_IN;
  assign n12081 = n12079 & n12078;
  assign n12080 = ~n14577 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P2_U3345 = ~n12081 | ~n12080;
  assign n13640 = ~P2_REG3_REG_11__SCAN_IN | ~P2_U3152;
  assign n12085 = ~P2_REG2_REG_10__SCAN_IN & ~n12088;
  assign n12086 = ~n12308 ^ n12307;
  assign n12087 = ~n12086 | ~n14882;
  assign n12097 = ~n13640 | ~n12087;
  assign n12095 = ~n14864 | ~P2_ADDR_REG_11__SCAN_IN;
  assign n12092 = ~P2_REG1_REG_10__SCAN_IN & ~n12088;
  assign n12301 = ~P2_REG1_REG_11__SCAN_IN ^ n12306;
  assign n12093 = ~n12302 ^ n12301;
  assign n12094 = ~n12093 | ~n11932;
  assign n12096 = ~n12095 | ~n12094;
  assign n12099 = ~n12097 & ~n12096;
  assign n12098 = ~n14887 | ~n12306;
  assign P2_U3256 = ~n12099 | ~n12098;
  assign n13819 = ~P1_U3084 | ~P1_REG3_REG_12__SCAN_IN;
  assign n12100 = ~n14837 | ~n12477;
  assign n12114 = ~n13819 | ~n12100;
  assign n12471 = ~P1_REG1_REG_12__SCAN_IN & ~n12477;
  assign n12470 = P1_REG1_REG_12__SCAN_IN & n12477;
  assign n12103 = ~n12471 & ~n12470;
  assign n12102 = ~n12105 | ~P1_REG1_REG_11__SCAN_IN;
  assign n12104 = n12103 ^ n12469;
  assign n12112 = ~n14333 | ~n12104;
  assign n12109 = ~n12105 & ~P1_REG2_REG_11__SCAN_IN;
  assign n12478 = ~P1_REG2_REG_12__SCAN_IN ^ n12477;
  assign n12110 = ~n12479 ^ n12478;
  assign n12111 = ~n12110 | ~n14325;
  assign n12113 = ~n12112 | ~n12111;
  assign n12116 = ~n12114 & ~n12113;
  assign n12115 = ~n14842 | ~P1_ADDR_REG_12__SCAN_IN;
  assign P1_U3253 = ~n12116 | ~n12115;
  assign n12119 = ~P1_DATAO_REG_28__SCAN_IN | ~n12117;
  assign n12118 = ~P1_U4006 | ~n17112;
  assign P1_U3583 = ~n12119 | ~n12118;
  assign n13289 = ~P2_REG3_REG_8__SCAN_IN | ~P2_U3152;
  assign n12122 = ~n12121 & ~n12120;
  assign n12124 = ~n12122 & ~n12924;
  assign n12125 = ~n12124 | ~n12123;
  assign n12134 = ~n13289 | ~n12125;
  assign n12132 = ~P2_ADDR_REG_8__SCAN_IN | ~n14864;
  assign n12128 = ~n12127 & ~n12126;
  assign n12917 = ~n11932;
  assign n12130 = ~n12128 & ~n12917;
  assign n12131 = ~n12130 | ~n12129;
  assign n12133 = ~n12132 | ~n12131;
  assign n12137 = ~n12134 & ~n12133;
  assign n12136 = ~n14887 | ~n12135;
  assign P2_U3253 = ~n12137 | ~n12136;
  assign n12141 = ~n12139 & ~n12138;
  assign ADD_1071_U61 = n12141 ^ n12140;
  assign n12143 = ~n12146 | ~n14582;
  assign n12142 = ~n13458 | ~P1_STATE_REG_SCAN_IN;
  assign n12145 = n12143 & n12142;
  assign n12144 = ~n14388 | ~P2_DATAO_REG_14__SCAN_IN;
  assign P1_U3339 = ~n12145 | ~n12144;
  assign n12148 = ~n12146 | ~n11059;
  assign n12147 = ~n13535 | ~P2_STATE_REG_SCAN_IN;
  assign n12150 = n12148 & n12147;
  assign n12149 = ~n14577 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P2_U3344 = ~n12150 | ~n12149;
  assign n12152 = ~P2_DATAO_REG_24__SCAN_IN | ~n13390;
  assign n12151 = ~P2_U3966 | ~n16363;
  assign P2_U3576 = ~n12152 | ~n12151;
  assign n12155 = n12154 | n12153;
  assign n12179 = ~P1_REG0_REG_1__SCAN_IN | ~n15801;
  assign n16558 = ~n16974;
  assign n12168 = ~n16558 & ~n16553;
  assign n12276 = ~n16554;
  assign n12159 = ~n12168 & ~n12276;
  assign n12161 = ~n12159 & ~n15738;
  assign n12160 = ~n16563 | ~n16974;
  assign n12166 = ~n12161 | ~n12160;
  assign n12162 = ~n12534;
  assign n12164 = ~n12162 & ~n15594;
  assign n12163 = ~n16562 & ~n15595;
  assign n12165 = ~n12164 & ~n12163;
  assign n12170 = ~n12166 | ~n12165;
  assign n12520 = ~n12168 ^ n12167;
  assign n12169 = ~n12520 & ~n15404;
  assign n12525 = ~n12170 & ~n12169;
  assign n12176 = ~n12520 & ~n15619;
  assign n12172 = ~n12560;
  assign n12171 = ~n12542 | ~n12282;
  assign n12519 = ~n12172 | ~n12171;
  assign n12174 = n12519 | n15185;
  assign n12173 = ~n12542 | ~n15793;
  assign n12175 = ~n12174 | ~n12173;
  assign n12177 = ~n12176 & ~n12175;
  assign n12183 = ~n12525 | ~n12177;
  assign n12178 = ~n15800 | ~n12183;
  assign P1_U3457 = ~n12179 | ~n12178;
  assign n12185 = ~P1_REG1_REG_1__SCAN_IN | ~n15806;
  assign n12184 = ~n15804 | ~n12183;
  assign P1_U3524 = ~n12185 | ~n12184;
  assign n12191 = n14882 & n12186;
  assign n12189 = ~n11932 | ~n12187;
  assign n12188 = ~n14887;
  assign n12190 = ~n12189 | ~n12188;
  assign n12192 = ~n12191 & ~n12190;
  assign n12196 = ~n12192 & ~n10261;
  assign n12194 = ~P2_ADDR_REG_0__SCAN_IN | ~n14864;
  assign n12193 = ~P2_REG3_REG_0__SCAN_IN | ~P2_U3152;
  assign n12195 = ~n12194 | ~n12193;
  assign n12201 = ~n12196 & ~n12195;
  assign n12198 = ~n11932 | ~P2_REG1_REG_0__SCAN_IN;
  assign n12197 = ~n14882 | ~P2_REG2_REG_0__SCAN_IN;
  assign n12199 = ~n12198 | ~n12197;
  assign n12200 = ~n12199 | ~n10261;
  assign P2_U3245 = ~n12201 | ~n12200;
  assign n12401 = ~P2_REG3_REG_3__SCAN_IN | ~P2_U3152;
  assign n12202 = ~n14864 | ~P2_ADDR_REG_3__SCAN_IN;
  assign n12216 = ~n12401 | ~n12202;
  assign n12205 = ~n12204 & ~n12203;
  assign n12207 = ~n12917 & ~n12205;
  assign n12214 = ~n12207 | ~n12206;
  assign n12210 = ~n12209 & ~n12208;
  assign n12212 = ~n12210 & ~n12924;
  assign n12213 = ~n12212 | ~n12211;
  assign n12215 = ~n12214 | ~n12213;
  assign n12219 = ~n12216 & ~n12215;
  assign n12218 = ~n14887 | ~n12217;
  assign P2_U3248 = ~n12219 | ~n12218;
  assign n12221 = ~P2_ADDR_REG_2__SCAN_IN | ~n14864;
  assign n12220 = ~P2_REG3_REG_2__SCAN_IN | ~P2_U3152;
  assign n12235 = ~n12221 | ~n12220;
  assign n12224 = ~n12223 & ~n12222;
  assign n12226 = ~n12917 & ~n12224;
  assign n12233 = ~n12226 | ~n12225;
  assign n12229 = ~n12228 & ~n12227;
  assign n12231 = ~n12229 & ~n12924;
  assign n12232 = ~n12231 | ~n12230;
  assign n12234 = ~n12233 | ~n12232;
  assign n12238 = ~n12235 & ~n12234;
  assign n12237 = ~n14887 | ~n12236;
  assign P2_U3247 = ~n12238 | ~n12237;
  assign n12241 = ~n12240 & ~n12239;
  assign n12243 = ~n12241 & ~n12924;
  assign n12245 = ~n12243 | ~n12242;
  assign n12244 = ~P2_REG3_REG_1__SCAN_IN | ~P2_U3152;
  assign n12254 = ~n12245 | ~n12244;
  assign n12252 = ~P2_ADDR_REG_1__SCAN_IN | ~n14864;
  assign n12248 = ~n12247 & ~n12246;
  assign n12250 = ~n12917 & ~n12248;
  assign n12251 = ~n12250 | ~n12249;
  assign n12253 = ~n12252 | ~n12251;
  assign n12257 = ~n12254 & ~n12253;
  assign n12256 = ~n14887 | ~n12255;
  assign P2_U3246 = ~n12257 | ~n12256;
  assign n13015 = ~P2_REG3_REG_6__SCAN_IN | ~P2_U3152;
  assign n12258 = ~n14864 | ~P2_ADDR_REG_6__SCAN_IN;
  assign n12272 = ~n13015 | ~n12258;
  assign n12261 = ~n12260 & ~n12259;
  assign n12263 = ~n12261 & ~n12917;
  assign n12270 = ~n12263 | ~n12262;
  assign n12266 = ~n12265 & ~n12264;
  assign n12268 = ~n12266 & ~n12924;
  assign n12269 = ~n12268 | ~n12267;
  assign n12271 = ~n12270 | ~n12269;
  assign n12275 = ~n12272 & ~n12271;
  assign n12274 = ~n14887 | ~n12273;
  assign P2_U3251 = ~n12275 | ~n12274;
  assign n12287 = ~P1_REG1_REG_0__SCAN_IN | ~n15806;
  assign n16975 = ~n12534 | ~n12934;
  assign n12936 = ~n12276 | ~n16975;
  assign n12277 = ~n15404 | ~n15738;
  assign n12279 = ~n12936 | ~n12277;
  assign n12278 = ~n12629 | ~n15636;
  assign n12942 = n12279 & n12278;
  assign n12280 = ~n15619;
  assign n12284 = ~n12936 | ~n12280;
  assign n12283 = ~n12282 | ~n12281;
  assign n12285 = n12284 & n12283;
  assign n12288 = ~n12942 | ~n12285;
  assign n12286 = ~n15804 | ~n12288;
  assign P1_U3523 = ~n12287 | ~n12286;
  assign n12290 = ~P1_REG0_REG_0__SCAN_IN | ~n15801;
  assign n12289 = ~n15800 | ~n12288;
  assign P1_U3454 = ~n12290 | ~n12289;
  assign n12292 = ~n12295 | ~n11059;
  assign n12291 = ~n13874 | ~P2_STATE_REG_SCAN_IN;
  assign n12294 = n12292 & n12291;
  assign n12293 = ~n14577 | ~P1_DATAO_REG_15__SCAN_IN;
  assign P2_U3343 = ~n12294 | ~n12293;
  assign n12297 = ~n12295 | ~n14582;
  assign n13771 = ~n13461;
  assign n12296 = ~n13771 | ~P1_STATE_REG_SCAN_IN;
  assign n12299 = n12297 & n12296;
  assign n12298 = ~n14388 | ~P2_DATAO_REG_15__SCAN_IN;
  assign P1_U3338 = ~n12299 | ~n12298;
  assign n14165 = ~P2_REG3_REG_12__SCAN_IN | ~P2_U3152;
  assign n12300 = ~n14864 | ~P2_ADDR_REG_12__SCAN_IN;
  assign n12316 = ~n14165 | ~n12300;
  assign n12304 = ~P2_REG1_REG_11__SCAN_IN & ~n12306;
  assign n12576 = P2_REG1_REG_12__SCAN_IN ^ n12311;
  assign n12305 = ~n12577 ^ n12576;
  assign n12314 = ~n12305 | ~n11932;
  assign n12310 = ~P2_REG2_REG_11__SCAN_IN & ~n12306;
  assign n12312 = ~n12583 ^ n12582;
  assign n12313 = ~n12312 | ~n14882;
  assign n12315 = ~n12314 | ~n12313;
  assign n12318 = ~n12316 & ~n12315;
  assign n12317 = ~n14887 | ~n12581;
  assign P2_U3257 = ~n12318 | ~n12317;
  assign n12322 = ~n12320 & ~n12319;
  assign ADD_1071_U60 = n12322 ^ n12321;
  assign n12333 = ~n14448 & ~n16090;
  assign n12324 = ~n15535 & ~n16076;
  assign n12323 = ~n15872 & ~n16081;
  assign n12331 = ~n12324 & ~n12323;
  assign n12328 = n12326 | n12325;
  assign n12329 = ~n12328 | ~n12327;
  assign n12330 = ~n15527 | ~n12329;
  assign n12332 = ~n12331 | ~n12330;
  assign n12336 = ~n12333 & ~n12332;
  assign n12420 = n12334 | n16486;
  assign n12335 = ~P2_REG3_REG_1__SCAN_IN | ~n12420;
  assign P2_U3224 = ~n12336 | ~n12335;
  assign n12358 = ~P2_REG1_REG_1__SCAN_IN | ~n16516;
  assign n15972 = ~n12346;
  assign n12337 = ~n16084;
  assign n12339 = ~n15972 | ~n12337;
  assign n12340 = ~n12339 | ~n12338;
  assign n12344 = ~n12340 | ~n15832;
  assign n12342 = ~n16081 & ~n16488;
  assign n12341 = ~n16076 & ~n15713;
  assign n12343 = ~n12342 & ~n12341;
  assign n12349 = ~n12344 | ~n12343;
  assign n12815 = ~n12346 ^ n12345;
  assign n12347 = ~n12815;
  assign n12348 = ~n12347 & ~n14769;
  assign n12811 = ~n12349 & ~n12348;
  assign n12350 = ~n12351 | ~n10645;
  assign n12807 = ~n12900 | ~n12350;
  assign n12355 = ~n12807 & ~n14995;
  assign n12353 = ~n12815 | ~n14993;
  assign n12352 = ~n12351 | ~n16502;
  assign n12354 = ~n12353 | ~n12352;
  assign n12356 = ~n12355 & ~n12354;
  assign n12359 = ~n12811 | ~n12356;
  assign n12357 = ~n16514 | ~n12359;
  assign P2_U3521 = ~n12358 | ~n12357;
  assign n12361 = ~P2_REG0_REG_1__SCAN_IN | ~n16511;
  assign n12360 = ~n16510 | ~n12359;
  assign P2_U3454 = ~n12361 | ~n12360;
  assign n12379 = ~P1_REG1_REG_5__SCAN_IN | ~n15806;
  assign n12363 = ~n16979 ^ n12362;
  assign n12367 = ~n12363 & ~n15738;
  assign n12365 = ~n12495 | ~n17091;
  assign n12364 = ~n16595 | ~n15636;
  assign n12366 = ~n12365 | ~n12364;
  assign n12444 = ~n12367 & ~n12366;
  assign n12368 = ~n12505 | ~n12794;
  assign n12369 = ~n12368 | ~n12435;
  assign n12371 = ~n12369 | ~n15791;
  assign n12439 = ~n12371 & ~n12370;
  assign n12438 = n12373 ^ n12372;
  assign n14935 = ~n15404 | ~n15619;
  assign n12375 = ~n12438 | ~n14935;
  assign n12374 = ~n12435 | ~n15793;
  assign n12376 = ~n12375 | ~n12374;
  assign n12377 = ~n12439 & ~n12376;
  assign n12380 = ~n12444 | ~n12377;
  assign n12378 = ~n15804 | ~n12380;
  assign P1_U3528 = ~n12379 | ~n12378;
  assign n12382 = ~P1_REG0_REG_5__SCAN_IN | ~n15801;
  assign n12381 = ~n15800 | ~n12380;
  assign P1_U3469 = ~n12382 | ~n12381;
  assign n12394 = ~P2_REG3_REG_0__SCAN_IN | ~n12420;
  assign n12392 = ~n14448 & ~n16071;
  assign n12384 = ~n12383 | ~n12806;
  assign n12385 = ~n12384 | ~n16071;
  assign n12387 = n12386 & n12385;
  assign n12390 = ~n15527 | ~n12387;
  assign n12389 = ~n15869 | ~n12388;
  assign n12391 = ~n12390 | ~n12389;
  assign n12393 = ~n12392 & ~n12391;
  assign P2_U3234 = ~n12394 | ~n12393;
  assign n12396 = ~n12427 & ~n14384;
  assign n12395 = ~n13774 & ~P1_U3084;
  assign n12398 = ~n12396 & ~n12395;
  assign n12397 = ~n14388 | ~P2_DATAO_REG_16__SCAN_IN;
  assign P1_U3337 = ~n12398 | ~n12397;
  assign n12404 = ~P2_REG3_REG_3__SCAN_IN & ~n15865;
  assign n12400 = ~n15535 & ~n12890;
  assign n12399 = ~n15872 & ~n16076;
  assign n12402 = ~n12400 & ~n12399;
  assign n12403 = ~n12402 | ~n12401;
  assign n12411 = ~n12404 & ~n12403;
  assign n12409 = ~n14448 & ~n16125;
  assign n12407 = ~n12406 ^ n12405;
  assign n12408 = ~n15861 & ~n12407;
  assign n12410 = ~n12409 & ~n12408;
  assign P2_U3220 = ~n12411 | ~n12410;
  assign n12413 = ~n15535 & ~n16124;
  assign n12412 = ~n15872 & ~n16070;
  assign n12426 = ~n12413 & ~n12412;
  assign n12417 = ~n12416 | ~n12415;
  assign n12419 = ~n12418 | ~n12417;
  assign n12424 = ~n15861 & ~n12419;
  assign n12422 = ~P2_REG3_REG_2__SCAN_IN | ~n12420;
  assign n12421 = ~n15867 | ~n16093;
  assign n12423 = ~n12422 | ~n12421;
  assign n12425 = ~n12424 & ~n12423;
  assign P2_U3239 = ~n12426 | ~n12425;
  assign n12430 = ~n12427 & ~n14094;
  assign n12428 = ~n14425;
  assign n12429 = ~n12428 & ~P2_U3152;
  assign n12432 = ~n12430 & ~n12429;
  assign n12431 = ~n14577 | ~P1_DATAO_REG_16__SCAN_IN;
  assign P2_U3342 = ~n12432 | ~n12431;
  assign n12434 = ~P2_DATAO_REG_25__SCAN_IN | ~n13390;
  assign n12433 = ~P2_U3966 | ~n15463;
  assign P2_U3577 = ~n12434 | ~n12433;
  assign n12437 = ~n12435 | ~n13968;
  assign n12436 = ~n15407 | ~n12818;
  assign n12443 = ~n12437 | ~n12436;
  assign n12441 = ~n12438 | ~n14655;
  assign n12440 = ~n12439 | ~n17072;
  assign n12442 = ~n12441 | ~n12440;
  assign n12445 = ~n12443 & ~n12442;
  assign n12446 = ~n12445 | ~n12444;
  assign n12448 = ~n15745 | ~n12446;
  assign n12447 = ~n15218 | ~P1_REG2_REG_5__SCAN_IN;
  assign P1_U3286 = ~n12448 | ~n12447;
  assign n12465 = ~P1_REG1_REG_4__SCAN_IN | ~n15806;
  assign n12450 = n16972 ^ n12449;
  assign n12455 = ~n12450 | ~n10774;
  assign n12453 = ~n16568 & ~n15594;
  assign n12452 = ~n12451 & ~n15595;
  assign n12454 = ~n12453 & ~n12452;
  assign n12458 = ~n12455 | ~n12454;
  assign n12790 = n16972 ^ n12456;
  assign n12457 = ~n12790 & ~n15404;
  assign n12788 = ~n12458 & ~n12457;
  assign n12462 = ~n12790 & ~n15619;
  assign n12801 = n12505 ^ n12794;
  assign n12460 = ~n12801 | ~n15791;
  assign n12459 = ~n12668 | ~n15793;
  assign n12461 = ~n12460 | ~n12459;
  assign n12463 = ~n12462 & ~n12461;
  assign n12466 = ~n12788 | ~n12463;
  assign n12464 = ~n15804 | ~n12466;
  assign P1_U3527 = ~n12465 | ~n12464;
  assign n12468 = ~P1_REG0_REG_4__SCAN_IN | ~n15801;
  assign n12467 = ~n15800 | ~n12466;
  assign P1_U3466 = ~n12468 | ~n12467;
  assign n12473 = P1_REG1_REG_13__SCAN_IN ^ n12983;
  assign n12476 = ~n12473 & ~n12474;
  assign n12475 = ~n14333 | ~n12984;
  assign n12491 = ~n12476 & ~n12475;
  assign n12482 = P1_REG2_REG_13__SCAN_IN ^ n12983;
  assign n12481 = ~P1_REG2_REG_12__SCAN_IN & ~n12477;
  assign n12485 = ~n12482 & ~n12483;
  assign n12484 = ~n12976 | ~n14325;
  assign n12487 = ~n12485 & ~n12484;
  assign n12486 = ~P1_REG3_REG_13__SCAN_IN;
  assign n13853 = ~n12486 & ~P1_STATE_REG_SCAN_IN;
  assign n12489 = ~n12487 & ~n13853;
  assign n12488 = ~n14837 | ~n12983;
  assign n12490 = ~n12489 | ~n12488;
  assign n12493 = ~n12491 & ~n12490;
  assign n12492 = ~P1_ADDR_REG_13__SCAN_IN | ~n14842;
  assign P1_U3254 = ~n12493 | ~n12492;
  assign n12515 = ~P1_REG0_REG_3__SCAN_IN | ~n15801;
  assign n12494 = ~n16896 ^ n16971;
  assign n12499 = ~n12494 & ~n15738;
  assign n12497 = ~n12495 | ~n15636;
  assign n12496 = ~n12721 | ~n17091;
  assign n12498 = ~n12497 | ~n12496;
  assign n12715 = ~n12499 & ~n12498;
  assign n12504 = ~n12500;
  assign n12503 = ~n12502 & ~n12501;
  assign n12714 = ~n12504 & ~n12503;
  assign n12512 = ~n12714 & ~n15789;
  assign n12508 = ~n12505;
  assign n12507 = ~n12506 | ~n12720;
  assign n12707 = ~n12508 | ~n12507;
  assign n12510 = n12707 | n15185;
  assign n12509 = ~n12720 | ~n15793;
  assign n12511 = ~n12510 | ~n12509;
  assign n12513 = ~n12512 & ~n12511;
  assign n12516 = ~n12715 | ~n12513;
  assign n12514 = ~n15800 | ~n12516;
  assign P1_U3463 = ~n12515 | ~n12514;
  assign n12518 = ~P1_REG1_REG_3__SCAN_IN | ~n15806;
  assign n12517 = ~n15804 | ~n12516;
  assign P1_U3526 = ~n12518 | ~n12517;
  assign n12531 = ~n15174 & ~n12519;
  assign n12524 = ~n12520 & ~n13107;
  assign n12523 = ~n12522 & ~n12521;
  assign n12526 = ~n12524 & ~n12523;
  assign n12527 = ~n12526 | ~n12525;
  assign n12529 = ~n15745 | ~n12527;
  assign n12528 = ~n15218 | ~P1_REG2_REG_1__SCAN_IN;
  assign n12530 = ~n12529 | ~n12528;
  assign n12533 = ~n12531 & ~n12530;
  assign n12532 = ~P1_REG3_REG_1__SCAN_IN | ~n15407;
  assign P1_U3290 = ~n12533 | ~n12532;
  assign n12536 = ~n17132 | ~n12721;
  assign n12535 = ~n15696 | ~n12534;
  assign n12546 = ~n12536 | ~n12535;
  assign n12540 = ~n12538 | ~n12537;
  assign n12541 = n12540 ^ n12539;
  assign n12544 = ~n12541 | ~n10132;
  assign n12543 = ~n15578 | ~n12542;
  assign n12545 = ~n12544 | ~n12543;
  assign n12548 = ~n12546 & ~n12545;
  assign n12547 = ~P1_REG3_REG_1__SCAN_IN | ~n12628;
  assign P1_U3220 = ~n12548 | ~n12547;
  assign n12567 = ~P1_REG0_REG_2__SCAN_IN | ~n15801;
  assign n12963 = n12549 ^ n16969;
  assign n12558 = ~n12963 & ~n15404;
  assign n12552 = ~n16568 & ~n15595;
  assign n12551 = ~n12550 & ~n15594;
  assign n12556 = ~n12552 & ~n12551;
  assign n12554 = ~n16969 ^ n12553;
  assign n12555 = ~n12554 | ~n10774;
  assign n12557 = ~n12556 | ~n12555;
  assign n12962 = ~n12558 & ~n12557;
  assign n12564 = ~n12963 & ~n15619;
  assign n12972 = n12560 ^ n12559;
  assign n12562 = ~n12972 | ~n15791;
  assign n12561 = ~n16561 | ~n15793;
  assign n12563 = ~n12562 | ~n12561;
  assign n12565 = ~n12564 & ~n12563;
  assign n12568 = ~n12962 | ~n12565;
  assign n12566 = ~n15800 | ~n12568;
  assign P1_U3460 = ~n12567 | ~n12566;
  assign n12570 = ~P1_REG1_REG_2__SCAN_IN | ~n15806;
  assign n12569 = ~n15804 | ~n12568;
  assign P1_U3525 = ~n12570 | ~n12569;
  assign n12574 = ~n12572 & ~n12571;
  assign ADD_1071_U59 = n12574 ^ n12573;
  assign n14243 = ~P2_REG3_REG_13__SCAN_IN | ~P2_U3152;
  assign n12575 = ~n14864 | ~P2_ADDR_REG_13__SCAN_IN;
  assign n12591 = ~n14243 | ~n12575;
  assign n12579 = ~P2_REG1_REG_12__SCAN_IN & ~n12581;
  assign n12580 = ~n12914 ^ n12913;
  assign n12589 = ~n12580 | ~n11932;
  assign n12585 = ~P2_REG2_REG_12__SCAN_IN & ~n12581;
  assign n12587 = ~n12921 ^ n12920;
  assign n12588 = ~n12587 | ~n14882;
  assign n12590 = ~n12589 | ~n12588;
  assign n12593 = ~n12591 & ~n12590;
  assign n12592 = ~n14887 | ~n12919;
  assign P2_U3258 = ~n12593 | ~n12592;
  assign n12609 = ~P2_REG0_REG_2__SCAN_IN | ~n16511;
  assign n15975 = n16076 ^ n13050;
  assign n12595 = ~n15975 ^ n12594;
  assign n12598 = ~n12595 & ~n15547;
  assign n13047 = n15975 ^ n12596;
  assign n12597 = ~n13047 & ~n14769;
  assign n12602 = ~n12598 & ~n12597;
  assign n12600 = ~n16124 & ~n15713;
  assign n12599 = ~n16070 & ~n16488;
  assign n12601 = ~n12600 & ~n12599;
  assign n13058 = ~n12602 | ~n12601;
  assign n13053 = ~n12900 ^ n13050;
  assign n12604 = ~n13053 | ~n16500;
  assign n12603 = ~n16093 | ~n16502;
  assign n12605 = ~n12604 | ~n12603;
  assign n12607 = ~n13058 & ~n12605;
  assign n12606 = n13047 | n16498;
  assign n12610 = ~n12607 | ~n12606;
  assign n12608 = ~n16510 | ~n12610;
  assign P2_U3457 = ~n12609 | ~n12608;
  assign n12612 = ~P2_REG1_REG_2__SCAN_IN | ~n16516;
  assign n12611 = ~n16514 | ~n12610;
  assign P2_U3522 = ~n12612 | ~n12611;
  assign n12614 = ~n15869 | ~n13014;
  assign n12616 = ~n12614 | ~n12613;
  assign n12615 = ~n15872 & ~n16124;
  assign n12623 = ~n12616 & ~n12615;
  assign n12620 = n12618 | n12617;
  assign n12621 = ~n12620 | ~n12619;
  assign n12622 = ~n15527 | ~n12621;
  assign n12625 = ~n12623 | ~n12622;
  assign n12624 = ~n14448 & ~n16115;
  assign n12627 = ~n12625 & ~n12624;
  assign n12626 = ~n12848 | ~n15530;
  assign P2_U3232 = ~n12627 | ~n12626;
  assign n12636 = ~P1_REG3_REG_0__SCAN_IN | ~n12628;
  assign n12634 = ~n17126 & ~n12934;
  assign n12632 = ~n17132 | ~n12629;
  assign n12631 = ~n10132 | ~n12630;
  assign n12633 = ~n12632 | ~n12631;
  assign n12635 = ~n12634 & ~n12633;
  assign P1_U3230 = ~n12636 | ~n12635;
  assign n12638 = ~P2_DATAO_REG_26__SCAN_IN | ~n13390;
  assign n12637 = ~P2_U3966 | ~n15557;
  assign P2_U3578 = ~n12638 | ~n12637;
  assign n12641 = ~n12680 & ~n14384;
  assign n12639 = ~n14627;
  assign n12640 = ~n12639 & ~P1_U3084;
  assign n12643 = ~n12641 & ~n12640;
  assign n12642 = ~n14388 | ~P2_DATAO_REG_17__SCAN_IN;
  assign P1_U3336 = ~n12643 | ~n12642;
  assign n12645 = ~n15532 | ~n16116;
  assign n12648 = ~n12645 | ~n12644;
  assign n12647 = ~n15535 & ~n12646;
  assign n12660 = ~n12648 & ~n12647;
  assign n12653 = ~n12649;
  assign n12652 = ~n12651 | ~n12650;
  assign n12654 = ~n12653 | ~n12652;
  assign n12658 = ~n15861 & ~n12654;
  assign n12656 = ~n15530 | ~n13075;
  assign n12655 = ~n15867 | ~n12876;
  assign n12657 = ~n12656 | ~n12655;
  assign n12659 = ~n12658 & ~n12657;
  assign P2_U3229 = ~n12660 | ~n12659;
  assign n12662 = ~P2_DATAO_REG_27__SCAN_IN | ~n13390;
  assign n12661 = ~P2_U3966 | ~n15704;
  assign P2_U3579 = ~n12662 | ~n12661;
  assign n12679 = ~n14853 | ~n12791;
  assign n12665 = ~n12664 | ~n12663;
  assign n12667 = ~n12665 | ~n10132;
  assign n12677 = ~n12667 & ~n12666;
  assign n12670 = ~n15578 | ~n12668;
  assign n12669 = ~n17132 | ~n12763;
  assign n12675 = ~n12670 | ~n12669;
  assign n12673 = ~n15696 | ~n12671;
  assign n12674 = ~n12673 | ~n12672;
  assign n12676 = n12675 | n12674;
  assign n12678 = ~n12677 & ~n12676;
  assign P1_U3228 = ~n12679 | ~n12678;
  assign n12683 = ~n12680 & ~n14094;
  assign n12682 = ~n12681 & ~P2_U3152;
  assign n12685 = ~n12683 & ~n12682;
  assign n12684 = ~n14577 | ~P1_DATAO_REG_17__SCAN_IN;
  assign P2_U3341 = ~n12685 | ~n12684;
  assign n12703 = ~P2_REG0_REG_4__SCAN_IN | ~n16511;
  assign n12686 = ~n12873 | ~n16500;
  assign n12853 = ~n12899 & ~n16115;
  assign n12690 = ~n12686 & ~n12853;
  assign n12859 = ~n13014 | ~n15549;
  assign n12688 = ~n12687 | ~n16502;
  assign n12689 = ~n12859 | ~n12688;
  assign n12701 = ~n12690 & ~n12689;
  assign n12847 = n15976 ^ n12691;
  assign n12699 = ~n12847 & ~n16498;
  assign n12693 = ~n14769 & ~n12847;
  assign n12692 = ~n16124 & ~n16488;
  assign n12698 = ~n12693 & ~n12692;
  assign n12696 = ~n12695 ^ n12694;
  assign n12697 = ~n15832 | ~n12696;
  assign n12856 = ~n12698 | ~n12697;
  assign n12700 = ~n12699 & ~n12856;
  assign n12704 = ~n12701 | ~n12700;
  assign n12702 = ~n16510 | ~n12704;
  assign P2_U3463 = ~n12703 | ~n12702;
  assign n12706 = ~P2_REG1_REG_4__SCAN_IN | ~n16516;
  assign n12705 = ~n16514 | ~n12704;
  assign P2_U3524 = ~n12706 | ~n12705;
  assign n12713 = ~P1_REG3_REG_3__SCAN_IN & ~n15766;
  assign n12709 = ~n15174 & ~n12707;
  assign n12708 = ~n15763 & ~n16567;
  assign n12711 = ~n12709 & ~n12708;
  assign n12710 = ~P1_REG2_REG_3__SCAN_IN | ~n15218;
  assign n12712 = ~n12711 | ~n12710;
  assign n12719 = ~n12713 & ~n12712;
  assign n13829 = ~n14655;
  assign n12716 = n12714 | n13829;
  assign n12717 = ~n12716 | ~n12715;
  assign n12718 = ~n12717 | ~n15745;
  assign P1_U3288 = ~n12719 | ~n12718;
  assign n12725 = ~n14796 & ~P1_REG3_REG_3__SCAN_IN;
  assign n12723 = ~n15578 | ~n12720;
  assign n12722 = ~n15696 | ~n12721;
  assign n12724 = ~n12723 | ~n12722;
  assign n12727 = ~n12725 & ~n12724;
  assign n12729 = ~n12727 | ~n12726;
  assign n12728 = ~n15689 & ~n12825;
  assign n12734 = ~n12729 & ~n12728;
  assign n12732 = ~n12731 ^ n12730;
  assign n12733 = ~n12732 | ~n10132;
  assign P1_U3216 = ~n12734 | ~n12733;
  assign n12744 = ~P1_REG1_REG_6__SCAN_IN | ~n15806;
  assign n12737 = ~n12735 | ~n15791;
  assign n12736 = ~n13114 | ~n15793;
  assign n12742 = n12737 & n12736;
  assign n12740 = ~n12738 & ~n15619;
  assign n12741 = ~n12740 & ~n12739;
  assign n12743 = ~n15804 | ~n12745;
  assign P1_U3529 = ~n12744 | ~n12743;
  assign n12747 = ~P1_REG0_REG_6__SCAN_IN | ~n15801;
  assign n12746 = ~n15800 | ~n12745;
  assign P1_U3472 = ~n12747 | ~n12746;
  assign n12750 = ~n12749 | ~n12748;
  assign n12752 = ~n12751 ^ n12750;
  assign n12760 = ~n12752 & ~n17147;
  assign n12754 = ~n17126 & ~n13424;
  assign n12753 = ~n17136 & ~n13371;
  assign n12758 = ~n12754 & ~n12753;
  assign n12756 = ~n15689 & ~n13366;
  assign n12757 = ~n12756 & ~n12755;
  assign n12759 = ~n12758 | ~n12757;
  assign n12762 = ~n12760 & ~n12759;
  assign n12761 = ~n14853 | ~n13420;
  assign P1_U3211 = ~n12762 | ~n12761;
  assign n12765 = ~n15578 | ~n13114;
  assign n12764 = ~n15696 | ~n12763;
  assign n12773 = ~n12765 | ~n12764;
  assign n12771 = ~n17132 | ~n13104;
  assign n12769 = ~n12766;
  assign n12768 = ~n14796 & ~n12767;
  assign n12770 = ~n12769 & ~n12768;
  assign n12772 = ~n12771 | ~n12770;
  assign n12787 = ~n12773 & ~n12772;
  assign n12820 = n12775 ^ n12776;
  assign n12778 = ~n12820 | ~n12774;
  assign n12777 = ~n12776 | ~n12775;
  assign n12784 = ~n12778 | ~n12777;
  assign n12782 = ~n12780 | ~n12779;
  assign n12783 = ~n12782 | ~n12781;
  assign n12785 = n12784 ^ n12783;
  assign n12786 = ~n12785 | ~n10132;
  assign P1_U3237 = ~n12787 | ~n12786;
  assign n12800 = ~n15218 & ~n12788;
  assign n15608 = ~n15745 | ~n12789;
  assign n12798 = n12790 | n15608;
  assign n12793 = ~n15218 | ~P1_REG2_REG_4__SCAN_IN;
  assign n12792 = ~n15407 | ~n12791;
  assign n12796 = ~n12793 | ~n12792;
  assign n12795 = ~n15763 & ~n12794;
  assign n12797 = ~n12796 & ~n12795;
  assign n12799 = ~n12798 | ~n12797;
  assign n12803 = ~n12800 & ~n12799;
  assign n12802 = ~n15762 | ~n12801;
  assign P1_U3287 = ~n12803 | ~n12802;
  assign n12805 = ~n15488 | ~P2_REG2_REG_1__SCAN_IN;
  assign n12804 = ~n15725 | ~P2_REG3_REG_1__SCAN_IN;
  assign n12814 = ~n12805 | ~n12804;
  assign n12809 = ~n12807 & ~n12806;
  assign n12808 = ~n16090 & ~n12855;
  assign n12810 = ~n12809 & ~n12808;
  assign n12812 = n12811 & n12810;
  assign n12813 = ~n15488 & ~n12812;
  assign n12817 = ~n12814 & ~n12813;
  assign n12816 = ~n14078 | ~n12815;
  assign P2_U3295 = ~n12817 | ~n12816;
  assign n12833 = ~n14853 | ~n12818;
  assign n12821 = ~n12820 ^ n12819;
  assign n12831 = ~n12821 & ~n17147;
  assign n12824 = ~n17126 & ~n12822;
  assign n12823 = ~n15689 & ~n13371;
  assign n12829 = ~n12824 & ~n12823;
  assign n12827 = ~n17136 & ~n12825;
  assign n12828 = ~n12827 & ~n12826;
  assign n12830 = ~n12829 | ~n12828;
  assign n12832 = ~n12831 & ~n12830;
  assign P1_U3225 = ~n12833 | ~n12832;
  assign n12837 = ~n12835 & ~n12834;
  assign ADD_1071_U58 = n12837 ^ n12836;
  assign n12839 = ~n12842 | ~n14582;
  assign n12838 = ~n14828 | ~P1_STATE_REG_SCAN_IN;
  assign n12841 = n12839 & n12838;
  assign n12840 = ~n14388 | ~P2_DATAO_REG_18__SCAN_IN;
  assign P1_U3335 = ~n12841 | ~n12840;
  assign n12844 = ~n12842 | ~n11059;
  assign n12843 = ~n14876 | ~P2_STATE_REG_SCAN_IN;
  assign n12846 = n12844 & n12843;
  assign n12845 = ~n14577 | ~P1_DATAO_REG_18__SCAN_IN;
  assign P2_U3340 = ~n12846 | ~n12845;
  assign n12852 = ~n15845 & ~n12847;
  assign n12850 = ~n15725 | ~n12848;
  assign n12849 = ~n15488 | ~P2_REG2_REG_4__SCAN_IN;
  assign n12851 = ~n12850 | ~n12849;
  assign n12864 = ~n12852 & ~n12851;
  assign n12854 = ~n12873 | ~n10888;
  assign n12861 = ~n12854 & ~n12853;
  assign n12857 = ~n16115 & ~n12855;
  assign n12858 = ~n12857 & ~n12856;
  assign n12860 = ~n12859 | ~n12858;
  assign n12862 = n12861 | n12860;
  assign n12863 = ~n12862 | ~n15720;
  assign P2_U3292 = ~n12864 | ~n12863;
  assign n12884 = ~P2_REG1_REG_5__SCAN_IN | ~n16516;
  assign n13085 = n12866 ^ n12865;
  assign n12868 = ~n13085 | ~n10644;
  assign n12867 = ~n16116 | ~n15550;
  assign n12872 = ~n12868 | ~n12867;
  assign n12870 = ~n15969 ^ n12869;
  assign n12871 = ~n12870 & ~n15547;
  assign n13073 = ~n12872 & ~n12871;
  assign n12881 = ~n13085 | ~n14993;
  assign n12875 = ~n13003;
  assign n12874 = ~n12873 | ~n12876;
  assign n13070 = ~n12875 | ~n12874;
  assign n12879 = ~n13070 & ~n14995;
  assign n13072 = ~n13251 | ~n15549;
  assign n12877 = ~n12876 | ~n16502;
  assign n12878 = ~n13072 | ~n12877;
  assign n12880 = ~n12879 & ~n12878;
  assign n12882 = n12881 & n12880;
  assign n12885 = ~n13073 | ~n12882;
  assign n12883 = ~n16514 | ~n12885;
  assign P2_U3525 = ~n12884 | ~n12883;
  assign n12887 = ~P2_REG0_REG_5__SCAN_IN | ~n16511;
  assign n12886 = ~n16510 | ~n12885;
  assign P2_U3466 = ~n12887 | ~n12886;
  assign n12909 = ~P2_REG1_REG_3__SCAN_IN | ~n16516;
  assign n13143 = n12889 ^ n12888;
  assign n12894 = ~n13143 | ~n10644;
  assign n12892 = ~n16076 & ~n16488;
  assign n12891 = ~n12890 & ~n15713;
  assign n12893 = ~n12892 & ~n12891;
  assign n12898 = ~n12894 | ~n12893;
  assign n12896 = ~n12895 ^ n15971;
  assign n12897 = ~n12896 & ~n15547;
  assign n13139 = ~n12898 & ~n12897;
  assign n12903 = n12899 | n14995;
  assign n12901 = ~n12900 & ~n16093;
  assign n12902 = ~n12901 & ~n16125;
  assign n13137 = ~n12903 & ~n12902;
  assign n12905 = ~n13143 | ~n14993;
  assign n12904 = ~n13144 | ~n16502;
  assign n12906 = ~n12905 | ~n12904;
  assign n12907 = ~n13137 & ~n12906;
  assign n12910 = ~n13139 | ~n12907;
  assign n12908 = ~n16514 | ~n12910;
  assign P2_U3523 = ~n12909 | ~n12908;
  assign n12912 = ~P2_REG0_REG_3__SCAN_IN | ~n16511;
  assign n12911 = ~n16510 | ~n12910;
  assign P2_U3460 = ~n12912 | ~n12911;
  assign n12916 = ~P2_REG1_REG_13__SCAN_IN & ~n12919;
  assign n12918 = n13531 ^ n13530;
  assign n12931 = ~n12918 & ~n12917;
  assign n12923 = ~P2_REG2_REG_13__SCAN_IN & ~n12919;
  assign n12925 = n13537 ^ n13536;
  assign n12927 = ~n12925 & ~n12924;
  assign n12929 = ~n12927 & ~n12926;
  assign n12928 = ~n14864 | ~P2_ADDR_REG_14__SCAN_IN;
  assign n12930 = ~n12929 | ~n12928;
  assign n12933 = ~n12931 & ~n12930;
  assign n12932 = ~n14887 | ~n13535;
  assign P2_U3259 = ~n12933 | ~n12932;
  assign n12935 = ~n15762 & ~n15313;
  assign n12941 = ~n12935 & ~n12934;
  assign n12937 = ~n15608;
  assign n12939 = ~n12937 | ~n12936;
  assign n12938 = ~P1_REG2_REG_0__SCAN_IN | ~n15218;
  assign n12940 = ~n12939 | ~n12938;
  assign n12946 = ~n12941 & ~n12940;
  assign n12943 = ~P1_REG3_REG_0__SCAN_IN | ~n15407;
  assign n12944 = ~n12943 | ~n12942;
  assign n12945 = ~n12944 | ~n15745;
  assign P1_U3291 = ~n12946 | ~n12945;
  assign n12950 = ~n13130 & ~n14796;
  assign n12948 = ~n15578 | ~n13223;
  assign n12947 = ~n15696 | ~n13104;
  assign n12949 = ~n12948 | ~n12947;
  assign n12952 = ~n12950 & ~n12949;
  assign n12954 = ~n12952 | ~n12951;
  assign n12953 = ~n15689 & ~n16629;
  assign n12961 = ~n12954 & ~n12953;
  assign n12958 = ~n12956 | ~n12955;
  assign n12959 = ~n12958 ^ n12957;
  assign n12960 = ~n12959 | ~n10132;
  assign P1_U3219 = ~n12961 | ~n12960;
  assign n12971 = ~n15218 & ~n12962;
  assign n12967 = ~n15608 & ~n12963;
  assign n12965 = ~n15313 | ~n16561;
  assign n12964 = ~n15218 | ~P1_REG2_REG_2__SCAN_IN;
  assign n12966 = ~n12965 | ~n12964;
  assign n12969 = ~n12967 & ~n12966;
  assign n12968 = ~P1_REG3_REG_2__SCAN_IN | ~n15407;
  assign n12970 = ~n12969 | ~n12968;
  assign n12974 = ~n12971 & ~n12970;
  assign n12973 = ~n15762 | ~n12972;
  assign P1_U3289 = ~n12974 | ~n12973;
  assign n14187 = ~P1_U3084 | ~P1_REG3_REG_14__SCAN_IN;
  assign n12975 = ~n14837 | ~n13458;
  assign n12982 = ~n14187 | ~n12975;
  assign n12980 = ~n14842 | ~P1_ADDR_REG_14__SCAN_IN;
  assign n12977 = ~P1_REG2_REG_13__SCAN_IN | ~n12983;
  assign n12978 = ~n13452 ^ n13451;
  assign n12979 = ~n12978 | ~n14325;
  assign n12981 = ~n12980 | ~n12979;
  assign n12992 = ~n12982 & ~n12981;
  assign n12985 = ~P1_REG1_REG_13__SCAN_IN | ~n12983;
  assign n12989 = ~P1_REG1_REG_14__SCAN_IN ^ n12986;
  assign n12987 = ~n12988 & ~n12989;
  assign n12990 = ~n12987 & ~n14833;
  assign n12991 = ~n12990 | ~n13459;
  assign P1_U3255 = ~n12992 | ~n12991;
  assign n13010 = ~P2_REG1_REG_6__SCAN_IN | ~n16516;
  assign n13039 = n15977 ^ n12993;
  assign n12998 = ~n13039 | ~n10644;
  assign n12996 = ~n13017 & ~n15713;
  assign n12995 = ~n12994 & ~n16488;
  assign n12997 = ~n12996 & ~n12995;
  assign n13002 = ~n12998 | ~n12997;
  assign n13000 = n15977 ^ n12999;
  assign n13001 = ~n13000 & ~n15547;
  assign n13044 = n13002 | n13001;
  assign n13038 = n13003 ^ n13032;
  assign n13005 = ~n13038 | ~n16500;
  assign n13004 = ~n13020 | ~n16502;
  assign n13006 = ~n13005 | ~n13004;
  assign n13008 = ~n13044 & ~n13006;
  assign n13007 = ~n13039 | ~n14993;
  assign n13009 = ~n16514 | ~n13011;
  assign P2_U3526 = ~n13010 | ~n13009;
  assign n13013 = ~P2_REG0_REG_6__SCAN_IN | ~n16511;
  assign n13012 = ~n16510 | ~n13011;
  assign P2_U3469 = ~n13013 | ~n13012;
  assign n13016 = ~n15532 | ~n13014;
  assign n13019 = ~n13016 | ~n13015;
  assign n13018 = ~n15535 & ~n13017;
  assign n13031 = ~n13019 & ~n13018;
  assign n13029 = ~n13033 & ~n15865;
  assign n13027 = ~n15867 | ~n13020;
  assign n13023 = ~n13022 | ~n13021;
  assign n13025 = n13024 ^ n13023;
  assign n13026 = ~n15527 | ~n13025;
  assign n13028 = ~n13027 | ~n13026;
  assign n13030 = ~n13029 & ~n13028;
  assign P2_U3241 = ~n13031 | ~n13030;
  assign n13035 = ~n15848 & ~n13032;
  assign n13034 = ~n15850 & ~n13033;
  assign n13037 = ~n13035 & ~n13034;
  assign n13036 = ~P2_REG2_REG_6__SCAN_IN | ~n15488;
  assign n13043 = ~n13037 | ~n13036;
  assign n13041 = ~n15847 | ~n13038;
  assign n13040 = ~n14078 | ~n13039;
  assign n13042 = ~n13041 | ~n13040;
  assign n13046 = ~n13043 & ~n13042;
  assign n13045 = ~n13044 | ~n15720;
  assign P2_U3290 = ~n13046 | ~n13045;
  assign n13057 = ~n15845 & ~n13047;
  assign n13049 = ~n15488 | ~P2_REG2_REG_2__SCAN_IN;
  assign n13048 = ~n15725 | ~P2_REG3_REG_2__SCAN_IN;
  assign n13052 = ~n13049 | ~n13048;
  assign n13051 = ~n15848 & ~n13050;
  assign n13055 = ~n13052 & ~n13051;
  assign n13054 = ~n15847 | ~n13053;
  assign n13056 = ~n13055 | ~n13054;
  assign n13060 = ~n13057 & ~n13056;
  assign n13059 = ~n13058 | ~n15720;
  assign P2_U3294 = ~n13060 | ~n13059;
  assign n13062 = ~n13065 | ~n14582;
  assign n13061 = ~n14836 | ~P1_STATE_REG_SCAN_IN;
  assign n13064 = n13062 & n13061;
  assign n13063 = ~n14388 | ~P2_DATAO_REG_19__SCAN_IN;
  assign P1_U3334 = ~n13064 | ~n13063;
  assign n13067 = ~n13065 | ~n11059;
  assign n13066 = ~n16472 | ~P2_STATE_REG_SCAN_IN;
  assign n13069 = n13067 & n13066;
  assign n13068 = ~n14577 | ~P1_DATAO_REG_19__SCAN_IN;
  assign P2_U3339 = ~n13069 | ~n13068;
  assign n13084 = ~n13071 & ~n13070;
  assign n13074 = ~n13073 | ~n13072;
  assign n13082 = ~n13074 | ~n15720;
  assign n13077 = ~n15488 | ~P2_REG2_REG_5__SCAN_IN;
  assign n13076 = ~n15725 | ~n13075;
  assign n13080 = ~n13077 | ~n13076;
  assign n13079 = ~n15848 & ~n13078;
  assign n13081 = ~n13080 & ~n13079;
  assign n13083 = ~n13082 | ~n13081;
  assign n13087 = ~n13084 & ~n13083;
  assign n13086 = ~n14078 | ~n13085;
  assign P2_U3291 = ~n13087 | ~n13086;
  assign n13089 = ~n15488 | ~P2_REG2_REG_0__SCAN_IN;
  assign n13088 = ~n15725 | ~P2_REG3_REG_0__SCAN_IN;
  assign n13092 = ~n13089 | ~n13088;
  assign n13090 = ~n15566 & ~n15847;
  assign n13091 = ~n13090 & ~n16071;
  assign n13098 = ~n13092 & ~n13091;
  assign n13096 = ~n15488 & ~n13093;
  assign n13095 = ~n15845 & ~n13094;
  assign n13097 = ~n13096 & ~n13095;
  assign P2_U3296 = ~n13098 | ~n13097;
  assign n16617 = ~n13223 | ~n13366;
  assign n13099 = ~n16596 | ~n13371;
  assign n13101 = ~n13114 | ~n16595;
  assign n13370 = ~n13102 | ~n13101;
  assign n13103 = ~n13424 | ~n13121;
  assign n13105 = ~n13364 | ~n13104;
  assign n13222 = ~n13106 | ~n13105;
  assign n13112 = ~n13160 & ~n13107;
  assign n13109 = ~n13365 | ~n13424;
  assign n13108 = ~n13109 | ~n13223;
  assign n13110 = ~n13108 | ~n15791;
  assign n13359 = ~n13109 & ~n13223;
  assign n13162 = n13110 | n13359;
  assign n13111 = ~n13162 & ~n14836;
  assign n13128 = ~n13112 & ~n13111;
  assign n13115 = ~n13113 | ~n16981;
  assign n13374 = ~n13115 | ~n16892;
  assign n16613 = ~n13364 | ~n13121;
  assign n13116 = ~n16613;
  assign n16899 = ~n13364 & ~n13121;
  assign n13119 = ~n13117 & ~n16899;
  assign n13118 = ~n13119 | ~n16985;
  assign n13120 = ~n13118 | ~n10774;
  assign n13125 = n13120 | n13350;
  assign n13123 = ~n16629 & ~n15595;
  assign n13122 = ~n13121 & ~n15594;
  assign n13124 = ~n13123 & ~n13122;
  assign n13127 = ~n13125 | ~n13124;
  assign n13126 = ~n13160 & ~n15404;
  assign n13129 = ~n13128 | ~n13166;
  assign n13136 = ~n13129 | ~n15745;
  assign n13134 = ~n15766 & ~n13130;
  assign n13132 = ~n15313 | ~n13223;
  assign n13131 = ~n15218 | ~P1_REG2_REG_8__SCAN_IN;
  assign n13133 = ~n13132 | ~n13131;
  assign n13135 = ~n13134 & ~n13133;
  assign P1_U3283 = ~n13136 | ~n13135;
  assign n13141 = ~P2_REG3_REG_3__SCAN_IN & ~n15850;
  assign n13138 = ~n13137 | ~n16038;
  assign n13140 = ~n13139 | ~n13138;
  assign n13142 = ~n13141 & ~n13140;
  assign n13148 = ~n15488 & ~n13142;
  assign n13146 = ~n14078 | ~n13143;
  assign n13145 = ~n15566 | ~n13144;
  assign n13150 = ~n13148 & ~n13147;
  assign n13149 = ~n15488 | ~P2_REG2_REG_3__SCAN_IN;
  assign P2_U3293 = ~n13150 | ~n13149;
  assign n13154 = ~n13155 | ~n14582;
  assign n13151 = n14388 & P2_DATAO_REG_20__SCAN_IN;
  assign n13153 = ~n13152 & ~n13151;
  assign P1_U3333 = ~n13154 | ~n13153;
  assign n13159 = ~n13155 | ~n11059;
  assign n13157 = ~n9039 & ~P2_U3152;
  assign n13156 = n14577 & P1_DATAO_REG_20__SCAN_IN;
  assign n13158 = ~n13157 & ~n13156;
  assign P2_U3338 = ~n13159 | ~n13158;
  assign n13168 = ~P1_REG1_REG_8__SCAN_IN | ~n15806;
  assign n13164 = ~n13160 & ~n15619;
  assign n13161 = ~n13223 | ~n15793;
  assign n13163 = ~n13162 | ~n13161;
  assign n13165 = ~n13164 & ~n13163;
  assign n13167 = ~n15804 | ~n13169;
  assign P1_U3531 = ~n13168 | ~n13167;
  assign n13171 = ~P1_REG0_REG_8__SCAN_IN | ~n15801;
  assign n13170 = ~n15800 | ~n13169;
  assign P1_U3478 = ~n13171 | ~n13170;
  assign n13177 = ~n13293 & ~n15850;
  assign n13175 = ~n14078 | ~n13399;
  assign n13174 = ~n15488 | ~P2_REG2_REG_8__SCAN_IN;
  assign n13194 = ~n13177 & ~n13176;
  assign n13179 = ~n13399 | ~n10644;
  assign n13178 = ~n13288 | ~n15550;
  assign n13183 = ~n13179 | ~n13178;
  assign n13181 = ~n15984 ^ n13180;
  assign n13182 = ~n13181 & ~n15547;
  assign n13186 = ~n13185 & ~n13184;
  assign n13187 = ~n13186 & ~n14995;
  assign n13395 = ~n13187 | ~n13309;
  assign n13190 = ~n13395 & ~n16472;
  assign n13188 = ~n16160 | ~n15285;
  assign n13393 = ~n16177 | ~n15549;
  assign n13189 = ~n13188 | ~n13393;
  assign n13191 = ~n13190 & ~n13189;
  assign n13192 = ~n13396 | ~n13191;
  assign n13193 = ~n13192 | ~n15720;
  assign P2_U3288 = ~n13194 | ~n13193;
  assign n13198 = ~n13196 & ~n13195;
  assign ADD_1071_U57 = n13198 ^ n13197;
  assign n13200 = ~n15532 | ~n13251;
  assign n13202 = ~n13200 | ~n13199;
  assign n13201 = ~n15535 & ~n13317;
  assign n13213 = ~n13202 & ~n13201;
  assign n13211 = ~n14448 & ~n13265;
  assign n13205 = ~n13204 | ~n13203;
  assign n13207 = n13206 ^ n13205;
  assign n13209 = ~n15527 | ~n13207;
  assign n13208 = ~n15530 | ~n13260;
  assign n13210 = ~n13209 | ~n13208;
  assign n13212 = ~n13211 & ~n13210;
  assign P2_U3215 = ~n13213 | ~n13212;
  assign n13215 = ~n15218 | ~P1_REG2_REG_9__SCAN_IN;
  assign n13214 = ~n13285 | ~n15407;
  assign n13219 = ~n13215 | ~n13214;
  assign n13238 = ~n13280 ^ n13359;
  assign n13217 = ~n13238 | ~n15762;
  assign n13216 = ~n15313 | ~n13280;
  assign n13218 = ~n13217 | ~n13216;
  assign n13236 = ~n13219 & ~n13218;
  assign n13588 = ~n16628 | ~n16629;
  assign n13590 = ~n13280 | ~n13474;
  assign n13220 = ~n13223;
  assign n13221 = ~n13220 | ~n13366;
  assign n13224 = ~n13223 | ~n13228;
  assign n13589 = ~n13225 | ~n13224;
  assign n13237 = n16987 ^ n13589;
  assign n13233 = n13237 | n13829;
  assign n13226 = ~n13350 & ~n16609;
  assign n13340 = ~n16987;
  assign n13227 = ~n13226 ^ n13340;
  assign n13232 = ~n13227 & ~n15738;
  assign n13230 = ~n13783 | ~n15636;
  assign n13229 = ~n13228 | ~n17091;
  assign n13231 = ~n13230 | ~n13229;
  assign n13234 = ~n13233 | ~n13244;
  assign n13235 = ~n13234 | ~n15745;
  assign P1_U3282 = ~n13236 | ~n13235;
  assign n13246 = ~P1_REG1_REG_9__SCAN_IN | ~n15806;
  assign n13242 = ~n13237 & ~n15789;
  assign n13240 = ~n13238 | ~n15791;
  assign n13239 = ~n13280 | ~n15793;
  assign n13241 = ~n13240 | ~n13239;
  assign n13243 = ~n13242 & ~n13241;
  assign n13245 = ~n15804 | ~n13247;
  assign P1_U3532 = ~n13246 | ~n13245;
  assign n13249 = ~P1_REG0_REG_9__SCAN_IN | ~n15801;
  assign n13248 = ~n15800 | ~n13247;
  assign P1_U3481 = ~n13249 | ~n13248;
  assign n13255 = n13438 & n10644;
  assign n13253 = ~n16161 | ~n15549;
  assign n13252 = ~n13251 | ~n15550;
  assign n13254 = ~n13253 | ~n13252;
  assign n13259 = ~n13255 & ~n13254;
  assign n13257 = ~n15981 ^ n13256;
  assign n13258 = ~n13257 | ~n15832;
  assign n13262 = ~n13443 | ~n15285;
  assign n13261 = ~n15725 | ~n13260;
  assign n13263 = ~n13262 | ~n13261;
  assign n13264 = ~n13442 & ~n13263;
  assign n13270 = ~n13264 & ~n15488;
  assign n13437 = ~n13266 ^ n13265;
  assign n13268 = ~n15847 | ~n13437;
  assign n13267 = ~n14078 | ~n13438;
  assign n13272 = ~n13270 & ~n13269;
  assign n13271 = ~n15488 | ~P2_REG2_REG_7__SCAN_IN;
  assign P2_U3289 = ~n13272 | ~n13271;
  assign n13275 = ~n13274 ^ n13273;
  assign n13284 = ~n13275 & ~n17147;
  assign n13277 = ~n17136 & ~n13366;
  assign n13279 = n13277 | n13276;
  assign n13278 = ~n15689 & ~n13594;
  assign n13282 = ~n13279 & ~n13278;
  assign n13281 = ~n15578 | ~n13280;
  assign n13283 = ~n13282 | ~n13281;
  assign n13287 = ~n13284 & ~n13283;
  assign n13286 = ~n14853 | ~n13285;
  assign P1_U3229 = ~n13287 | ~n13286;
  assign n13290 = ~n15532 | ~n13288;
  assign n13292 = ~n13290 | ~n13289;
  assign n13291 = ~n15535 & ~n16209;
  assign n13304 = ~n13292 & ~n13291;
  assign n13302 = ~n13293 & ~n15865;
  assign n13300 = ~n15867 | ~n16160;
  assign n13296 = ~n13295 | ~n13294;
  assign n13298 = n13297 ^ n13296;
  assign n13299 = ~n15527 | ~n13298;
  assign n13301 = ~n13300 | ~n13299;
  assign n13303 = ~n13302 & ~n13301;
  assign P2_U3223 = ~n13304 | ~n13303;
  assign n13306 = ~n15848 & ~n16199;
  assign n13305 = ~n15850 & ~n13549;
  assign n13308 = ~n13306 & ~n13305;
  assign n13307 = ~P2_REG2_REG_9__SCAN_IN | ~n15488;
  assign n13316 = ~n13308 | ~n13307;
  assign n13490 = n16176 ^ n13309;
  assign n13314 = ~n15847 | ~n13490;
  assign n13311 = ~n15888;
  assign n13310 = ~n15890;
  assign n13313 = ~n14078 | ~n13495;
  assign n13315 = ~n13314 | ~n13313;
  assign n13326 = ~n13316 & ~n13315;
  assign n13321 = ~n13495 | ~n10644;
  assign n13319 = ~n13642 & ~n15713;
  assign n13318 = ~n13317 & ~n16488;
  assign n13320 = ~n13319 & ~n13318;
  assign n13324 = ~n13321 | ~n13320;
  assign n13322 = n15986 ^ n15887;
  assign n13323 = ~n13322 & ~n15547;
  assign n13494 = n13324 | n13323;
  assign n13325 = ~n13494 | ~n15720;
  assign P2_U3287 = ~n13326 | ~n13325;
  assign n13328 = ~P2_DATAO_REG_29__SCAN_IN | ~n13390;
  assign n13327 = ~P2_U3966 | ~n16427;
  assign P2_U3581 = ~n13328 | ~n13327;
  assign n13333 = ~n13334 | ~n14582;
  assign n13331 = ~n13329 & ~P1_U3084;
  assign n13330 = n14388 & P2_DATAO_REG_21__SCAN_IN;
  assign n13332 = ~n13331 & ~n13330;
  assign P1_U3332 = ~n13333 | ~n13332;
  assign n13339 = ~n13334 | ~n11059;
  assign n13337 = ~n16031 & ~P2_U3152;
  assign n13336 = ~n14962 & ~n13335;
  assign n13338 = ~n13337 & ~n13336;
  assign P2_U3337 = ~n13339 | ~n13338;
  assign n13341 = ~n13589 | ~n13340;
  assign n16991 = ~n16624;
  assign n13348 = ~n13407 & ~n15608;
  assign n13344 = ~n13595 & ~n15763;
  assign n13343 = ~n15766 & ~n13473;
  assign n13346 = ~n13344 & ~n13343;
  assign n13345 = ~P1_REG2_REG_10__SCAN_IN | ~n15218;
  assign n13347 = ~n13346 | ~n13345;
  assign n13363 = ~n13348 & ~n13347;
  assign n13349 = ~n16628 | ~n13474;
  assign n13351 = ~n13350 & ~n16934;
  assign n16910 = ~n16628 & ~n13474;
  assign n13580 = ~n13351 & ~n16910;
  assign n13352 = ~n16624 ^ n13580;
  assign n13356 = ~n13352 | ~n10774;
  assign n13354 = ~n16629 & ~n15594;
  assign n13353 = ~n13598 & ~n15595;
  assign n13355 = ~n13354 & ~n13353;
  assign n13357 = ~n13407 & ~n15404;
  assign n13610 = ~n16628 | ~n13359;
  assign n13408 = n13611 ^ n13610;
  assign n13360 = ~n13408 | ~n14237;
  assign n13361 = ~n13414 | ~n13360;
  assign n13362 = ~n13361 | ~n15745;
  assign P1_U3281 = ~n13363 | ~n13362;
  assign n13382 = ~P1_REG1_REG_7__SCAN_IN | ~n15806;
  assign n13434 = ~n13365 ^ n13364;
  assign n13369 = ~n13434 | ~n15791;
  assign n13367 = ~n13424 & ~n15422;
  assign n13426 = ~n13366 & ~n15595;
  assign n13368 = ~n13367 & ~n13426;
  assign n13380 = n13369 & n13368;
  assign n13423 = ~n16983 ^ n13370;
  assign n13378 = ~n13423 & ~n15619;
  assign n13373 = ~n13423 & ~n15404;
  assign n13372 = ~n13371 & ~n15594;
  assign n13377 = ~n13373 & ~n13372;
  assign n13375 = ~n16606 ^ n13374;
  assign n13376 = ~n13375 | ~n10774;
  assign n13379 = ~n13378 & ~n13425;
  assign n13381 = ~n15804 | ~n13383;
  assign P1_U3530 = ~n13382 | ~n13381;
  assign n13385 = ~P1_REG0_REG_7__SCAN_IN | ~n15801;
  assign n13384 = ~n15800 | ~n13383;
  assign P1_U3475 = ~n13385 | ~n13384;
  assign n13389 = ~n13387 & ~n13386;
  assign ADD_1071_U56 = n13389 ^ n13388;
  assign n13392 = ~P2_DATAO_REG_28__SCAN_IN | ~n13390;
  assign n13391 = ~P2_U3966 | ~n15868;
  assign P2_U3580 = ~n13392 | ~n13391;
  assign n13403 = ~P2_REG0_REG_8__SCAN_IN | ~n16511;
  assign n13394 = ~n16160 | ~n16502;
  assign n13398 = ~n13394 | ~n13393;
  assign n13400 = ~n13399 | ~n14993;
  assign n13402 = ~n16510 | ~n13404;
  assign P2_U3475 = ~n13403 | ~n13402;
  assign n13406 = ~P2_REG1_REG_8__SCAN_IN | ~n16516;
  assign n13405 = ~n16514 | ~n13404;
  assign P2_U3528 = ~n13406 | ~n13405;
  assign n13416 = ~P1_REG0_REG_10__SCAN_IN | ~n15801;
  assign n13412 = ~n13407 & ~n15619;
  assign n13410 = ~n13408 | ~n15791;
  assign n13409 = ~n13611 | ~n15793;
  assign n13411 = ~n13410 | ~n13409;
  assign n13413 = ~n13412 & ~n13411;
  assign n13415 = ~n15800 | ~n13417;
  assign P1_U3484 = ~n13416 | ~n13415;
  assign n13419 = ~P1_REG1_REG_10__SCAN_IN | ~n15806;
  assign n13418 = ~n15804 | ~n13417;
  assign P1_U3533 = ~n13419 | ~n13418;
  assign n13422 = ~n15218 | ~P1_REG2_REG_7__SCAN_IN;
  assign n13421 = ~n13420 | ~n15407;
  assign n13433 = ~n13422 | ~n13421;
  assign n13431 = n13423 | n15608;
  assign n13429 = ~n15763 & ~n13424;
  assign n13427 = ~n13426 & ~n13425;
  assign n13428 = ~n15218 & ~n13427;
  assign n13430 = ~n13429 & ~n13428;
  assign n13432 = ~n13431 | ~n13430;
  assign n13436 = ~n13433 & ~n13432;
  assign n13435 = ~n15762 | ~n13434;
  assign P1_U3284 = ~n13436 | ~n13435;
  assign n13447 = ~P2_REG0_REG_7__SCAN_IN | ~n16511;
  assign n13440 = ~n13437 | ~n16500;
  assign n13439 = ~n13438 | ~n14993;
  assign n13441 = ~n13440 | ~n13439;
  assign n13445 = ~n13442 & ~n13441;
  assign n13444 = ~n13443 | ~n16502;
  assign n13446 = ~n16510 | ~n13448;
  assign P2_U3472 = ~n13447 | ~n13446;
  assign n13450 = ~P2_REG1_REG_7__SCAN_IN | ~n16516;
  assign n13449 = ~n16514 | ~n13448;
  assign P2_U3527 = ~n13450 | ~n13449;
  assign n13454 = ~n13458 & ~P1_REG2_REG_14__SCAN_IN;
  assign n13457 = ~n13455 & ~P1_REG2_REG_15__SCAN_IN;
  assign n13456 = ~n13772 | ~n14325;
  assign n13470 = ~n13457 & ~n13456;
  assign n13460 = ~n13458 | ~P1_REG1_REG_14__SCAN_IN;
  assign n13464 = ~n13462 & ~P1_REG1_REG_15__SCAN_IN;
  assign n13463 = ~n14333 | ~n13760;
  assign n13466 = ~n13464 & ~n13463;
  assign n13468 = ~n13466 & ~n13465;
  assign n13467 = ~n14837 | ~n13771;
  assign n13469 = ~n13468 | ~n13467;
  assign n13472 = ~n13470 & ~n13469;
  assign n13471 = ~n14842 | ~P1_ADDR_REG_15__SCAN_IN;
  assign P1_U3256 = ~n13472 | ~n13471;
  assign n13478 = ~n13473 & ~n14796;
  assign n13476 = ~n13611 | ~n15578;
  assign n13475 = ~n15696 | ~n13474;
  assign n13477 = ~n13476 | ~n13475;
  assign n13480 = ~n13478 & ~n13477;
  assign n13482 = ~n13480 | ~n13479;
  assign n13481 = ~n15689 & ~n13598;
  assign n13489 = ~n13482 & ~n13481;
  assign n13487 = ~n13486 ^ n13485;
  assign n13488 = ~n13487 | ~n10132;
  assign P1_U3215 = ~n13489 | ~n13488;
  assign n13499 = ~P2_REG1_REG_9__SCAN_IN | ~n16516;
  assign n13492 = ~n13490 | ~n16500;
  assign n13491 = ~n16176 | ~n16502;
  assign n13493 = ~n13492 | ~n13491;
  assign P2_U3529 = ~n13499 | ~n13498;
  assign n13502 = ~P2_REG0_REG_9__SCAN_IN | ~n16511;
  assign P2_U3478 = ~n13502 | ~n13501;
  assign n13505 = ~n13508 & ~n14384;
  assign n17093 = ~n13503;
  assign n13504 = ~n17093 & ~P1_U3084;
  assign n13507 = ~n13505 & ~n13504;
  assign n13506 = ~n14388 | ~P2_DATAO_REG_22__SCAN_IN;
  assign P1_U3331 = ~n13507 | ~n13506;
  assign n13510 = ~n13508 & ~n14094;
  assign n13509 = ~n16491 & ~P2_U3152;
  assign n13512 = ~n13510 & ~n13509;
  assign n13511 = ~n14577 | ~P1_DATAO_REG_22__SCAN_IN;
  assign P2_U3336 = ~n13512 | ~n13511;
  assign n13514 = ~n15532 | ~n16177;
  assign n13516 = ~n13514 | ~n13513;
  assign n13515 = ~n15535 & ~n16192;
  assign n13527 = ~n13516 & ~n13515;
  assign n13525 = ~n13683 & ~n15865;
  assign n13523 = ~n15867 | ~n16205;
  assign n13519 = ~n13518 | ~n13517;
  assign n13521 = n13520 ^ n13519;
  assign n13522 = ~n15527 | ~n13521;
  assign n13526 = ~n13525 & ~n13524;
  assign P2_U3219 = ~n13527 | ~n13526;
  assign n13528 = ~n14864 | ~P2_ADDR_REG_15__SCAN_IN;
  assign n13544 = ~n13529 | ~n13528;
  assign n13533 = ~P2_REG1_REG_14__SCAN_IN & ~n13535;
  assign n13534 = ~P2_REG1_REG_15__SCAN_IN ^ n13875;
  assign n13542 = ~n13534 | ~n11932;
  assign n13539 = ~P2_REG2_REG_14__SCAN_IN & ~n13535;
  assign n13540 = ~P2_REG2_REG_15__SCAN_IN ^ n13865;
  assign n13541 = ~n13540 | ~n14882;
  assign n13546 = ~n13544 & ~n13543;
  assign n13545 = ~n14887 | ~n13874;
  assign P2_U3260 = ~n13546 | ~n13545;
  assign ADD_1071_U55 = ~n13548 ^ n13547;
  assign n13562 = ~n15865 & ~n13549;
  assign n13551 = ~n15532 | ~n16161;
  assign n13553 = ~n13551 | ~n13550;
  assign n13552 = ~n15535 & ~n13642;
  assign n13560 = ~n13553 & ~n13552;
  assign n13557 = n13555 | n13554;
  assign n13558 = ~n13557 | ~n13556;
  assign n13559 = ~n15527 | ~n13558;
  assign n13564 = ~n13562 & ~n13561;
  assign n13563 = ~n15867 | ~n16176;
  assign P2_U3233 = ~n13564 | ~n13563;
  assign n13579 = ~n14853 | ~n13842;
  assign n13567 = ~n13566 | ~n13565;
  assign n13569 = n13568 ^ n13567;
  assign n13577 = ~n13569 & ~n17147;
  assign n13571 = ~n17136 & ~n13594;
  assign n13573 = n13571 | n13570;
  assign n13572 = ~n15689 & ~n13961;
  assign n13575 = ~n13573 & ~n13572;
  assign n13574 = ~n15578 | ~n13837;
  assign n13576 = ~n13575 | ~n13574;
  assign n13578 = ~n13577 & ~n13576;
  assign P1_U3234 = ~n13579 | ~n13578;
  assign n13781 = ~n13581 | ~n16935;
  assign n13582 = ~n13781 | ~n16914;
  assign n13585 = ~n14146 & ~n15595;
  assign n13584 = ~n13598 & ~n15594;
  assign n13586 = ~n13585 & ~n13584;
  assign n13591 = ~n13611 | ~n13783;
  assign n13789 = ~n13597 | ~n13596;
  assign n13788 = ~n13789 | ~n16989;
  assign n13609 = ~n15218 & ~n13664;
  assign n13605 = ~n13657 & ~n15608;
  assign n13603 = ~n13973 | ~n15313;
  assign n13602 = ~n15218 | ~P1_REG2_REG_12__SCAN_IN;
  assign n13604 = ~n13603 | ~n13602;
  assign n13607 = ~n13605 & ~n13604;
  assign n13606 = ~n13811 | ~n15407;
  assign n13613 = ~n13609 & ~n13608;
  assign n13793 = ~n13611 & ~n13610;
  assign n13658 = n13974 ^ n13973;
  assign n13612 = ~n13658 | ~n15762;
  assign P1_U3279 = ~n13613 | ~n13612;
  assign n13615 = ~n13614;
  assign n13617 = ~n15988;
  assign n13624 = n13670 | n14769;
  assign n13622 = ~n16226 & ~n15713;
  assign n13621 = ~n13642 & ~n16488;
  assign n13623 = ~n13622 & ~n13621;
  assign n13636 = ~n15488 & ~n13677;
  assign n13632 = ~n15845 & ~n13670;
  assign n13630 = ~n15566 | ~n16188;
  assign n13629 = ~n15725 | ~n13654;
  assign n13631 = ~n13630 | ~n13629;
  assign n13634 = ~n13632 & ~n13631;
  assign n13633 = ~n15488 | ~P2_REG2_REG_11__SCAN_IN;
  assign n13639 = ~n13636 & ~n13635;
  assign n13671 = n13637 ^ n16188;
  assign n13638 = ~n15847 | ~n13671;
  assign P2_U3285 = ~n13639 | ~n13638;
  assign n13641 = ~n15869 | ~n16230;
  assign n13644 = ~n13641 | ~n13640;
  assign n13643 = ~n15872 & ~n13642;
  assign n13651 = ~n13644 & ~n13643;
  assign n13647 = ~n13646 | ~n13645;
  assign n13649 = n13648 ^ n13647;
  assign n13652 = ~n14448 & ~n16203;
  assign n13655 = ~n13654 | ~n15530;
  assign P2_U3238 = ~n13656 | ~n13655;
  assign n13666 = ~P1_REG0_REG_12__SCAN_IN | ~n15801;
  assign n13662 = ~n13657 & ~n15619;
  assign n13660 = ~n13658 | ~n15791;
  assign n13659 = ~n13973 | ~n15793;
  assign n13661 = ~n13660 | ~n13659;
  assign P1_U3490 = ~n13666 | ~n13665;
  assign n13669 = ~P1_REG1_REG_12__SCAN_IN | ~n15806;
  assign P1_U3535 = ~n13669 | ~n13668;
  assign n13679 = ~P2_REG0_REG_11__SCAN_IN | ~n16511;
  assign n13675 = ~n13670 & ~n16498;
  assign n13673 = ~n13671 | ~n16500;
  assign n13672 = ~n16188 | ~n16502;
  assign n13674 = ~n13673 | ~n13672;
  assign P2_U3484 = ~n13679 | ~n13678;
  assign n13682 = ~P2_REG1_REG_11__SCAN_IN | ~n16516;
  assign P2_U3531 = ~n13682 | ~n13681;
  assign n13685 = ~n15848 & ~n13738;
  assign n13684 = ~n15850 & ~n13683;
  assign n13687 = ~n13685 & ~n13684;
  assign n13686 = ~P2_REG2_REG_10__SCAN_IN | ~n15488;
  assign n13694 = ~n13687 | ~n13686;
  assign n13739 = ~n16205 ^ n13688;
  assign n13692 = ~n15847 | ~n13739;
  assign n13691 = ~n14078 | ~n13740;
  assign n13693 = ~n13692 | ~n13691;
  assign n13704 = ~n13694 & ~n13693;
  assign n13698 = ~n16177 | ~n15550;
  assign n13697 = n13696 | n15547;
  assign n13699 = ~n16192 & ~n15713;
  assign n13703 = ~n13737 | ~n15720;
  assign P2_U3286 = ~n13704 | ~n13703;
  assign n13706 = ~n14388 | ~P2_DATAO_REG_23__SCAN_IN;
  assign P1_U3330 = ~n13707 | ~n13706;
  assign n13711 = ~n14577 | ~P1_DATAO_REG_23__SCAN_IN;
  assign P2_U3335 = ~n13712 | ~n13711;
  assign n13716 = ~n14164 & ~n15850;
  assign n13714 = ~n15566 | ~n16229;
  assign n13713 = ~n15488 | ~P2_REG2_REG_12__SCAN_IN;
  assign n13736 = ~n13716 & ~n13715;
  assign n13718 = ~n15902;
  assign n13724 = n13890 & n15272;
  assign n13721 = ~n16225 & ~n13720;
  assign n13722 = ~n13721 & ~n14995;
  assign n13723 = ~n13893 & ~n16472;
  assign n13733 = ~n13724 & ~n13723;
  assign n13726 = ~n16192 & ~n16488;
  assign n13725 = ~n14167 & ~n15713;
  assign n13727 = ~n13726 & ~n13725;
  assign P2_U3284 = ~n13736 | ~n13735;
  assign n13748 = ~P2_REG0_REG_10__SCAN_IN | ~n16511;
  assign n13744 = ~n13738 & ~n15451;
  assign n13742 = ~n16500 | ~n13739;
  assign n13741 = ~n14993 | ~n13740;
  assign P2_U3481 = ~n13748 | ~n13747;
  assign n13751 = ~P2_REG1_REG_10__SCAN_IN | ~n16516;
  assign P2_U3530 = ~n13751 | ~n13750;
  assign n13755 = ~n13753 & ~P1_U3084;
  assign n13754 = n14388 & P2_DATAO_REG_24__SCAN_IN;
  assign n13756 = ~n13755 & ~n13754;
  assign P1_U3329 = ~n13757 | ~n13756;
  assign n14528 = ~P1_REG3_REG_16__SCAN_IN | ~P1_U3084;
  assign n13758 = ~n14837 | ~n14328;
  assign n13769 = ~n14528 | ~n13758;
  assign n13767 = ~n14842 | ~P1_ADDR_REG_16__SCAN_IN;
  assign n13764 = ~P1_REG1_REG_16__SCAN_IN ^ n13774;
  assign n13762 = ~n13763 & ~n13764;
  assign n13765 = ~n13762 & ~n14833;
  assign n13766 = ~n13765 | ~n14329;
  assign n13768 = ~n13767 | ~n13766;
  assign n13780 = ~n13769 & ~n13768;
  assign n13777 = ~P1_REG2_REG_16__SCAN_IN ^ n13774;
  assign n13775 = ~n13776 & ~n13777;
  assign n13778 = ~n13775 & ~n14825;
  assign n13779 = ~n13778 | ~n14321;
  assign P1_U3257 = ~n13780 | ~n13779;
  assign n13801 = ~P1_REG1_REG_11__SCAN_IN | ~n15806;
  assign n13785 = ~n15636 | ~n13855;
  assign n13784 = ~n17091 | ~n13783;
  assign n13786 = ~n13785 | ~n13784;
  assign n13791 = ~n13788;
  assign n13790 = ~n13789 & ~n16989;
  assign n13798 = ~n13830 & ~n15789;
  assign n13794 = ~n13793 & ~n13792;
  assign n13795 = ~n13794 & ~n15185;
  assign n13831 = ~n13795 | ~n13974;
  assign n13796 = ~n13837 | ~n15793;
  assign n13797 = ~n13831 | ~n13796;
  assign n13799 = ~n13798 & ~n13797;
  assign P1_U3534 = ~n13801 | ~n13800;
  assign n13804 = ~P1_REG0_REG_11__SCAN_IN | ~n15801;
  assign P1_U3487 = ~n13804 | ~n13803;
  assign n13807 = ~n13806 & ~P2_U3152;
  assign n13809 = ~n14577 | ~P1_DATAO_REG_24__SCAN_IN;
  assign P2_U3334 = ~n13810 | ~n13809;
  assign n13828 = ~n14853 | ~n13811;
  assign n13816 = ~n13812 & ~n13845;
  assign n13813 = ~n13846;
  assign n13814 = ~n13813 & ~n13845;
  assign n13815 = ~n9042 & ~n13814;
  assign n13824 = ~n13973 | ~n15578;
  assign n13822 = ~n15689 & ~n14146;
  assign n13820 = ~n15696 | ~n13818;
  assign n13821 = ~n13820 | ~n13819;
  assign n13823 = ~n13822 & ~n13821;
  assign n13825 = ~n13824 | ~n13823;
  assign P1_U3222 = ~n13828 | ~n13827;
  assign n13835 = ~n13830 & ~n13829;
  assign n13833 = n13831 | n14836;
  assign n13836 = ~n13835 & ~n13834;
  assign n13841 = ~n15218 & ~n13836;
  assign n13839 = ~n13837 | ~n15313;
  assign n13838 = ~n15218 | ~P1_REG2_REG_11__SCAN_IN;
  assign n13840 = ~n13839 | ~n13838;
  assign n13843 = ~n13842 | ~n15407;
  assign P1_U3280 = ~n13844 | ~n13843;
  assign n13863 = ~n14853 | ~n13979;
  assign n13849 = ~n9042 & ~n13845;
  assign n13848 = ~n13847 | ~n13846;
  assign n13850 = ~n13849 & ~n13848;
  assign n13851 = ~n13850 & ~n17147;
  assign n13859 = ~n14159 & ~n17126;
  assign n13854 = ~n15689 & ~n14151;
  assign n13857 = ~n13854 & ~n13853;
  assign n13856 = ~n15696 | ~n13855;
  assign n13858 = ~n13857 | ~n13856;
  assign n13860 = ~n13859 & ~n13858;
  assign P1_U3232 = ~n13863 | ~n13862;
  assign n13868 = ~P2_REG2_REG_16__SCAN_IN;
  assign n13870 = ~n14425 ^ n13868;
  assign n13872 = ~n13869 & ~n13870;
  assign n13871 = ~n14882 | ~n14426;
  assign n13887 = ~n13872 & ~n13871;
  assign n13879 = P2_REG1_REG_16__SCAN_IN ^ n14425;
  assign n13881 = ~n13878 & ~n13879;
  assign n13880 = ~n14416 | ~n11932;
  assign n13883 = ~n13881 & ~n13880;
  assign n14449 = ~P2_STATE_REG_SCAN_IN & ~n13882;
  assign n13885 = ~n13883 & ~n14449;
  assign n13884 = ~n14864 | ~P2_ADDR_REG_16__SCAN_IN;
  assign n13888 = ~n14887 | ~n14425;
  assign P2_U3261 = ~n13889 | ~n13888;
  assign n13898 = ~P2_REG1_REG_12__SCAN_IN | ~n16516;
  assign n13891 = ~n16225 & ~n15451;
  assign P2_U3532 = ~n13898 | ~n13897;
  assign n13901 = ~P2_REG0_REG_12__SCAN_IN | ~n16511;
  assign P2_U3487 = ~n13901 | ~n13900;
  assign n13904 = ~n16230 | ~n15550;
  assign n13903 = ~n16248 | ~n15549;
  assign n13905 = ~n13904 | ~n13903;
  assign n13912 = ~n13911 | ~n14261;
  assign n13913 = ~n13912 | ~n16500;
  assign n13933 = n13913 | n14002;
  assign n13914 = ~n14261 | ~n16502;
  assign n13919 = ~n16516 | ~P2_REG1_REG_13__SCAN_IN;
  assign P2_U3533 = ~n13920 | ~n13919;
  assign n13922 = ~n16511 | ~P2_REG0_REG_13__SCAN_IN;
  assign P2_U3490 = ~n13923 | ~n13922;
  assign n13926 = ~n15566 | ~n14261;
  assign n13925 = ~n15725 | ~n13924;
  assign n13929 = ~n13927 & ~n15488;
  assign n13928 = ~n15720 & ~P2_REG2_REG_13__SCAN_IN;
  assign n13930 = ~n13929 & ~n13928;
  assign n13935 = ~n15845 & ~n13932;
  assign n13934 = ~n14079 & ~n13933;
  assign n13936 = ~n13935 & ~n13934;
  assign P2_U3283 = ~n13937 | ~n13936;
  assign n13939 = ~n13938 & ~P1_U3084;
  assign n13941 = ~n14388 | ~P2_DATAO_REG_25__SCAN_IN;
  assign P1_U3328 = ~n13942 | ~n13941;
  assign n13945 = ~n14962 & ~n13944;
  assign n13948 = ~n13947 | ~P2_STATE_REG_SCAN_IN;
  assign P2_U3333 = ~n13949 | ~n13948;
  assign n13951 = ~n13961 & ~n15594;
  assign n13950 = ~n14151 & ~n15595;
  assign n13959 = ~n13951 & ~n13950;
  assign n13953 = ~n13952 & ~n14144;
  assign n13956 = ~n13953 & ~n16643;
  assign n13954 = ~n16668 | ~n16666;
  assign n13964 = ~n13960 | ~n16994;
  assign n13962 = ~n13973;
  assign n13966 = ~n13964 | ~n13963;
  assign n14131 = ~n13966 | ~n13965;
  assign n13967 = n13966 | n13965;
  assign n13970 = ~n14024 | ~n14655;
  assign n13969 = ~n16668 | ~n13968;
  assign n14025 = n16668 ^ n14158;
  assign n13976 = n14025 | n15174;
  assign n13975 = ~n15218 | ~P1_REG2_REG_13__SCAN_IN;
  assign n13977 = ~n13976 | ~n13975;
  assign n13980 = ~n13979 | ~n15407;
  assign P1_U3278 = ~n13981 | ~n13980;
  assign n13987 = n13983 & n13994;
  assign n13984 = ~n13994 & ~n16251;
  assign n13990 = ~n16265 | ~n15549;
  assign n13989 = ~n13988 | ~n15550;
  assign n13991 = ~n13990 | ~n13989;
  assign n13998 = ~n15725 | ~n13997;
  assign n13999 = ~n15720 | ~n13998;
  assign n14000 = ~n15720 & ~P2_REG2_REG_14__SCAN_IN;
  assign n14009 = n14001 | n14000;
  assign n14004 = ~n15566 | ~n16247;
  assign n14003 = ~n15847 | ~n14012;
  assign n14006 = ~n15845 & ~n14011;
  assign P2_U3282 = ~n14009 | ~n14008;
  assign n14013 = ~n16247 | ~n16502;
  assign n14019 = ~n16511 | ~P2_REG0_REG_14__SCAN_IN;
  assign P2_U3493 = ~n14020 | ~n14019;
  assign n14022 = ~n16516 | ~P2_REG1_REG_14__SCAN_IN;
  assign P2_U3534 = ~n14023 | ~n14022;
  assign n14033 = ~P1_REG1_REG_13__SCAN_IN | ~n15806;
  assign n14029 = ~n14025 & ~n15185;
  assign n14027 = ~n14159 & ~n15422;
  assign n14028 = n14027 | n14026;
  assign P1_U3536 = ~n14033 | ~n14032;
  assign n14036 = ~P1_REG0_REG_13__SCAN_IN | ~n15801;
  assign P1_U3493 = ~n14036 | ~n14035;
  assign n14040 = ~n14038 & ~P1_U3084;
  assign n14039 = n14388 & P2_DATAO_REG_26__SCAN_IN;
  assign n14041 = ~n14040 & ~n14039;
  assign P1_U3327 = ~n14042 | ~n14041;
  assign n14044 = ~n15848 & ~n14447;
  assign n14043 = n15725 & n14432;
  assign n14046 = ~n14044 & ~n14043;
  assign n14045 = ~n15847 | ~n14117;
  assign n14056 = ~n16265 | ~n15550;
  assign n14055 = ~n16051 | ~n15549;
  assign n14057 = ~n14056 | ~n14055;
  assign n14059 = n15720 | P2_REG2_REG_16__SCAN_IN;
  assign P2_U3280 = ~n14062 | ~n14061;
  assign n14065 = ~n16285 & ~n15713;
  assign n14064 = ~n16244 & ~n16488;
  assign n14066 = ~n14065 & ~n14064;
  assign n14075 = ~P2_REG2_REG_15__SCAN_IN;
  assign n14076 = ~n15488 | ~n14075;
  assign n14084 = ~n14079;
  assign n14081 = ~n16266 | ~n14080;
  assign n14085 = ~n14084 | ~n14106;
  assign n14089 = ~n15566 | ~n16266;
  assign n14088 = ~n15725 | ~n14087;
  assign n14090 = ~n14089 | ~n14088;
  assign P2_U3281 = ~n14093 | ~n14092;
  assign n14097 = ~n14962 & ~n14096;
  assign n14100 = ~n14099 | ~P2_STATE_REG_SCAN_IN;
  assign P2_U3332 = ~n14101 | ~n14100;
  assign n14105 = ~n14104 & ~n15451;
  assign n14107 = n14106 | n14105;
  assign n14111 = ~n16516 | ~P2_REG1_REG_15__SCAN_IN;
  assign P2_U3535 = ~n14112 | ~n14111;
  assign n14114 = ~n16511 | ~P2_REG0_REG_15__SCAN_IN;
  assign P2_U3496 = ~n14115 | ~n14114;
  assign n14118 = ~n16280 | ~n16502;
  assign n14124 = ~n16511 | ~P2_REG0_REG_16__SCAN_IN;
  assign P2_U3499 = ~n14125 | ~n14124;
  assign n14127 = ~n16516 | ~P2_REG1_REG_16__SCAN_IN;
  assign P2_U3536 = ~n14128 | ~n14127;
  assign n14135 = ~n14133 | ~n14132;
  assign n14134 = ~n16657 | ~n16678;
  assign n14280 = ~n14135 | ~n14134;
  assign n14138 = ~n16700 & ~n15763;
  assign n14137 = ~n15766 & ~n14136;
  assign n14140 = ~n14138 & ~n14137;
  assign n14139 = ~P1_REG2_REG_15__SCAN_IN | ~n15218;
  assign n14141 = ~n14140 | ~n14139;
  assign n16671 = ~n16668 | ~n14146;
  assign n14143 = ~n16637;
  assign n16653 = ~n14144 & ~n14143;
  assign n14145 = ~n16653;
  assign n16650 = ~n16668 & ~n14146;
  assign n14265 = ~n14225 | ~n16931;
  assign n14153 = ~n14151 & ~n15594;
  assign n14152 = ~n16689 & ~n15595;
  assign n14154 = ~n14153 & ~n14152;
  assign n14295 = ~n14296 ^ n14275;
  assign n14160 = ~n14295 | ~n14237;
  assign P1_U3276 = ~n14163 | ~n14162;
  assign n14179 = ~n15865 & ~n14164;
  assign n14166 = ~n15532 | ~n16189;
  assign n14169 = ~n14166 | ~n14165;
  assign n14168 = ~n15535 & ~n14167;
  assign n14177 = ~n14169 & ~n14168;
  assign n14174 = ~n14170 & ~n14247;
  assign n14249 = ~n14171;
  assign n14172 = ~n14249 & ~n14247;
  assign n14173 = ~n14248 & ~n14172;
  assign n14180 = ~n15867 | ~n16229;
  assign P2_U3226 = ~n14181 | ~n14180;
  assign n14196 = n14796 | n14218;
  assign n14185 = ~n14183 | ~n14182;
  assign n14192 = ~n16657 | ~n15578;
  assign n14190 = ~n15689 & ~n16701;
  assign n14188 = ~n15696 | ~n16666;
  assign n14189 = ~n14188 | ~n14187;
  assign n14191 = ~n14190 & ~n14189;
  assign n14193 = ~n14192 | ~n14191;
  assign P1_U3213 = ~n14196 | ~n14195;
  assign n14200 = ~n16487 & ~P2_U3152;
  assign n14199 = ~n14962 & ~n14198;
  assign n14201 = ~n14200 & ~n14199;
  assign P2_U3331 = ~n14202 | ~n14201;
  assign n14210 = ~n16516 | ~P2_REG1_REG_17__SCAN_IN;
  assign P2_U3537 = ~n14211 | ~n14210;
  assign n14213 = ~n16511 | ~P2_REG0_REG_17__SCAN_IN;
  assign P2_U3502 = ~n14214 | ~n14213;
  assign n14224 = ~n14391 & ~n15608;
  assign n14220 = ~n14217 & ~n15763;
  assign n14219 = ~n15766 & ~n14218;
  assign n14222 = ~n14220 & ~n14219;
  assign n14221 = ~P1_REG2_REG_14__SCAN_IN | ~n15218;
  assign n14223 = ~n14222 | ~n14221;
  assign n14231 = ~n16701 & ~n15595;
  assign n14232 = ~n16666 | ~n17091;
  assign n14392 = n16657 ^ n14236;
  assign n14238 = ~n14392 | ~n14237;
  assign n14240 = ~n14239 | ~n15745;
  assign P1_U3277 = ~n14241 | ~n14240;
  assign n14260 = ~n15865 & ~n14242;
  assign n14244 = ~n15532 | ~n16230;
  assign n14246 = ~n14244 | ~n14243;
  assign n14245 = ~n15535 & ~n16244;
  assign n14258 = ~n14246 & ~n14245;
  assign n14250 = ~n14248 & ~n14247;
  assign n14253 = ~n14251;
  assign n14254 = ~n14253 | ~n14252;
  assign n14262 = ~n15867 | ~n14261;
  assign P2_U3236 = ~n14263 | ~n14262;
  assign n14346 = ~n14265 | ~n16922;
  assign n14268 = ~n14266 | ~n16884;
  assign n14286 = ~n14267 & ~n16880;
  assign n14269 = n14268 | n14286;
  assign n14272 = ~n16544 & ~n15595;
  assign n14271 = ~n16689 & ~n15594;
  assign n14273 = ~n14272 & ~n14271;
  assign n14276 = ~n16716 | ~n15793;
  assign n14282 = ~n14280 | ~n14279;
  assign n14281 = ~n14296 | ~n14527;
  assign n14356 = ~n14282 | ~n14281;
  assign n14285 = ~n14356 | ~n14283;
  assign n14481 = ~n14285 | ~n14284;
  assign n14289 = ~n15806 | ~P1_REG1_REG_17__SCAN_IN;
  assign P1_U3540 = ~n14290 | ~n14289;
  assign n14292 = ~n15801 | ~P1_REG0_REG_17__SCAN_IN;
  assign P1_U3505 = ~n14293 | ~n14292;
  assign n14304 = ~P1_REG0_REG_15__SCAN_IN | ~n15801;
  assign n14298 = ~n14295 | ~n15791;
  assign n14297 = ~n14296 | ~n15793;
  assign P1_U3499 = ~n14304 | ~n14303;
  assign n14307 = ~P1_REG1_REG_15__SCAN_IN | ~n15806;
  assign P1_U3538 = ~n14307 | ~n14306;
  assign n14309 = ~n15745 & ~P1_REG2_REG_17__SCAN_IN;
  assign n14315 = ~n14311 | ~n15762;
  assign n14313 = ~n16712 & ~n15763;
  assign n14312 = n15407 & n14544;
  assign n14314 = ~n14313 & ~n14312;
  assign P1_U3274 = ~n14320 | ~n14319;
  assign n14324 = P1_REG2_REG_17__SCAN_IN ^ n14627;
  assign n14322 = ~n14328 | ~P1_REG2_REG_16__SCAN_IN;
  assign n14327 = ~n14324 & ~n14323;
  assign n14326 = ~n14628 | ~n14325;
  assign n14341 = ~n14327 & ~n14326;
  assign n14332 = P1_REG1_REG_17__SCAN_IN ^ n14627;
  assign n14330 = ~n14328 | ~P1_REG1_REG_16__SCAN_IN;
  assign n14335 = ~n14332 & ~n14331;
  assign n14334 = ~n14333 | ~n14617;
  assign n14337 = ~n14335 & ~n14334;
  assign n14546 = ~P1_STATE_REG_SCAN_IN & ~n14336;
  assign n14339 = ~n14337 & ~n14546;
  assign n14338 = ~n14837 | ~n14627;
  assign n14342 = ~n14842 | ~P1_ADDR_REG_17__SCAN_IN;
  assign P1_U3258 = ~n14343 | ~n14342;
  assign n14345 = ~n14344;
  assign n14351 = ~n16713 & ~n15595;
  assign n14350 = ~n16701 & ~n15594;
  assign n14352 = ~n14351 & ~n14350;
  assign n14361 = ~n14378 | ~n15745;
  assign n14359 = ~P1_REG2_REG_16__SCAN_IN;
  assign n14360 = ~n15218 | ~n14359;
  assign n14372 = n16692 ^ n14362;
  assign n14366 = ~n14372 | ~n15762;
  assign n14364 = ~n16687 & ~n15763;
  assign n14363 = ~n15766 & ~n14536;
  assign n14365 = ~n14364 & ~n14363;
  assign n14367 = ~n14366 | ~n14365;
  assign P1_U3275 = ~n14370 | ~n14369;
  assign n14374 = ~n14372 | ~n15791;
  assign n14373 = ~n16692 | ~n15793;
  assign n14379 = ~n15801 | ~P1_REG0_REG_16__SCAN_IN;
  assign P1_U3502 = ~n14380 | ~n14379;
  assign n14382 = ~n15806 | ~P1_REG1_REG_16__SCAN_IN;
  assign P1_U3539 = ~n14383 | ~n14382;
  assign n14389 = ~n14388 | ~P2_DATAO_REG_27__SCAN_IN;
  assign P1_U3326 = ~n14390 | ~n14389;
  assign n14400 = ~P1_REG0_REG_14__SCAN_IN | ~n15801;
  assign n14394 = ~n14392 | ~n15791;
  assign n14393 = ~n16657 | ~n15793;
  assign P1_U3496 = ~n14400 | ~n14399;
  assign n14403 = ~P1_REG1_REG_14__SCAN_IN | ~n15806;
  assign P1_U3537 = ~n14403 | ~n14402;
  assign n14406 = ~n14404 & ~P2_U3152;
  assign n14405 = n14577 & P1_DATAO_REG_28__SCAN_IN;
  assign n14407 = ~n14406 & ~n14405;
  assign P2_U3330 = ~n14408 | ~n14407;
  assign n14410 = ~n14585 & ~n14409;
  assign n14412 = ~n14411 & ~n14410;
  assign P1_U3325 = ~n14413 | ~n14412;
  assign n14414 = ~n14864 | ~P2_ADDR_REG_17__SCAN_IN;
  assign n14423 = ~n14415 | ~n14414;
  assign n14559 = ~P2_REG1_REG_17__SCAN_IN & ~n14424;
  assign n14558 = P2_REG1_REG_17__SCAN_IN & n14424;
  assign n14418 = ~n14559 & ~n14558;
  assign n14417 = ~P2_REG1_REG_16__SCAN_IN | ~n14425;
  assign n14419 = n14418 ^ n14557;
  assign n14420 = ~n14887 | ~n14424;
  assign n14431 = ~n14423 & ~n14422;
  assign n14564 = ~P2_REG2_REG_17__SCAN_IN & ~n14424;
  assign n14563 = P2_REG2_REG_17__SCAN_IN & n14424;
  assign n14428 = ~n14564 & ~n14563;
  assign n14427 = ~P2_REG2_REG_16__SCAN_IN | ~n14425;
  assign n14429 = n14428 ^ n14562;
  assign n14430 = ~n14882 | ~n14429;
  assign P2_U3262 = ~n14431 | ~n14430;
  assign n14446 = ~n15530 | ~n14432;
  assign n14438 = ~n14437;
  assign n14441 = ~n14439 | ~n14438;
  assign n14454 = ~n14448 & ~n14447;
  assign n14450 = ~n15535 & ~n16054;
  assign n14452 = ~n14450 & ~n14449;
  assign n14451 = ~n15532 | ~n16265;
  assign n14453 = ~n14452 | ~n14451;
  assign n14455 = ~n14454 & ~n14453;
  assign P2_U3228 = ~n14456 | ~n14455;
  assign n14460 = n14458 | n14995;
  assign n14465 = ~n16511 | ~P2_REG0_REG_18__SCAN_IN;
  assign P2_U3505 = ~n14466 | ~n14465;
  assign n14468 = ~n16516 | ~P2_REG1_REG_18__SCAN_IN;
  assign P2_U3538 = ~n14469 | ~n14468;
  assign n14473 = ~n16531 & ~n15595;
  assign n14472 = ~n16713 & ~n15594;
  assign n14474 = ~n14473 & ~n14472;
  assign n14477 = ~n14797 | ~n15793;
  assign n14483 = ~n14481 | ~n14480;
  assign n14604 = ~n14483 | ~n14482;
  assign n14487 = ~n15806 | ~P1_REG1_REG_18__SCAN_IN;
  assign P1_U3541 = ~n14488 | ~n14487;
  assign n14490 = ~n15801 | ~P1_REG0_REG_18__SCAN_IN;
  assign P1_U3508 = ~n14491 | ~n14490;
  assign n14493 = ~n15745 & ~P1_REG2_REG_18__SCAN_IN;
  assign n14499 = ~n14495 | ~n15762;
  assign n14497 = ~n16728 & ~n15763;
  assign n14496 = ~n14795 & ~n15766;
  assign n14498 = ~n14497 & ~n14496;
  assign P1_U3273 = ~n14504 | ~n14503;
  assign n14514 = n15530 & n14505;
  assign n14507 = ~n15869 | ~n14506;
  assign n14556 = ~P2_REG3_REG_18__SCAN_IN | ~P2_U3152;
  assign n14509 = ~n14507 | ~n14556;
  assign n14508 = ~n15872 & ~n16054;
  assign n14512 = ~n14509 & ~n14508;
  assign n14511 = ~n15867 | ~n14510;
  assign n14513 = ~n14512 | ~n14511;
  assign n14521 = ~n14514 & ~n14513;
  assign P2_U3240 = ~n14521 | ~n14520;
  assign n14533 = ~n16692 | ~n15578;
  assign n14531 = ~n15689 & ~n16713;
  assign n14529 = ~n15696 | ~n14527;
  assign n14530 = ~n14529 | ~n14528;
  assign n14532 = ~n14531 & ~n14530;
  assign n14534 = ~n14533 | ~n14532;
  assign n14537 = n14796 | n14536;
  assign P1_U3224 = ~n14538 | ~n14537;
  assign n14552 = ~n16712 & ~n17126;
  assign n14550 = ~n14605 | ~n17132;
  assign n14548 = ~n17136 & ~n16689;
  assign n14545 = n14853 & n14544;
  assign n14547 = n14546 | n14545;
  assign n14549 = ~n14548 & ~n14547;
  assign n14551 = ~n14550 | ~n14549;
  assign n14553 = ~n14552 & ~n14551;
  assign P1_U3226 = ~n14554 | ~n14553;
  assign n14555 = ~n14864 | ~P2_ADDR_REG_18__SCAN_IN;
  assign n14571 = ~n14556 | ~n14555;
  assign n14867 = P2_REG1_REG_18__SCAN_IN ^ n14566;
  assign n14874 = P2_REG2_REG_18__SCAN_IN ^ n14566;
  assign n14572 = ~n14887 | ~n14876;
  assign P2_U3263 = ~n14573 | ~n14572;
  assign n14579 = ~n14576 & ~P2_U3152;
  assign n14578 = n14577 & P1_DATAO_REG_29__SCAN_IN;
  assign n14580 = ~n14579 & ~n14578;
  assign P2_U3329 = ~n14581 | ~n14580;
  assign n14587 = ~n14583 & ~P1_U3084;
  assign n14584 = ~P2_DATAO_REG_29__SCAN_IN;
  assign n14586 = ~n14585 & ~n14584;
  assign n14588 = ~n14587 & ~n14586;
  assign P1_U3324 = ~n14589 | ~n14588;
  assign n14668 = ~n14590 & ~n16881;
  assign n14595 = ~n14850 & ~n15595;
  assign n14594 = ~n16544 & ~n15594;
  assign n14596 = ~n14595 & ~n14594;
  assign n14602 = ~n16548 | ~n15793;
  assign n14607 = ~n14604 | ~n16540;
  assign n14683 = ~n14607 | ~n14606;
  assign n14611 = ~n15801 | ~P1_REG0_REG_19__SCAN_IN;
  assign P1_U3510 = ~n14612 | ~n14611;
  assign n14614 = ~n15806 | ~P1_REG1_REG_19__SCAN_IN;
  assign P1_U3542 = ~n14615 | ~n14614;
  assign n14798 = ~P1_REG3_REG_18__SCAN_IN | ~P1_U3084;
  assign n14616 = ~n14837 | ~n14828;
  assign n14626 = ~n14798 | ~n14616;
  assign n14624 = ~n14842 | ~P1_ADDR_REG_18__SCAN_IN;
  assign n14618 = ~P1_REG1_REG_17__SCAN_IN | ~n14627;
  assign n14630 = ~n14828;
  assign n14621 = ~P1_REG1_REG_18__SCAN_IN ^ n14630;
  assign n14619 = ~n14620 & ~n14621;
  assign n14622 = ~n14619 & ~n14833;
  assign n14636 = ~n14626 & ~n14625;
  assign n14629 = ~P1_REG2_REG_17__SCAN_IN | ~n14627;
  assign n14633 = ~P1_REG2_REG_18__SCAN_IN ^ n14630;
  assign n14631 = ~n14632 & ~n14633;
  assign n14634 = ~n14631 & ~n14825;
  assign n14635 = ~n14634 | ~n14822;
  assign P1_U3259 = ~n14636 | ~n14635;
  assign n14648 = n15530 & n14640;
  assign n14641 = ~n15869 | ~n16299;
  assign n14866 = ~P2_REG3_REG_19__SCAN_IN | ~P2_U3152;
  assign n14644 = ~n14641 | ~n14866;
  assign n14643 = ~n15872 & ~n14642;
  assign n14646 = ~n14644 & ~n14643;
  assign n14645 = ~n15867 | ~n15914;
  assign n14649 = ~n14648 & ~n14647;
  assign P2_U3221 = ~n14650 | ~n14649;
  assign n14652 = n14651 | n14836;
  assign n14653 = ~n14652 | ~n15745;
  assign n14660 = ~n15218 | ~n14659;
  assign n14663 = ~n16548 | ~n15313;
  assign n14662 = ~n14852 | ~n15407;
  assign P1_U3272 = n14665 | n14664;
  assign n14730 = ~n14669 & ~n17005;
  assign n14672 = ~n14924 & ~n15595;
  assign n14671 = ~n16531 & ~n15594;
  assign n14673 = ~n14672 & ~n14671;
  assign n14675 = ~n15745 & ~P1_REG2_REG_20__SCAN_IN;
  assign n14678 = ~n14948 & ~n15763;
  assign n14677 = ~n14947 & ~n15766;
  assign n14679 = ~n14678 & ~n14677;
  assign n14685 = ~n14683 | ~n16537;
  assign n14747 = ~n14685 | ~n14684;
  assign P1_U3271 = ~n14687 | ~n14686;
  assign n14696 = ~n15806 | ~P1_REG1_REG_20__SCAN_IN;
  assign P1_U3543 = ~n14697 | ~n14696;
  assign n14699 = ~n15801 | ~P1_REG0_REG_20__SCAN_IN;
  assign P1_U3511 = ~n14700 | ~n14699;
  assign n14710 = ~n16516 | ~P2_REG1_REG_19__SCAN_IN;
  assign P2_U3539 = ~n14711 | ~n14710;
  assign n14713 = ~n16511 | ~P2_REG0_REG_19__SCAN_IN;
  assign P2_U3507 = ~n14714 | ~n14713;
  assign n14727 = n15530 & n14780;
  assign n14721 = ~n15869 | ~n16322;
  assign n14720 = ~P2_REG3_REG_20__SCAN_IN | ~P2_U3152;
  assign n14723 = ~n14721 | ~n14720;
  assign n14722 = ~n15872 & ~n15913;
  assign n14725 = ~n14723 & ~n14722;
  assign P2_U3235 = ~n14729 | ~n14728;
  assign n16877 = ~n15087 & ~n16739;
  assign n17012 = ~n16867 & ~n16877;
  assign n14907 = ~n14731 | ~n16875;
  assign n14734 = ~n14906 & ~n15595;
  assign n14733 = ~n14850 & ~n15594;
  assign n14735 = ~n14734 & ~n14733;
  assign n14737 = ~n15745 & ~P1_REG2_REG_21__SCAN_IN;
  assign n14741 = ~n15087 & ~n15763;
  assign n14740 = ~n15085 & ~n15766;
  assign n14742 = ~n14741 & ~n14740;
  assign n14750 = ~n14747 | ~n14746;
  assign n14923 = ~n14750 | ~n14749;
  assign P1_U3270 = ~n14752 | ~n14751;
  assign n14755 = ~n14753 | ~n15791;
  assign n14761 = ~n15806 | ~P1_REG1_REG_21__SCAN_IN;
  assign P1_U3544 = ~n14762 | ~n14761;
  assign n14764 = ~n15801 | ~P1_REG0_REG_21__SCAN_IN;
  assign P1_U3512 = ~n14765 | ~n14764;
  assign n14773 = ~n15913 & ~n16488;
  assign n14772 = ~n15031 & ~n15713;
  assign n14774 = ~n14773 & ~n14772;
  assign n14778 = n15720 | P2_REG2_REG_20__SCAN_IN;
  assign n14782 = ~n15848 & ~n16302;
  assign n14781 = n15725 & n14780;
  assign n14785 = ~n14782 & ~n14781;
  assign P2_U3276 = ~n14789 | ~n14788;
  assign n14793 = ~n14791 | ~n14790;
  assign n14805 = ~n14796 & ~n14795;
  assign n14803 = ~n14797 | ~n15578;
  assign n14801 = ~n16531 & ~n15689;
  assign n14799 = ~n15696 | ~n16717;
  assign n14800 = ~n14799 | ~n14798;
  assign n14802 = ~n14801 & ~n14800;
  assign n14806 = ~n14805 & ~n14804;
  assign P1_U3236 = ~n14807 | ~n14806;
  assign n14816 = ~n16511 | ~P2_REG0_REG_20__SCAN_IN;
  assign P2_U3508 = ~n14817 | ~n14816;
  assign n14819 = ~n16516 | ~P2_REG1_REG_20__SCAN_IN;
  assign P2_U3540 = ~n14820 | ~n14819;
  assign n14824 = n17072 ^ P1_REG2_REG_19__SCAN_IN;
  assign n14821 = ~n14828 | ~P1_REG2_REG_18__SCAN_IN;
  assign n14851 = ~P1_STATE_REG_SCAN_IN & ~n14827;
  assign n14832 = ~n17072 ^ P1_REG1_REG_19__SCAN_IN;
  assign n14829 = ~n14828 | ~P1_REG1_REG_18__SCAN_IN;
  assign n14838 = ~n14837 | ~n14836;
  assign n14843 = ~P1_ADDR_REG_19__SCAN_IN | ~n14842;
  assign P1_U3260 = ~n14844 | ~n14843;
  assign n14861 = ~n14850 & ~n15689;
  assign n14857 = ~n16544 & ~n17136;
  assign n14855 = ~n14851;
  assign n14854 = ~n14853 | ~n14852;
  assign n14856 = ~n14855 | ~n14854;
  assign n14858 = ~n14857 & ~n14856;
  assign P1_U3217 = ~n14863 | ~n14862;
  assign n14865 = ~P2_ADDR_REG_19__SCAN_IN | ~n14864;
  assign n14886 = ~n14866 | ~n14865;
  assign n14872 = n16472 ^ P2_REG1_REG_19__SCAN_IN;
  assign n14869 = ~P2_REG1_REG_18__SCAN_IN & ~n14876;
  assign n14880 = n16472 ^ P2_REG2_REG_19__SCAN_IN;
  assign n14877 = ~P2_REG2_REG_18__SCAN_IN & ~n14876;
  assign n14888 = ~n14887 | ~n16472;
  assign P2_U3264 = ~n14889 | ~n14888;
  assign n14903 = n15530 & n14895;
  assign n14897 = ~n15869 | ~n16334;
  assign n14896 = ~P2_REG3_REG_21__SCAN_IN | ~P2_U3152;
  assign n14899 = ~n14897 | ~n14896;
  assign n16311 = ~n16299;
  assign n14898 = ~n15872 & ~n16311;
  assign n14901 = ~n14899 & ~n14898;
  assign P2_U3225 = ~n14905 | ~n14904;
  assign n17014 = ~n16754 | ~n16866;
  assign n14967 = ~n14908 & ~n16867;
  assign n14911 = ~n15582 & ~n15595;
  assign n14910 = ~n14924 & ~n15594;
  assign n14912 = ~n14911 & ~n14910;
  assign n14914 = ~n15745 & ~P1_REG2_REG_22__SCAN_IN;
  assign n14918 = ~n15231 & ~n15763;
  assign n14917 = n15230 & n15407;
  assign n14919 = ~n14918 & ~n14917;
  assign n14926 = ~n14923 & ~n17012;
  assign P1_U3269 = ~n14929 | ~n14928;
  assign n14932 = ~n14930 | ~n15791;
  assign n14939 = ~n15806 | ~P1_REG1_REG_22__SCAN_IN;
  assign P1_U3545 = ~n14940 | ~n14939;
  assign n14942 = ~n15801 | ~P1_REG0_REG_22__SCAN_IN;
  assign P1_U3513 = ~n14943 | ~n14942;
  assign n14956 = ~n15086 & ~n14947;
  assign n14954 = ~n16739 | ~n17132;
  assign n14950 = ~n16534 | ~n15696;
  assign n14949 = ~P1_REG3_REG_20__SCAN_IN | ~P1_U3084;
  assign n14951 = ~n14950 | ~n14949;
  assign P1_U3231 = ~n14958 | ~n14957;
  assign n14959 = ~P2_IR_REG_31__SCAN_IN | ~P2_STATE_REG_SCAN_IN;
  assign n14960 = n14959 | P2_IR_REG_30__SCAN_IN;
  assign n14964 = ~n14961 & ~n14960;
  assign n15370 = ~P1_DATAO_REG_31__SCAN_IN;
  assign n14963 = ~n14962 & ~n15370;
  assign n14965 = ~n14964 & ~n14963;
  assign P2_U3327 = ~n14966 | ~n14965;
  assign n17016 = ~n16865 & ~n16762;
  assign n15153 = ~n14968 | ~n16754;
  assign n14971 = ~n15697 | ~n15636;
  assign n14970 = ~n15512 | ~n17091;
  assign n14972 = ~n14971 | ~n14970;
  assign n15158 = ~n14979 | ~n14978;
  assign n14988 = ~n15063 | ~n15762;
  assign n14985 = n15510 & n15407;
  assign P1_U3268 = ~n14992 | ~n14991;
  assign n14999 = ~n14996 & ~n14995;
  assign n15006 = n15003 | n15002;
  assign n15004 = ~n16516 | ~P2_REG1_REG_21__SCAN_IN;
  assign P2_U3541 = ~n15005 | ~n15004;
  assign n15007 = ~n16511 | ~P2_REG0_REG_21__SCAN_IN;
  assign P2_U3509 = ~n15008 | ~n15007;
  assign n15021 = n15530 & n15040;
  assign n15015 = ~n15532 | ~n16322;
  assign n15014 = ~P2_REG3_REG_22__SCAN_IN | ~P2_U3152;
  assign n15017 = ~n15015 | ~n15014;
  assign n15016 = ~n15535 & ~n15030;
  assign n15019 = ~n15017 & ~n15016;
  assign P2_U3237 = ~n15023 | ~n15022;
  assign n15026 = ~n15025 & ~n16012;
  assign n15050 = ~n15027 & ~n15026;
  assign n15033 = ~n15030 & ~n15713;
  assign n15032 = ~n15031 & ~n16488;
  assign n15034 = ~n15033 & ~n15032;
  assign n15038 = n15720 | P2_REG2_REG_22__SCAN_IN;
  assign n15042 = ~n15848 & ~n16337;
  assign n15041 = n15725 & n15040;
  assign n15045 = ~n15042 & ~n15041;
  assign P2_U3274 = ~n15049 | ~n15048;
  assign n15058 = ~n16516 | ~P2_REG1_REG_22__SCAN_IN;
  assign P2_U3542 = ~n15059 | ~n15058;
  assign n15061 = ~n16511 | ~P2_REG0_REG_22__SCAN_IN;
  assign P2_U3510 = ~n15062 | ~n15061;
  assign n15064 = ~n15160 | ~n15793;
  assign n15073 = n15070 | n15069;
  assign n15071 = ~n15806 | ~P1_REG1_REG_23__SCAN_IN;
  assign P1_U3546 = ~n15072 | ~n15071;
  assign n15074 = ~n15801 | ~P1_REG0_REG_23__SCAN_IN;
  assign P1_U3514 = ~n15075 | ~n15074;
  assign n15079 = ~n15077 & ~n15076;
  assign n15096 = ~n15086 & ~n15085;
  assign n15090 = ~n15088 | ~n15696;
  assign n15089 = ~P1_REG3_REG_21__SCAN_IN | ~P1_U3084;
  assign n15091 = ~n15090 | ~n15089;
  assign n15093 = ~n15512 | ~n17132;
  assign P1_U3221 = ~n15098 | ~n15097;
  assign n15102 = ~n15101 & ~n15100;
  assign n15124 = ~n15103 & ~n15102;
  assign n15107 = ~n16367 & ~n15713;
  assign n15106 = ~n16338 & ~n16488;
  assign n15108 = ~n15107 & ~n15106;
  assign n15112 = n15720 | P2_REG2_REG_23__SCAN_IN;
  assign n15117 = ~n15115 & ~n15848;
  assign n15116 = n15725 & n15142;
  assign P2_U3273 = ~n15123 | ~n15122;
  assign n15126 = ~n16348 | ~n16502;
  assign n15132 = ~n16516 | ~P2_REG1_REG_23__SCAN_IN;
  assign P2_U3543 = ~n15133 | ~n15132;
  assign n15135 = ~n16511 | ~P2_REG0_REG_23__SCAN_IN;
  assign P2_U3511 = ~n15136 | ~n15135;
  assign n15150 = n15530 & n15142;
  assign n15144 = ~n15532 | ~n16334;
  assign n15143 = ~P2_REG3_REG_23__SCAN_IN | ~P2_U3152;
  assign n15146 = ~n15144 | ~n15143;
  assign n15145 = ~n15535 & ~n16367;
  assign n15148 = ~n15146 & ~n15145;
  assign n15147 = ~n15867 | ~n16348;
  assign P2_U3218 = ~n15152 | ~n15151;
  assign n15297 = ~n15154 | ~n16768;
  assign n15156 = ~n15159 | ~n17091;
  assign n15162 = ~n15158 & ~n17016;
  assign n15305 = ~n15162 & ~n15161;
  assign n15164 = ~n16781 | ~n15636;
  assign n15192 = ~n15167 & ~n15166;
  assign n15168 = n15745 | P1_REG2_REG_24__SCAN_IN;
  assign n15176 = ~n15175 & ~n15763;
  assign n15178 = ~n15585 | ~n15407;
  assign P1_U3267 = ~n15183 | ~n15182;
  assign n15188 = n15186 | n15185;
  assign n15187 = ~n15579 | ~n15793;
  assign n15193 = ~n15801 | ~P1_REG0_REG_24__SCAN_IN;
  assign P1_U3515 = ~n15194 | ~n15193;
  assign n15196 = ~n15806 | ~P1_REG1_REG_24__SCAN_IN;
  assign P1_U3547 = ~n15197 | ~n15196;
  assign n15199 = ~n15254 | ~n15212;
  assign n15200 = ~n15214 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n16520 = ~n15201 | ~n15200;
  assign n15204 = ~n15202 | ~n15212;
  assign n15760 = ~n16520 & ~n15205;
  assign n15207 = ~n15218 | ~P1_REG2_REG_30__SCAN_IN;
  assign n15206 = ~n17087 | ~P1_B_REG_SCAN_IN;
  assign n15740 = ~n15636 | ~n15206;
  assign n15219 = ~n15745 | ~n15360;
  assign n15208 = ~n15207 | ~n15219;
  assign P1_U3262 = ~n15211 | ~n15210;
  assign n15216 = ~n15213 | ~n15212;
  assign n15215 = ~n15214 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n16836 = ~n15216 | ~n15215;
  assign n15220 = ~n15218 | ~P1_REG2_REG_31__SCAN_IN;
  assign n15221 = ~n15220 | ~n15219;
  assign P1_U3261 = ~n15224 | ~n15223;
  assign n15228 = ~n15226 & ~n15225;
  assign n15237 = ~n17130 | ~n15230;
  assign n15233 = ~n16739 | ~n15696;
  assign n15232 = ~P1_REG3_REG_22__SCAN_IN | ~P1_U3084;
  assign n15234 = ~n15233 | ~n15232;
  assign n15238 = ~n15582 & ~n15689;
  assign P1_U3233 = ~n15241 | ~n15240;
  assign n15243 = ~n16362 | ~n16502;
  assign n15249 = ~n16516 | ~P2_REG1_REG_24__SCAN_IN;
  assign P2_U3544 = ~n15250 | ~n15249;
  assign n15252 = ~n16511 | ~P2_REG0_REG_24__SCAN_IN;
  assign P2_U3512 = ~n15253 | ~n15252;
  assign n15255 = ~n15258 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n15260 = ~n15257 | ~n10310;
  assign n15259 = ~n15258 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n16411 = ~n16503;
  assign n15962 = ~n15967;
  assign n15262 = ~n15261 | ~P2_B_REG_SCAN_IN;
  assign n15835 = ~n15549 | ~n15262;
  assign n15377 = ~n15720 | ~n15452;
  assign n15263 = ~n15488 | ~P2_REG2_REG_30__SCAN_IN;
  assign n15264 = ~n15377 | ~n15263;
  assign P2_U3266 = ~n15267 | ~n15266;
  assign n15462 = ~n15269 | ~n15268;
  assign n16018 = ~n15271 & ~n15270;
  assign n15273 = n10644 | n15272;
  assign n15277 = ~n15275 | ~n15274;
  assign n15479 = ~n15277 | ~n15276;
  assign n15280 = ~n16367 & ~n16488;
  assign n15279 = ~n16393 & ~n15713;
  assign n15284 = n15337 | n16472;
  assign n15286 = ~n15725 | ~n15529;
  assign n15290 = n15289 | n15288;
  assign n15294 = ~n15488 | ~P2_REG2_REG_25__SCAN_IN;
  assign P2_U3271 = ~n15295 | ~n15294;
  assign n15391 = ~n15298 | ~n16771;
  assign n16857 = ~n16781 & ~n16778;
  assign n15302 = ~n16816 & ~n15595;
  assign n15301 = ~n15509 & ~n15594;
  assign n15303 = ~n15302 & ~n15301;
  assign n15307 = ~n15305 | ~n17018;
  assign n15401 = ~n15307 | ~n15306;
  assign n15329 = ~n15309 & ~n15308;
  assign n15310 = n15745 | P1_REG2_REG_25__SCAN_IN;
  assign n15317 = n15691 & n15407;
  assign n15315 = ~n15323 | ~n15762;
  assign n15318 = n15317 | n15316;
  assign P1_U3266 = ~n15321 | ~n15320;
  assign n15324 = ~n16782 | ~n15793;
  assign n15332 = ~n15329 | ~n15328;
  assign n15330 = ~n15801 | ~P1_REG0_REG_25__SCAN_IN;
  assign P1_U3516 = ~n15331 | ~n15330;
  assign n15333 = ~n15806 | ~P1_REG1_REG_25__SCAN_IN;
  assign P1_U3548 = ~n15334 | ~n15333;
  assign n15340 = n15338 | n15337;
  assign n15339 = ~n15531 | ~n16502;
  assign n15347 = ~n15344 | ~n15343;
  assign n15345 = ~n16511 | ~P2_REG0_REG_25__SCAN_IN;
  assign P2_U3513 = ~n15346 | ~n15345;
  assign n15348 = ~n16516 | ~P2_REG1_REG_25__SCAN_IN;
  assign P2_U3545 = ~n15349 | ~n15348;
  assign n15356 = ~n15353 | ~n15352;
  assign n15354 = ~n15806 | ~P1_REG1_REG_30__SCAN_IN;
  assign P1_U3553 = ~n15355 | ~n15354;
  assign n15357 = ~n15801 | ~P1_REG0_REG_30__SCAN_IN;
  assign P1_U3521 = ~n15358 | ~n15357;
  assign n15366 = ~n15363 | ~n15362;
  assign n15364 = ~n15806 | ~P1_REG1_REG_31__SCAN_IN;
  assign P1_U3554 = ~n15365 | ~n15364;
  assign n15367 = ~n15801 | ~P1_REG0_REG_31__SCAN_IN;
  assign P1_U3522 = ~n15368 | ~n15367;
  assign n15373 = ~n15369 & ~n9036;
  assign n15376 = ~n15488 | ~P2_REG2_REG_31__SCAN_IN;
  assign n15378 = ~n15377 | ~n15376;
  assign P2_U3265 = ~n15381 | ~n15380;
  assign n15388 = ~n15385 | ~n15384;
  assign n15386 = ~n16516 | ~P2_REG1_REG_30__SCAN_IN;
  assign P2_U3550 = ~n15387 | ~n15386;
  assign n15389 = ~n16511 | ~P2_REG0_REG_30__SCAN_IN;
  assign P2_U3518 = ~n15390 | ~n15389;
  assign n15392 = ~n15391 & ~n17024;
  assign n16864 = ~n16787 | ~n16814;
  assign n17026 = ~n15393 & ~n16856;
  assign n15592 = ~n15395 | ~n17026;
  assign n15398 = ~n16777 & ~n15594;
  assign n15397 = ~n17135 & ~n15595;
  assign n15399 = ~n15398 & ~n15397;
  assign n15403 = ~n15401 | ~n17024;
  assign n15601 = ~n15403 | ~n15402;
  assign n15428 = ~n15406 & ~n15405;
  assign n15413 = n15812 & n15407;
  assign n15415 = n15745 | P1_REG2_REG_26__SCAN_IN;
  assign P1_U3265 = ~n15420 | ~n15419;
  assign n15425 = n15424 | n15423;
  assign n15431 = ~n15428 | ~n15427;
  assign n15429 = ~n15806 | ~P1_REG1_REG_26__SCAN_IN;
  assign P1_U3549 = ~n15430 | ~n15429;
  assign n15432 = ~n15801 | ~P1_REG0_REG_26__SCAN_IN;
  assign P1_U3517 = ~n15433 | ~n15432;
  assign n15437 = ~n15435 | ~n15434;
  assign n15447 = n15530 & n15439;
  assign n15441 = ~n15532 | ~n16347;
  assign n15440 = ~P2_REG3_REG_24__SCAN_IN | ~P2_U3152;
  assign n15443 = ~n15441 | ~n15440;
  assign n15442 = ~n15535 & ~n16379;
  assign n15444 = ~n15443 & ~n15442;
  assign P2_U3231 = ~n15449 | ~n15448;
  assign n15458 = ~n15455 | ~n15454;
  assign n15456 = ~n16511 | ~P2_REG0_REG_31__SCAN_IN;
  assign P2_U3519 = ~n15457 | ~n15456;
  assign n15459 = ~n16516 | ~P2_REG1_REG_31__SCAN_IN;
  assign P2_U3551 = ~n15460 | ~n15459;
  assign n15560 = ~n15465 & ~n15464;
  assign n15942 = ~n15558 & ~n16393;
  assign n15470 = ~n15492 | ~n15847;
  assign n15469 = ~n15558 | ~n15566;
  assign n15477 = n15472 | n15471;
  assign n15475 = ~n15725 | ~n15473;
  assign n15474 = ~n15488 | ~P2_REG2_REG_26__SCAN_IN;
  assign n15476 = ~n15475 | ~n15474;
  assign n15480 = ~n15479 | ~n16018;
  assign n15545 = ~n15480 | ~n15938;
  assign n15498 = ~n15487 & ~n15486;
  assign n15489 = n15498 | n15488;
  assign P2_U3270 = ~n15490 | ~n15489;
  assign n15501 = ~n15498 | ~n15497;
  assign n15499 = ~n16511 | ~P2_REG0_REG_26__SCAN_IN;
  assign P2_U3514 = ~n15500 | ~n15499;
  assign n15502 = ~n16516 | ~P2_REG1_REG_26__SCAN_IN;
  assign P2_U3546 = ~n15503 | ~n15502;
  assign n15507 = ~n15505 & ~n15504;
  assign n15520 = ~n15509 & ~n15689;
  assign n15518 = ~n17130 | ~n15510;
  assign n15514 = ~n15512 | ~n15696;
  assign n15513 = ~P1_REG3_REG_23__SCAN_IN | ~P1_U3084;
  assign n15515 = ~n15514 | ~n15513;
  assign P1_U3214 = ~n15522 | ~n15521;
  assign n15541 = n15530 & n15529;
  assign n15534 = ~n15532 | ~n16363;
  assign n15533 = ~P2_REG3_REG_25__SCAN_IN | ~P2_U3152;
  assign n15537 = ~n15534 | ~n15533;
  assign n15536 = ~n15535 & ~n16393;
  assign n15538 = ~n15537 & ~n15536;
  assign P2_U3227 = ~n15543 | ~n15542;
  assign n16030 = ~n15544 & ~n15828;
  assign n15546 = ~n15545 & ~n15940;
  assign n15551 = ~n15557 | ~n15550;
  assign n15664 = ~n15554 & ~n15553;
  assign n15555 = n15720 | P2_REG2_REG_27__SCAN_IN;
  assign n15706 = ~n15562 & ~n15561;
  assign n15866 = ~n15564;
  assign n15570 = ~n15866 & ~n15850;
  assign n15567 = ~n16436 | ~n15566;
  assign n15571 = n15570 | n15569;
  assign P2_U3269 = ~n15574 | ~n15573;
  assign n15589 = ~n16777 & ~n15689;
  assign n15580 = ~P1_REG3_REG_24__SCAN_IN | ~P1_U3084;
  assign n15583 = ~n15582 & ~n17136;
  assign n15586 = ~n17130 | ~n15585;
  assign P1_U3227 = ~n15591 | ~n15590;
  assign n15633 = ~n15592 | ~n16864;
  assign n15597 = ~n16816 & ~n15594;
  assign n15596 = ~n15752 & ~n15595;
  assign n15603 = ~n15601 | ~n15600;
  assign n15644 = ~n15603 | ~n15602;
  assign n15627 = ~n15605 & ~n15604;
  assign n15606 = n15745 | P1_REG2_REG_27__SCAN_IN;
  assign n15614 = ~n15621 | ~n15762;
  assign n15612 = ~n16854 & ~n15763;
  assign n15611 = ~n15766 & ~n15610;
  assign P1_U3264 = ~n15618 | ~n15617;
  assign n15630 = ~n15627 | ~n15626;
  assign n15628 = ~n15801 | ~P1_REG0_REG_27__SCAN_IN;
  assign P1_U3518 = ~n15629 | ~n15628;
  assign n15631 = ~n15806 | ~P1_REG1_REG_27__SCAN_IN;
  assign P1_U3550 = ~n15632 | ~n15631;
  assign n16947 = ~n16854 | ~n16853;
  assign n15734 = ~n15634 | ~n16947;
  assign n15638 = ~n17131 | ~n15636;
  assign n15637 = ~n16853 | ~n17091;
  assign n15678 = ~n15640 & ~n15639;
  assign n15641 = n15745 | P1_REG2_REG_28__SCAN_IN;
  assign n15649 = ~n15766 & ~n17128;
  assign P1_U3263 = ~n15656 | ~n15655;
  assign n15668 = ~n15665 | ~n15664;
  assign n15666 = ~n16511 | ~P2_REG0_REG_27__SCAN_IN;
  assign P2_U3515 = ~n15667 | ~n15666;
  assign n15669 = ~n16516 | ~P2_REG1_REG_27__SCAN_IN;
  assign P2_U3547 = ~n15670 | ~n15669;
  assign n15681 = ~n15678 | ~n15677;
  assign n15679 = ~n15801 | ~P1_REG0_REG_28__SCAN_IN;
  assign P1_U3519 = ~n15680 | ~n15679;
  assign n15682 = ~n15806 | ~P1_REG1_REG_28__SCAN_IN;
  assign P1_U3551 = ~n15683 | ~n15682;
  assign n15701 = ~n16816 & ~n15689;
  assign n15693 = P1_STATE_REG_SCAN_IN | n15690;
  assign n15692 = ~n15691 | ~n17130;
  assign n15694 = ~n15693 | ~n15692;
  assign n15698 = ~n15697 | ~n15696;
  assign P1_U3223 = ~n15703 | ~n15702;
  assign n15823 = ~n15708 & ~n15707;
  assign n16406 = ~n15777 | ~n15834;
  assign n16414 = ~n15777 & ~n15834;
  assign n16022 = ~n16413 & ~n16414;
  assign n15715 = ~n16405 & ~n16488;
  assign n15714 = ~n16410 & ~n15713;
  assign n15783 = ~n15719 & ~n15718;
  assign n15721 = n15720 | P2_REG2_REG_28__SCAN_IN;
  assign n15726 = n15725 & n15724;
  assign P2_U3268 = ~n15733 | ~n15732;
  assign n16861 = ~n17110 | ~n15752;
  assign n15735 = ~n15734 | ~n16861;
  assign n15737 = ~n15735 | ~n16794;
  assign n17064 = ~n16520 | ~n15736;
  assign n16951 = ~n16520 & ~n15736;
  assign n17023 = ~n16801 & ~n16951;
  assign n15744 = ~n15739 & ~n15738;
  assign n15742 = n17062 | n15740;
  assign n15741 = ~n17112 | ~n17091;
  assign n15798 = ~n15744 & ~n15743;
  assign n15746 = n15745 | P1_REG2_REG_29__SCAN_IN;
  assign n15750 = ~n15751 & ~n15752;
  assign n15753 = ~n15748 | ~n17110;
  assign n15749 = ~n15753 | ~n17023;
  assign n15757 = n15750 | n15749;
  assign n15755 = ~n15751 & ~n17023;
  assign n15754 = ~n15753 | ~n15752;
  assign n15756 = ~n15755 | ~n15754;
  assign n15772 = ~n15790 & ~n15758;
  assign n15767 = ~n15766 & ~n15765;
  assign P1_U3355 = ~n15774 | ~n15773;
  assign n15786 = ~n15783 | ~n15782;
  assign n15784 = ~n16511 | ~P2_REG0_REG_28__SCAN_IN;
  assign P2_U3516 = ~n15785 | ~n15784;
  assign n15787 = ~n16516 | ~P2_REG1_REG_28__SCAN_IN;
  assign P2_U3548 = ~n15788 | ~n15787;
  assign n15797 = ~n15790 & ~n15789;
  assign n15799 = ~n15797 & ~n15796;
  assign n15803 = ~n15805 | ~n15800;
  assign n15802 = ~n15801 | ~P1_REG0_REG_29__SCAN_IN;
  assign n15808 = ~n15805 | ~n15804;
  assign n15807 = ~n15806 | ~P1_REG1_REG_29__SCAN_IN;
  assign n15818 = ~n15812 | ~n17130;
  assign n15814 = ~n17132 | ~n16853;
  assign n15813 = ~P1_REG3_REG_26__SCAN_IN | ~P1_U3084;
  assign n15815 = ~n15814 | ~n15813;
  assign n15819 = ~n16777 & ~n17136;
  assign P1_U3238 = ~n15822 | ~n15821;
  assign n15827 = ~n15826 & ~n15825;
  assign n16499 = n15827 ^ n16024;
  assign n15842 = ~n16499 & ~n14769;
  assign n15947 = ~n15828 & ~n16413;
  assign n15831 = ~n15830 | ~n16425;
  assign n15838 = ~n15834 & ~n16488;
  assign n15836 = ~n16452;
  assign n15837 = ~n15836 & ~n15835;
  assign n15841 = ~n15840 | ~n15839;
  assign n16509 = ~n15842 & ~n15841;
  assign n15844 = ~n16509 | ~n15720;
  assign n15843 = n15720 | P2_REG2_REG_29__SCAN_IN;
  assign n15856 = ~n16499 & ~n15845;
  assign n15851 = ~n15850 & ~n15849;
  assign P2_U3267 = ~n15858 | ~n15857;
  assign n15862 = ~n15860 & ~n15859;
  assign n15864 = ~n15862 & ~n15861;
  assign n15880 = ~n15863 | ~n15864;
  assign n15878 = ~n15866 & ~n15865;
  assign n15871 = ~n15869 | ~n15868;
  assign n15870 = ~P2_REG3_REG_27__SCAN_IN | ~P2_U3152;
  assign n15874 = ~n15871 | ~n15870;
  assign n15873 = ~n15872 & ~n16393;
  assign n15875 = ~n15874 & ~n15873;
  assign P2_U3216 = ~n15880 | ~n15879;
  assign n16462 = ~n15961 | ~n15967;
  assign n16305 = ~n16294 & ~n15881;
  assign n15885 = ~n15883 | ~n15882;
  assign n15886 = ~n15885 | ~n15884;
  assign n15911 = ~n16293 & ~n15886;
  assign n15896 = ~n15895 & ~n15894;
  assign n15898 = ~n16203 & ~n16189;
  assign n15900 = ~n15899 & ~n15898;
  assign n15903 = ~n16252 & ~n15902;
  assign n15908 = ~n16063 & ~n15907;
  assign n16308 = ~n15914 | ~n15913;
  assign n15921 = ~n15919 & ~n15918;
  assign n15923 = ~n15921 | ~n15920;
  assign n15927 = ~n15925 & ~n15924;
  assign n15933 = ~n15931 | ~n15930;
  assign n15937 = ~n15935 & ~n15934;
  assign n15939 = ~n15937 | ~n15936;
  assign n15944 = ~n15943 & ~n15942;
  assign n15950 = ~n15947 | ~n15946;
  assign n15956 = ~n15950 | ~n15949;
  assign n15951 = ~n15956 | ~n15953;
  assign n15952 = ~n15951 | ~n16449;
  assign n15957 = ~n15967 | ~n16452;
  assign n15963 = ~n15960 | ~n15959;
  assign n16463 = ~n15968 | ~n15962;
  assign n16041 = ~n15963 | ~n16463;
  assign n15964 = ~n16452 | ~n16031;
  assign n16482 = ~n16041 & ~n15966;
  assign n16033 = n16482 | n16031;
  assign n15974 = ~n15970 & ~n15969;
  assign n15973 = ~n15972 & ~n15971;
  assign n15980 = ~n15974 | ~n15973;
  assign n15978 = ~n15976 & ~n15975;
  assign n15979 = ~n15978 | ~n15977;
  assign n15982 = ~n15980 & ~n15979;
  assign n15983 = ~n15982 | ~n15981;
  assign n15985 = ~n15984 & ~n15983;
  assign n15987 = ~n15986 | ~n15985;
  assign n15990 = ~n15988 & ~n15987;
  assign n15991 = ~n15990 | ~n15989;
  assign n15993 = ~n15992 & ~n15991;
  assign n15995 = ~n15994 | ~n15993;
  assign n15999 = ~n15996 & ~n15995;
  assign n15998 = ~n15997;
  assign n16000 = ~n15999 | ~n15998;
  assign n16002 = ~n16001 & ~n16000;
  assign n16004 = ~n16003 | ~n16002;
  assign n16005 = ~n16067 & ~n16004;
  assign n16007 = ~n16006 | ~n16005;
  assign n16009 = ~n16008 & ~n16007;
  assign n16011 = ~n16010 | ~n16009;
  assign n16013 = ~n16012 & ~n16011;
  assign n16015 = ~n16014 | ~n16013;
  assign n16017 = ~n16016 & ~n16015;
  assign n16035 = ~n16032 | ~n16031;
  assign n16034 = ~n16033 | ~n16035;
  assign n16047 = ~n16037 | ~n16036;
  assign n16040 = ~n16039 & ~n16038;
  assign n16042 = ~n9039;
  assign n16050 = ~n16405 | ~n16461;
  assign n16049 = ~n16048 | ~n16391;
  assign n16052 = ~n16051 | ~n16461;
  assign n16058 = ~n16053 | ~n16052;
  assign n16055 = ~n16054 | ~n16391;
  assign n16057 = ~n16056 | ~n16055;
  assign n16059 = ~n16058 | ~n16057;
  assign n16060 = ~n16067 & ~n16059;
  assign n16065 = ~n16062 & ~n16391;
  assign n16064 = ~n16063 & ~n16461;
  assign n16066 = ~n16065 & ~n16064;
  assign n16069 = ~n16090 | ~n16461;
  assign n16068 = ~n16070 | ~n16391;
  assign n16100 = ~n16087;
  assign n16072 = ~n16100 & ~n16070;
  assign n16075 = ~n16073 & ~n16461;
  assign n16074 = ~n16093 & ~n16391;
  assign n16092 = ~n16075 & ~n16074;
  assign n16077 = ~n16092 | ~n16076;
  assign n16078 = ~n16077 | ~n16461;
  assign n16089 = ~n16079 & ~n16078;
  assign n16083 = ~n16082 ^ n16081;
  assign n16086 = ~n16083 & ~n10645;
  assign n16085 = ~n16084 & ~n16471;
  assign n16099 = ~n16086 & ~n16085;
  assign n16088 = ~n16091 | ~n16070;
  assign n16098 = ~n16089 | ~n16088;
  assign n16096 = ~n16091 | ~n16090;
  assign n16105 = ~n16092;
  assign n16094 = ~n16105 & ~n16093;
  assign n16095 = ~n16094 & ~n16461;
  assign n16097 = ~n16096 | ~n16095;
  assign n16103 = ~n16098 | ~n16097;
  assign n16101 = ~n16099;
  assign n16107 = ~n16103 | ~n16102;
  assign n16123 = ~n16107 | ~n16106;
  assign n16109 = ~n16124 | ~n16391;
  assign n16108 = ~n16125 | ~n16461;
  assign n16122 = ~n16109 | ~n16108;
  assign n16121 = ~n16123 & ~n16122;
  assign n16113 = ~n16110 & ~n16391;
  assign n16112 = ~n16111 & ~n16461;
  assign n16114 = ~n16113 & ~n16112;
  assign n16139 = ~n16116 | ~n16115;
  assign n16118 = ~n16139 | ~n16391;
  assign n16117 = ~n16143 | ~n16461;
  assign n16119 = ~n16118 | ~n16117;
  assign n16120 = ~n16145 | ~n16119;
  assign n16131 = ~n16121 & ~n16120;
  assign n16129 = ~n16123 | ~n16122;
  assign n16127 = ~n16124 | ~n16461;
  assign n16126 = ~n16125 | ~n16391;
  assign n16128 = ~n16127 | ~n16126;
  assign n16130 = ~n16129 | ~n16128;
  assign n16159 = ~n16131 | ~n16130;
  assign n16133 = ~n16132;
  assign n16134 = ~n16133 & ~n16391;
  assign n16138 = ~n16135 | ~n16134;
  assign n16137 = ~n16151 & ~n16136;
  assign n16142 = ~n16138 & ~n16137;
  assign n16140 = ~n16139;
  assign n16141 = ~n16145 | ~n16140;
  assign n16157 = ~n16142 | ~n16141;
  assign n16144 = ~n16143;
  assign n16155 = ~n16145 | ~n16144;
  assign n16149 = ~n16147 & ~n16461;
  assign n16153 = ~n16149 | ~n16148;
  assign n16152 = ~n16151 & ~n16150;
  assign n16154 = ~n16153 & ~n16152;
  assign n16156 = ~n16155 | ~n16154;
  assign n16158 = ~n16157 | ~n16156;
  assign n16172 = ~n16159 | ~n16158;
  assign n16163 = ~n16160 & ~n16461;
  assign n16162 = ~n16161 & ~n16391;
  assign n16182 = ~n16163 & ~n16162;
  assign n16170 = ~n16182 & ~n16164;
  assign n16168 = ~n16165 | ~n16461;
  assign n16167 = ~n16166 | ~n16391;
  assign n16169 = ~n16168 | ~n16167;
  assign n16171 = ~n16170 & ~n16169;
  assign n16187 = ~n16172 | ~n16171;
  assign n16174 = ~n16205 & ~n16391;
  assign n16173 = ~n16195 & ~n16461;
  assign n16179 = ~n16176 & ~n16461;
  assign n16178 = ~n16177 & ~n16391;
  assign n16210 = ~n16179 & ~n16178;
  assign n16184 = ~n16210 | ~n16180;
  assign n16183 = ~n16182 | ~n16181;
  assign n16185 = ~n16184 | ~n16183;
  assign n16186 = ~n16198 & ~n16185;
  assign n16218 = ~n16187 | ~n16186;
  assign n16191 = ~n16188 & ~n16391;
  assign n16190 = ~n16189 & ~n16461;
  assign n16193 = ~n16219 | ~n16192;
  assign n16197 = ~n16193 | ~n16461;
  assign n16196 = ~n16206 & ~n16195;
  assign n16202 = ~n16197 & ~n16196;
  assign n16200 = ~n16210 & ~n16199;
  assign n16201 = ~n16212 | ~n16200;
  assign n16216 = ~n16202 | ~n16201;
  assign n16204 = ~n16219 | ~n16203;
  assign n16208 = ~n16204 | ~n16391;
  assign n16207 = ~n16206 & ~n16205;
  assign n16214 = ~n16208 & ~n16207;
  assign n16211 = ~n16210 & ~n16209;
  assign n16213 = ~n16212 | ~n16211;
  assign n16215 = ~n16214 | ~n16213;
  assign n16224 = ~n16218 | ~n16217;
  assign n16222 = ~n16219;
  assign n16221 = ~n16220;
  assign n16223 = ~n16222 | ~n16221;
  assign n16234 = ~n16224 | ~n16223;
  assign n16228 = ~n16225 | ~n16391;
  assign n16227 = ~n16226 | ~n16461;
  assign n16232 = ~n16229 & ~n16391;
  assign n16231 = ~n16230 & ~n16461;
  assign n16237 = ~n16232 & ~n16231;
  assign n16233 = ~n16238 | ~n16237;
  assign n16242 = ~n16234 | ~n16233;
  assign n16236 = ~n16251 & ~n16461;
  assign n16235 = ~n16252 & ~n16391;
  assign n16240 = ~n16236 & ~n16235;
  assign n16239 = ~n16238 & ~n16237;
  assign n16241 = ~n16240 & ~n16239;
  assign n16258 = ~n16242 | ~n16241;
  assign n16246 = ~n16243 | ~n16461;
  assign n16245 = ~n16244 | ~n16391;
  assign n16250 = ~n16247 & ~n16461;
  assign n16249 = ~n16248 & ~n16391;
  assign n16256 = ~n16260 & ~n16259;
  assign n16254 = ~n16251 & ~n16391;
  assign n16253 = ~n16252 & ~n16461;
  assign n16255 = ~n16254 & ~n16253;
  assign n16262 = ~n16258 | ~n16257;
  assign n16261 = ~n16260 | ~n16259;
  assign n16269 = ~n16262 | ~n16261;
  assign n16264 = ~n16266 & ~n16391;
  assign n16263 = ~n16265 & ~n16461;
  assign n16271 = ~n16264 & ~n16263;
  assign n16267 = ~n16266 | ~n16265;
  assign n16268 = ~n16271 | ~n16267;
  assign n16276 = ~n16269 | ~n16268;
  assign n16274 = ~n16271 & ~n16270;
  assign n16283 = ~n16276 | ~n16275;
  assign n16278 = ~n16277 | ~n16391;
  assign n16281 = ~n16279 | ~n16278;
  assign n16284 = ~n16280 | ~n16391;
  assign n16282 = ~n16281 | ~n16284;
  assign n16288 = ~n16283 | ~n16282;
  assign n16286 = ~n16284;
  assign n16287 = ~n16286 | ~n16285;
  assign n16289 = ~n16288 | ~n16287;
  assign n16291 = ~n16290 | ~n16289;
  assign n16307 = ~n16292 | ~n16291;
  assign n16297 = ~n16307 & ~n16293;
  assign n16295 = ~n16294;
  assign n16296 = ~n16295 | ~n16391;
  assign n16304 = ~n16297 & ~n16296;
  assign n16301 = ~n16298 | ~n16461;
  assign n16300 = ~n16299 | ~n16391;
  assign n16303 = ~n16317 | ~n16302;
  assign n16315 = ~n16304 | ~n16303;
  assign n16310 = ~n16307 & ~n16306;
  assign n16309 = ~n16308 | ~n16461;
  assign n16313 = ~n16310 & ~n16309;
  assign n16314 = ~n16313 | ~n16312;
  assign n16327 = ~n16315 | ~n16314;
  assign n16330 = ~n16317 & ~n16316;
  assign n16320 = ~n16327 & ~n16330;
  assign n16319 = ~n16321 & ~n16391;
  assign n16318 = ~n16322 & ~n16461;
  assign n16326 = ~n16320 & ~n16328;
  assign n16324 = ~n16321 & ~n16461;
  assign n16323 = ~n16322 & ~n16391;
  assign n16325 = ~n16324 & ~n16323;
  assign n16344 = ~n16326 & ~n16325;
  assign n16332 = ~n16327;
  assign n16331 = ~n16330 & ~n16329;
  assign n16336 = ~n16333 & ~n16391;
  assign n16335 = ~n16334 & ~n16461;
  assign n16340 = ~n16337 | ~n16391;
  assign n16339 = ~n16338 | ~n16461;
  assign n16343 = ~n16342 | ~n16341;
  assign n16357 = ~n16344 & ~n16343;
  assign n16346 = ~n16348 & ~n16461;
  assign n16345 = ~n16347 & ~n16391;
  assign n16349 = ~n16348 | ~n16347;
  assign n16352 = ~n16351;
  assign n16361 = ~n16357 & ~n16356;
  assign n16360 = ~n16359 & ~n16358;
  assign n16371 = ~n16361 & ~n16360;
  assign n16365 = ~n16362 & ~n16391;
  assign n16364 = ~n16363 & ~n16461;
  assign n16369 = ~n16366 | ~n16391;
  assign n16368 = ~n16367 | ~n16461;
  assign n16377 = ~n16371 | ~n16370;
  assign n16384 = ~n16377 | ~n16376;
  assign n16381 = ~n16378 | ~n16391;
  assign n16380 = ~n16379 | ~n16461;
  assign n16402 = ~n16384 | ~n16383;
  assign n16389 = ~n16392 | ~n16461;
  assign n16388 = ~n16393 | ~n16391;
  assign n16397 = ~n16390 | ~n16400;
  assign n16395 = ~n16392 | ~n16391;
  assign n16394 = ~n16393 | ~n16461;
  assign n16396 = ~n16395 | ~n16394;
  assign n16404 = ~n16397 | ~n16396;
  assign n16440 = ~n16404 | ~n16403;
  assign n16438 = ~n16439 | ~n16440;
  assign n16407 = ~n16438 | ~n16405;
  assign n16419 = ~n16407 | ~n16406;
  assign n16409 = ~n16411 | ~n16461;
  assign n16408 = ~n16410 | ~n16391;
  assign n16428 = ~n16409 | ~n16408;
  assign n16412 = ~n16411 & ~n16410;
  assign n16418 = ~n16428 & ~n16412;
  assign n16416 = ~n16413 & ~n16391;
  assign n16445 = ~n16418 & ~n16417;
  assign n16424 = ~n16419 | ~n16445;
  assign n16420 = ~n16428 | ~n16503;
  assign n16421 = ~n16420 | ~n16391;
  assign n16435 = ~n16424 | ~n16423;
  assign n16431 = ~n16426 & ~n16425;
  assign n16430 = ~n16429 | ~n16461;
  assign n16433 = ~n16431 & ~n16430;
  assign n16448 = ~n16435 | ~n16434;
  assign n16437 = ~n16436 & ~n16391;
  assign n16441 = ~n16440;
  assign n16456 = ~n16448 | ~n16447;
  assign n16460 = ~n16456 | ~n16455;
  assign n16475 = ~n16467 | ~n16466;
  assign n16470 = ~n16469 & ~n16468;
  assign n16473 = ~n16471 | ~n16491;
  assign n16476 = ~n16475 | ~n16474;
  assign n16480 = ~n16479 | ~n9039;
  assign n16484 = ~n16481 | ~n16480;
  assign n16483 = ~n16482 | ~n10888;
  assign n16485 = ~n16484 | ~n16483;
  assign n16497 = ~n16485 | ~n16492;
  assign n16490 = ~n16486;
  assign n16489 = ~n16488 & ~n16487;
  assign n16495 = ~n16490 | ~n16489;
  assign n16493 = ~n16492 | ~n16491;
  assign n16494 = n16493 & P2_B_REG_SCAN_IN;
  assign n16496 = ~n16495 | ~n16494;
  assign P2_U3244 = ~n16497 | ~n16496;
  assign n16507 = ~n16499 & ~n16498;
  assign n16508 = ~n16507 & ~n16506;
  assign n16515 = ~n16509 | ~n16508;
  assign n16513 = ~n16515 | ~n16510;
  assign n16512 = ~n16511 | ~P2_REG0_REG_29__SCAN_IN;
  assign P2_U3517 = ~n16513 | ~n16512;
  assign n16518 = ~n16515 | ~n16514;
  assign n16517 = ~n16516 | ~P2_REG1_REG_29__SCAN_IN;
  assign P2_U3549 = ~n16518 | ~n16517;
  assign n16519 = ~n17131 & ~n16688;
  assign n16522 = ~n16951 & ~n16519;
  assign n16521 = ~n16520 & ~n16688;
  assign n16800 = ~n16522 & ~n16521;
  assign n16526 = ~n16524 ^ n16843;
  assign n16525 = ~n16853 ^ n16688;
  assign n16821 = ~n16800 & ~n16529;
  assign n16533 = ~n16530 | ~n16843;
  assign n16688 = ~n16843;
  assign n16532 = ~n16531 | ~n16688;
  assign n16536 = ~n16535 & ~n16688;
  assign n16542 = ~n16549 | ~n16537;
  assign n16539 = ~n16728 | ~n16843;
  assign n16538 = ~n16544 | ~n16688;
  assign n16541 = ~n16543 | ~n16540;
  assign n16550 = ~n16549 & ~n16548;
  assign n16551 = ~n16550 & ~n16843;
  assign n16556 = ~n16553 & ~n16574;
  assign n16555 = ~n16554 | ~n16974;
  assign n16557 = ~n16556 | ~n16555;
  assign n16560 = ~n16557 | ~n16843;
  assign n16559 = ~n16558 | ~n16688;
  assign n16566 = ~n16560 | ~n16559;
  assign n16571 = ~n16562 & ~n16561;
  assign n16564 = ~n16563 & ~n16571;
  assign n16565 = ~n16564 & ~n16843;
  assign n16578 = ~n16566 & ~n16565;
  assign n16570 = ~n16568 & ~n16567;
  assign n16573 = ~n16570 & ~n16569;
  assign n17038 = ~n16571;
  assign n16572 = ~n17038 & ~n16688;
  assign n16576 = ~n16573 & ~n16572;
  assign n16575 = ~n16574 | ~n16688;
  assign n16577 = ~n16576 | ~n16575;
  assign n16586 = ~n16578 & ~n16577;
  assign n16580 = ~n16579 | ~n16901;
  assign n16584 = ~n16580 | ~n16843;
  assign n16582 = ~n16888 | ~n16581;
  assign n16583 = ~n16582 | ~n16688;
  assign n16585 = ~n16584 | ~n16583;
  assign n16594 = ~n16586 & ~n16585;
  assign n16588 = ~n16888 & ~n16688;
  assign n16587 = ~n16901 & ~n16843;
  assign n16592 = ~n16588 & ~n16587;
  assign n16591 = ~n16590 | ~n16589;
  assign n16593 = ~n16592 | ~n16591;
  assign n16602 = ~n16594 & ~n16593;
  assign n16893 = ~n16596 | ~n16595;
  assign n16597 = ~n16893 | ~n16890;
  assign n16600 = ~n16597 | ~n16688;
  assign n16900 = ~n16892 | ~n16598;
  assign n16599 = ~n16900 | ~n16843;
  assign n16601 = ~n16600 | ~n16599;
  assign n16608 = ~n16602 & ~n16601;
  assign n16604 = ~n16893 & ~n16688;
  assign n16603 = ~n16892 & ~n16843;
  assign n16605 = ~n16604 & ~n16603;
  assign n16607 = ~n16606 | ~n16605;
  assign n16612 = ~n16608 & ~n16607;
  assign n16610 = ~n16609 & ~n16899;
  assign n16611 = ~n16610 & ~n16843;
  assign n16615 = ~n16612 & ~n16611;
  assign n16907 = ~n16617 | ~n16613;
  assign n16614 = ~n16907 | ~n16843;
  assign n16621 = ~n16615 | ~n16614;
  assign n16619 = ~n16616 & ~n16688;
  assign n16618 = ~n16617 & ~n16843;
  assign n16620 = ~n16619 & ~n16618;
  assign n16623 = ~n16628 | ~n16843;
  assign n16622 = ~n16629 | ~n16688;
  assign n16626 = ~n16623 | ~n16622;
  assign n16625 = ~n16627 & ~n16626;
  assign n16635 = ~n16625 & ~n16624;
  assign n16633 = ~n16627 | ~n16626;
  assign n16631 = ~n16628 | ~n16688;
  assign n16630 = ~n16629 | ~n16843;
  assign n16632 = ~n16631 | ~n16630;
  assign n16634 = ~n16633 | ~n16632;
  assign n16642 = ~n16635 | ~n16634;
  assign n16636 = ~n16915;
  assign n16638 = ~n16636 | ~n16688;
  assign n16640 = ~n16638 | ~n16637;
  assign n16639 = ~n16935 & ~n16688;
  assign n16641 = ~n16640 & ~n16639;
  assign n16646 = ~n16914;
  assign n16644 = ~n16643 & ~n16646;
  assign n16647 = ~n16646 | ~n16688;
  assign n16649 = ~n16666 & ~n16688;
  assign n16652 = ~n16650 & ~n16649;
  assign n16651 = ~n16668 & ~n16688;
  assign n16665 = ~n16652 & ~n16651;
  assign n16654 = ~n16653 & ~n16843;
  assign n16655 = ~n16665 & ~n16654;
  assign n16681 = ~n16657 & ~n16688;
  assign n16658 = ~n16681 | ~n16678;
  assign n16663 = ~n16660 & ~n16688;
  assign n16662 = ~n16661 & ~n16843;
  assign n16664 = ~n16663 & ~n16662;
  assign n16670 = ~n16665 & ~n16664;
  assign n16667 = ~n16666 | ~n16843;
  assign n16669 = ~n16668 & ~n16667;
  assign n16675 = ~n16670 & ~n16669;
  assign n16674 = ~n16673 | ~n16688;
  assign n16676 = ~n16675 | ~n16674;
  assign n16679 = ~n16678 & ~n16688;
  assign n16682 = ~n16680 & ~n16679;
  assign n16683 = ~n16682 & ~n16681;
  assign n16686 = ~n16700 | ~n16843;
  assign n16685 = ~n16701 | ~n16688;
  assign n16691 = ~n16687 | ~n16843;
  assign n16690 = ~n16689 | ~n16688;
  assign n16695 = ~n16692 & ~n16843;
  assign n16694 = ~n16693 & ~n16688;
  assign n16703 = ~n16700 | ~n16688;
  assign n16702 = ~n16701 | ~n16843;
  assign n16704 = ~n16703 | ~n16702;
  assign n16710 = ~n16709 | ~n16708;
  assign n16715 = ~n16712 | ~n16688;
  assign n16714 = ~n16713 | ~n16843;
  assign n16719 = ~n16716 & ~n16688;
  assign n16718 = ~n16717 & ~n16843;
  assign n16722 = ~n16719 & ~n16718;
  assign n16725 = ~n16722;
  assign n16724 = ~n16723;
  assign n16730 = ~n16729 | ~n16728;
  assign n16733 = ~n16732;
  assign n16740 = ~n16739 | ~n16738;
  assign n16743 = ~n16879 & ~n16688;
  assign n16742 = ~n16875 & ~n16843;
  assign n16751 = ~n16869 | ~n16843;
  assign n16750 = ~n16866 & ~n16843;
  assign n16761 = ~n16749 & ~n16750;
  assign n16753 = ~n16867 & ~n16843;
  assign n16755 = ~n16877 & ~n16688;
  assign n16766 = ~n16865 | ~n16688;
  assign n16769 = ~n16874 | ~n16688;
  assign n16773 = ~n17051 & ~n16843;
  assign n16772 = ~n16771 & ~n16688;
  assign n16774 = ~n16773 & ~n16772;
  assign n16780 = ~n16777 | ~n16688;
  assign n16779 = ~n16778 | ~n16843;
  assign n16784 = ~n16781 & ~n16688;
  assign n16783 = ~n16782 & ~n16843;
  assign n16809 = ~n16784 & ~n16783;
  assign n16791 = ~n16786 & ~n16785;
  assign n16790 = ~n16787 ^ n16688;
  assign n16789 = ~n16788 ^ n16843;
  assign n16792 = ~n17135 | ~n16688;
  assign n16793 = ~n16854 & ~n16792;
  assign n16795 = ~n16950 | ~n16843;
  assign n16797 = ~n16861 & ~n16843;
  assign n16802 = ~n16951 | ~n16843;
  assign n16833 = ~n16825 & ~n16824;
  assign n16954 = ~n16837 & ~n17062;
  assign n16826 = ~n16954 | ~n16843;
  assign n16831 = n16833 | n16832;
  assign n16828 = ~n16954 | ~n16688;
  assign n16838 = ~n16837;
  assign n17036 = ~n16839 & ~n16838;
  assign n17031 = ~n16842 & ~n17036;
  assign n16850 = ~n16840 | ~n17031;
  assign n16848 = ~n16850 | ~n16846;
  assign n16852 = ~n16848 | ~n16847;
  assign n16966 = ~n16852 | ~n16851;
  assign n16855 = ~n16854 & ~n16853;
  assign n16858 = ~n16864 | ~n16857;
  assign n16871 = ~n16870 | ~n16869;
  assign n16876 = ~n16875;
  assign n16927 = ~n16877 & ~n16876;
  assign n16883 = ~n16879 | ~n16878;
  assign n17004 = ~n16881 & ~n16880;
  assign n16882 = ~n16887 & ~n17004;
  assign n16930 = ~n16883 & ~n16882;
  assign n16886 = ~n16885 | ~n16884;
  assign n17008 = ~n16887 & ~n16886;
  assign n16889 = ~n16899;
  assign n16895 = ~n16889 | ~n16888;
  assign n16891 = ~n16890;
  assign n16894 = ~n16892 | ~n16891;
  assign n16898 = ~n16894 | ~n16893;
  assign n16932 = ~n16895 & ~n16898;
  assign n16897 = ~n16896 & ~n17043;
  assign n16906 = ~n16932 | ~n16897;
  assign n16904 = ~n16899 & ~n16898;
  assign n16902 = ~n16900;
  assign n16903 = ~n16902 | ~n16901;
  assign n16905 = ~n16904 | ~n16903;
  assign n16908 = ~n16906 | ~n16905;
  assign n16909 = ~n16908 & ~n16907;
  assign n16911 = ~n16909 & ~n16934;
  assign n16913 = ~n16911 & ~n16910;
  assign n16912 = ~n16935;
  assign n16917 = ~n16913 & ~n16912;
  assign n16916 = ~n16915 | ~n16914;
  assign n16918 = ~n16917 & ~n16916;
  assign n16920 = ~n16919 | ~n16918;
  assign n16921 = ~n16931 | ~n16920;
  assign n16923 = ~n16922 | ~n16921;
  assign n16924 = ~n16940 | ~n16923;
  assign n16925 = ~n17008 | ~n16924;
  assign n16926 = ~n16930 | ~n16925;
  assign n16928 = ~n16927 | ~n16926;
  assign n17048 = ~n16929 & ~n16928;
  assign n16942 = ~n16930;
  assign n16938 = ~n16931;
  assign n16933 = ~n16932;
  assign n16936 = ~n16934 & ~n16933;
  assign n16937 = ~n16936 | ~n16935;
  assign n16939 = ~n16938 & ~n16937;
  assign n16941 = ~n16940 | ~n16939;
  assign n16943 = ~n17041 | ~n17046;
  assign n16944 = ~n17048 | ~n16943;
  assign n16948 = ~n16947 | ~n16946;
  assign n16952 = n17058 | n16949;
  assign n16968 = ~n16966 | ~n16965;
  assign n17083 = ~n16968 | ~n16967;
  assign n16970 = ~n16969;
  assign n16973 = ~n16971 | ~n16970;
  assign n16978 = ~n16973 & ~n16972;
  assign n17040 = ~n16975 | ~n16974;
  assign n16977 = ~n16976 & ~n17040;
  assign n16980 = ~n16978 | ~n16977;
  assign n16982 = ~n16980 & ~n16979;
  assign n16984 = ~n16982 | ~n16981;
  assign n16986 = n16984 | n16983;
  assign n16988 = ~n16986 & ~n16985;
  assign n16990 = ~n16988 | ~n16987;
  assign n16992 = ~n16990 & ~n16989;
  assign n16993 = ~n16992 | ~n16991;
  assign n16995 = ~n16994 & ~n16993;
  assign n16997 = ~n16996 | ~n16995;
  assign n16999 = ~n16998 & ~n16997;
  assign n17001 = ~n17000 | ~n16999;
  assign n17003 = ~n17002 & ~n17001;
  assign n17006 = ~n17004 | ~n17003;
  assign n17007 = ~n17006 & ~n17005;
  assign n17009 = ~n17008 | ~n17007;
  assign n17011 = ~n17010 & ~n17009;
  assign n17015 = ~n17014 & ~n17013;
  assign n17017 = ~n17016 | ~n17015;
  assign n17019 = ~n17018 & ~n17017;
  assign n17039 = ~n17038 | ~n17037;
  assign n17042 = ~n17040 & ~n17039;
  assign n17044 = ~n17042 & ~n17041;
  assign n17045 = ~n17044 & ~n17043;
  assign n17047 = ~n17046 | ~n17045;
  assign n17068 = n17067 | n17066;
  assign n17074 = ~n17073;
  assign n17082 = ~n17081 & ~n17080;
  assign n17085 = ~n17083 | ~n17082;
  assign n17101 = ~n17085 | ~n17084;
  assign n17088 = ~n17087 | ~n17086;
  assign n17090 = ~n17089 & ~n17088;
  assign n17095 = ~n17091 | ~n17090;
  assign n17094 = ~n17093 | ~n17092;
  assign n17098 = ~n17095 | ~n17094;
  assign n17097 = ~n17096 & ~P1_U3084;
  assign n17099 = ~n17098 | ~n17097;
  assign n17100 = ~n17099 | ~P1_B_REG_SCAN_IN;
  assign P1_U3240 = ~n17101 | ~n17100;
  assign n17105 = ~n17112 | ~n17104;
  assign n17113 = ~n17112 | ~n17111;
  assign n17129 = ~n17128;
  assign n17140 = ~n17130 | ~n17129;
  assign n17134 = ~n17132 | ~n17131;
  assign n17133 = ~P1_U3084 | ~P1_REG3_REG_28__SCAN_IN;
  assign n17138 = ~n17134 | ~n17133;
  assign n17137 = ~n17136 & ~n17135;
  assign n17139 = ~n17138 & ~n17137;
  assign n17141 = ~n17140 | ~n17139;
  assign n17152 = ~n17146 & ~n17145;
  assign n17151 = ~n17150 | ~n17149;
  assign P1_U3218 = ~n17152 | ~n17151;
endmodule


