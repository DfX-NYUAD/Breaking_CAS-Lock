// Benchmark "b14_C" written by ABC on Sat Feb  8 17:46:26 2020

module b14_C ( 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN,
    REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN,
    REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN,
    REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN,
    REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN,
    REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN,
    REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN,
    REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN,
    IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN,
    IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN,
    IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN,
    IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN,
    IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN,
    IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN,
    IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN,
    IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN,
    IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN,
    IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN,
    IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, D_REG_1__SCAN_IN,
    D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
    D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
    D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
    D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
    D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
    D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
    D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
    D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
    D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
    D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
    REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
    REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
    REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
    REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
    REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
    REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
    REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
    REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
    REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
    REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
    REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
    REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
    REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
    REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
    REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
    REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
    REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
    REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
    REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
    REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
    REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
    REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
    REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
    REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
    REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
    REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
    REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
    REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
    REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
    REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
    REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
    REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
    ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
    ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
    ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
    ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
    ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
    ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
    DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
    DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
    DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
    DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
    DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
    DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
    DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
    DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
    DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
    DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
    DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
    REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
    REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
    REG3_REG_22__SCAN_IN,
    U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
    U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
    U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
    U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
    U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
    U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
    U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
    U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
    U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
    U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
    U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
    U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
    U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
    U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
    U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
    U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
    U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
    U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
    U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
    U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
    U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
    U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
    U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
    U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
    U3211, U3210, U3149, U3148, U4043  );
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
    REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
    REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
    REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
    REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
    REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
    REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
    REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
    IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
    IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
    IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
    IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
    IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
    IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
    IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
    IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
    IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
    IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
    IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
    D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN,
    D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
    D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
    D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
    D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
    D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
    D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
    D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
    D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
    D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
    REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
    REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
    REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
    REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
    REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
    REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
    REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
    REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
    REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
    REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
    REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
    REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
    REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
    REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
    REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
    REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
    REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
    REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
    REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
    REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
    REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
    REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
    REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
    REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
    REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
    REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
    REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
    REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
    REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
    REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
    REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
    REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
    ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
    ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
    ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
    ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
    ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
    ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
    ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
    DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
    DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
    DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
    DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
    DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
    DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
    DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
    DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
    DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
    B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
    REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
    REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
    U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
    U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
    U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
    U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
    U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
    U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
    U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
    U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
    U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
    U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
    U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
    U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
    U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
    U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
    U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
    U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
    U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
    U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
    U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
    U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
    U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
    U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
    U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
    U3211, U3210, U3149, U3148, U4043;
  wire n7769, n7764, n7743, n7056, n5826, n7777, n5209, n5392, n6996, n6127,
    n7501, n4415, n4506, n4444, n4633, n4948, n4396, n6698, n5436, n7746,
    n4584, n7533, n6832, n6422, n7767, n7763, n6193, n7595, n7677, n7666,
    n7676, n7683, n7593, n7609, n7603, n7450, n7608, n7602, n7447, n7320,
    n7317, n7483, n7345, n7348, n7495, n7444, n7482, n7256, n7556, n7376,
    n7690, n7314, n6913, n7330, n7375, n6910, n7554, n7253, n7492, n7519,
    n6886, n6883, n6911, n7304, n7353, n7498, n7313, n7423, n6982, n7732,
    n7245, n6907, n7255, n7484, n6760, n6903, n6973, n6763, n6981, n6881,
    n7265, n6739, n7475, n6736, n6777, n6947, n7377, n6761, n6877, n6811,
    n6805, n6958, n6980, n6814, n7262, n6774, n7404, n6758, n6803, n6737,
    n5198, n6941, n6891, n7369, n7715, n6813, n5041, n6802, n6810, n6930,
    n7264, n6772, n6734, n6827, n6800, n7112, n6824, n6730, n5091, n6927,
    n6786, n6933, n6852, n6743, n6809, n6667, n6798, n6843, n6670, n6926,
    n7111, n6931, n7587, n6642, n6669, n6922, n6620, n7291, n7334, n5090,
    n6901, n7105, n6851, n6645, n6618, n5079, n6753, n7101, n6921, n6848,
    n6492, n6854, n6617, n6661, n6729, n6711, n6747, n6495, n6595, n6584,
    n6603, n7290, n6728, n6592, n6704, n7095, n6615, n6745, n6640, n7094,
    n6420, n6491, n6594, n6526, n6591, n6657, n6413, n6720, n6487, n7092,
    n6635, n6419, n5067, n6522, n6801, n6521, n6656, n6590, n6580, n5168,
    n6538, n6417, n7091, n6411, n6490, n6536, n6579, n6581, n4901, n6534,
    n4900, n6616, n6484, n7080, n6560, n6652, n6577, n6481, n6403, n6461,
    n6533, n6455, n7544, n7547, n6438, n6558, n6479, n7509, n7546, n6434,
    n6572, n7512, n7827, n6525, n6460, n6410, n6454, n6409, n7835, n7511,
    n6380, n6448, n6555, n5064, n7674, n7825, n7069, n6433, n7753, n6430,
    n7067, n6301, n6379, n7834, n6329, n7681, n6570, n7607, n7481, n6387,
    n7471, n7759, n6443, n7063, n6300, n6326, n7751, n6377, n7374, n7443,
    n5061, n7606, n6234, n6245, n6192, n6298, n7461, n6381, n6347, n6299,
    n7490, n7329, n6325, n6242, n6278, n7399, n7459, n7470, n6426, n7230,
    n7469, n6188, n6231, n6274, n7458, n7398, n7400, n7623, n6179, n7466,
    n6875, n7396, n6215, n7227, n6241, n6272, n7455, n5154, n5196, n6866,
    n7467, n6184, n5057, n5195, n6119, n7393, n7225, n6176, n7223, n6946,
    n7250, n7464, n6169, n6823, n6874, n6252, n6864, n7394, n6694, n6691,
    n6863, n7220, n7381, n6108, n6873, n5054, n6059, n6160, n7218, n6771,
    n6056, n7246, n6116, n6690, n5988, n6515, n6692, n7389, n7380, n6770,
    n6687, n6732, n4768, n6506, n5985, n7211, n6504, n6370, n6513, n7052,
    n6503, n6639, n6367, n7209, n7051, n6673, n6366, n6588, n6682, n6674,
    n6364, n6368, n6321, n6598, n6312, n7031, n6459, n6396, n6309, n5046,
    n7217, n6349, n7030, n7104, n6359, n6383, n7215, n6350, n5242, n5241,
    n6281, n7660, n5045, n7097, n7555, n5218, n5217, n7655, n7517, n6216,
    n7641, n7691, n7102, n7713, n4881, n5298, n6315, n5237, n7552, n7692,
    n7776, n6073, n6204, n7592, n7436, n7549, n7785, n7731, n6172, n7640,
    n7257, n7714, n5844, n7735, n5613, n6155, n5235, n6696, n5184, n5230,
    n4909, n4972, n6552, n4648, n5214, n4623, n4818, n6549, n4744, n4715,
    n6424, n4767, n6474, n4621, n7717, n7716, n4674, n5229, n7643, n5232,
    n7551, n7514, n7658, n6404, n7289, n5176, n5183, n7733, n5001, n7575,
    n5260, n5310, n6372, n7778, n4675, n4696, n5314, n5252, n4906, n4816,
    n4712, n7586, n4793, n5063, n5060, n7582, n4769, n7791, n6799, n7034,
    n5289, n7003, n5240, n6141, n6153, n5175, n4622, n4945, n7525, n7789,
    n4647, n7288, n7261, n5179, n4591, n7020, n6203, n5000, n5295, n5286,
    n7068, n4919, n4966, n5273, n4943, n7333, n5292, n4546, n6719, n5148,
    n4970, n4544, n4883, n7430, n7168, n7574, n7439, n4875, n4999, n5251,
    n4879, n5825, n4861, n5239, n5236, n7431, n4840, n5160, n4836, n5231,
    n4815, n4791, n7403, n7530, n4811, n5164, n5110, n6150, n5163, n5158,
    n5152, n4941, n6632, n7496, n4694, n4566, n5171, n6134, n5155, n4691,
    n7166, n7747, n7667, n6713, n7201, n6290, n7336, n5153, n5169, n7057,
    n5145, n5123, n6471, n4671, n4619, n6092, n7138, n6441, n7120, n7793,
    n4667, n5137, n6439, n6607, n4646, n4642, n7521, n4760, n5142, n7007,
    n4998, n4764, n5014, n5126, n4994, n7008, n4742, n7698, n7252, n7823,
    n4788, n5019, n4737, n7087, n7121, n5151, n5149, n4709, n5156, n5118,
    n7283, n5208, n4713, n5876, n7829, n6540, n7072, n5139, n5894, n6341,
    n7010, n6543, n7140, n6706, n6261, n6944, n7628, n6974, n5136, n7532,
    n6819, n5906, n6467, n7143, n7177, n7123, n5811, n7013, n4996, n5078,
    n6740, n5221, n5068, n5233, n7084, n7196, n6928, n5187, n5226, n7808,
    n6407, n5182, n5246, n7073, n5238, n4850, n7178, n5532, n7085, n7414,
    n7620, n7462, n5269, n7081, n7504, n7527, n4800, n7082, n5940, n7079,
    n6889, n5327, n6162, n7392, n6196, n5994, n6937, n5009, n7397, n7411,
    n6199, n4683, n4895, n4728, n4932, n5892, n4954, n4659, n7632, n5904,
    n7268, n4753, n4799, n4777, n4703, n6731, n6068, n6663, n4776, n6621,
    n4982, n4888, n5262, n5326, n5280, n4825, n4556, n6436, n5104, n4501,
    n6382, n5305, n4514, n4575, n5937, n4849, n4632, n4898, n4536, n5207,
    n4532, n4929, n4574, n4891, n7506, n4508, n4892, n6029, n5253, n4533,
    n4752, n5087, n4845, n6016, n5206, n4631, n4702, n4981, n4928, n4727,
    n5115, n5277, n5278, n5077, n4951, n5031, n4775, n4821, n7559, n5097,
    n4658, n4651, n4555, n5901, n5003, n5302, n4950, n5004, n4682, n5303,
    n7726, n6109, n5400, n4657, n4553, n4851, n5481, n4549, n4629, n4630,
    n5470, n7699, n7308, n5028, n5261, n5267, n5266, n7538, n5024, n5102,
    n7273, n4956, n5101, n5070, n5074, n6964, n5116, n5086, n5085, n5081,
    n5467, n4625, n4983, n4496, n5503, n7668, n5114, n5200, n5466, n5694,
    n4491, n5015, n5096, n7234, n5080, n5113, n5502, n7661, n5521, n7779,
    n4510, n7650, n4886, n5388, n5501, n7757, n5026, n5396, n5711, n5465,
    n5112, n6500, n5005, n7647, n5474, n4430, n4490, n5272, n4492, n4974,
    n7775, n4486, n5095, n6779, n4451, n6083, n5105, n5518, n4949, n4528,
    n6093, n5499, n6357, n4527, n5517, n4868, n7224, n7226, n4927, n6091,
    n4961, n6316, n4539, n4890, n6306, n5902, n4959, n7485, n4505, n5500,
    n7387, n4855, n5519, n4780, n5779, n5778, n4489, n5515, n5769, n4989,
    n6151, n4936, n6680, n4988, n4755, n5514, n6062, n4685, n5557, n4794,
    n5562, n5495, n4636, n4731, n4771, n5626, n4699, n5635, n5856, n4986,
    n4388, n4718, n5632, n7395, n4504, n5623, n4804, n4442, n4866, n6355,
    n4436, n5381, n4435, n4802, n4512, n5301, n4847, n4679, n4778, n4426,
    n4935, n4853, n4960, n6914, n4914, n6624, n4803, n4893, n5032, n4394,
    n4912, n4389, n4534, n4397, n7754, n7615, n7612, n7604, n7689, n7686,
    n7662, n7675, n7682, n5339, n7583, n7711, n7445, n7570, n7535, n7315,
    n7557, n7531, n7343, n7493, n7526, n7298, n5299, n7297, n6953, n7491,
    n6950, n7293, n5199, n6908, n7244, n7663, n7656, n6948, n7233, n5119,
    n7231, n7254, n7408, n6826, n7646, n5111, n7590, n5197, n7114, n7435,
    n5094, n6880, n6890, n6856, n7342, n6733, n6853, n6757, n6785, n6818,
    n7433, n7258, n6902, n6816, n6807, n7301, n6666, n5185, n6644, n6641,
    n6846, n7096, n6494, n6845, n6613, n6602, n6583, n6660, n6638, n6462,
    n6486, n6465, n6464, n6789, n6519, n6415, n6589, n7090, n6582, n6391,
    n6516, n6388, n7078, n6390, n7070, n6530, n6605, n6453, n6327, n6303,
    n7543, n4885, n7639, n6330, n6571, n6478, n4882, n7508, n7634, n6428,
    n6246, n6235, n7633, n7680, n6243, n6405, n7599, n7635, n6442, n6386,
    n7402, n6286, n7061, n7630, n6535, n6296, n7598, n6189, n6285, n7670,
    n7478, n6260, n7228, n5058, n6258, n7489, n7626, n4819, n6177, n7371,
    n7229, n6339, n6323, n6180, n7619, n7328, n6120, n7617, n6187, n6117,
    n7442, n6230, n7486, n6212, n7310, n6240, n7384, n6232, n6255, n7307,
    n6978, n6222, n7385, n6876, n7249, n6822, n6175, n5193, n6820, n5191,
    n7214, n6104, n6871, n7379, n7388, n6861, n6756, n6045, n6784, n5053,
    n7212, n6850, n6677, n6685, n6101, n6808, n6755, n6765, n7113, n5982,
    n6783, n6686, n6601, n6514, n6678, n5918, n5052, n6764, n6037, n6664,
    n6781, n7032, n5912, n6665, n6599, n5049, n6501, n6511, n5961, n6362,
    n5048, n6354, n6310, n6363, n5869, n6397, n5047, n6307, n7815, n7810,
    n5814, n7693, n6475, n7103, n7213, n7812, n6423, n7060, n5297, n5755,
    n7739, n7125, n6695, n7162, n6551, n6449, n4595, n5316, n7062, n7718,
    n7550, n5997, n5216, n7119, n7585, n7089, n7066, n7645, n6110, n4594,
    n7736, n6152, n7259, n5928, n4673, n7432, n7058, n6940, n7041, n7130,
    n7133, n7053, n6658, n5213, n4695, n6984, n5161, n7059, n6456, n4670,
    n7064, n4672, n6488, n5177, n6440, n7644, n6113, n7158, n5666, n5166,
    n6030, n6012, n7132, n4940, n7071, n7074, n5133, n7323, n7055, n4968,
    n7174, n7036, n4965, n7149, n7093, n4693, n5534, n4860, n6788, n5309,
    n5288, n4863, n4810, n7124, n7011, n5312, n5172, n4874, n5285, n6999,
    n6742, n4618, n4877, n6559, n4838, n4542, n4835, n5971, n7285, n4790,
    n7038, n4921, n7159, n5328, n4813, n5129, n7752, n7299, n4918, n5275,
    n4614, n5131, n5255, n7144, n5258, n4690, n4666, n5640, n7296, n4669,
    n5271, n7024, n7148, n7086, n6817, n7001, n7054, n5017, n5144, n6920,
    n6925, n4711, n4708, n7579, n7015, n4589, n4759, n5141, n4787, n4762,
    n4993, n4955, n6923, n5281, n5871, n7826, n5965, n7833, n5307, n7136,
    n6122, n6712, n4896, n4515, n7665, n5306, n4736, n6520, n6887, n4826,
    n5250, n6716, n7117, n5257, n7287, n4933, n4739, n7560, n4537, n7474,
    n5121, n7368, n5254, n5282, n5220, n5181, n4789, n4834, n4995, n4837,
    n5891, n4859, n5245, n4862, n4873, n5228, n4992, n7813, n4876, n5225,
    n4545, n4917, n4920, n4942, n7460, n7832, n6865, n4665, n4668, n5903,
    n4689, n4707, n5248, n4710, n4735, n4738, n4761, n4758, n4692, n6659,
    n6833, n4509, n4678, n4822, n4846, n4796, n6457, n5323, n4698, n5065,
    n4541, n4812, n4964, n4786, n4939, n4747, n4772, n7383, n4809, n4967,
    n4677, n4795, n5816, n5132, n4697, n5529, n4746, n5227, n5008, n4650,
    n5244, n5224, n5268, n5076, n5103, n4526, n5247, n5088, n5030, n5321,
    n4681, n4751, n4726, n4725, n4773, n4701, n5007, n5780, n4979, n4978,
    n7359, n5203, n7722, n4721, n5029, n5075, n6787, n4554, n5777, n6878,
    n5698, n4494, n4507, n4488, n5520, n4493, n5716, n4487, n5714, n6510,
    n7312, n4484, n5402, n5709, n4403, n5590, n7678, n4540, n4483, n5594,
    n5390, n7465, n4869, n7454, n4543, n5498, n7238, n7616, n4782, n5737,
    n5729, n4867, n7624, n4416, n5497, n5516, n6860, n6870, n4958, n5496,
    n4844, n4779, n4830, n4913, n4686, n4820, n4806, n5559, n4852, n4829,
    n4720, n4634, n4684, n5513, n4749, n5494, n6688, n7629, n4390, n4384,
    n4608, n4393, n4984, n4557, n4411, n4449, n5581, n4432, n6123, n6130,
    n6985, n4741, n4763, n4839, n4908, n6573, n5051, n4740, n6085, n6502,
    n4716, n4714, n4854, n4754, n7175, n7173, n6997, n6569, n5018, n4864,
    n5178, n5174, n5162, n5059, n6444, n5147, n5050, n4905, n4792, n4817,
    n7786, n7774, n7782, n4766, n5287, n5294, n5284, n4676, n4880, n4884,
    n4841, n4842, n4617, n4969, n6916, n4997, n7100, n7050, n7108, n4655,
    n5624, n5727, n5708, n5713, n5692, n5696, n5895, n7282, n6797, n7065,
    n6612, n7335, n7327, n6932, n5186, n6905, n6655, n6653, n6662, n5165,
    n6563, n6458, n4732, n5962, n4743, n4903, n6333, n7406, n7405, n4923,
    n4947, n4831, n5315, n5320, n4723, n4717, n4724, n5633, n5735, n5504,
    n5907, n6095, n6318, n6512, n7627, n7625, n5066, n7758, n6527, n6237,
    n6249, n4911, n4828, n4729, n4606, n4719, n7805, n4870, n6087, n6148,
    n6146, n6505, n7621, n7077, n7204, n7088, n7083, n7004, n7193, n4878,
    n4814, n5293, n5270, n7207, n7208, n7029, n7192, n7581, n6892, n6744,
    n6650, n6373, n6163, n5042, n4865, n5259, n5256, n4745, n4582, n5234,
    n5219, n5222, n5223, n4944, n7515, n4645, n6267, n5533, n5249, n4609,
    n5135, n4495, n5290, n5313, n4922, n4924, n4907, n5771, n6144, n6308,
    n6361, n6684, n6862, n7391, n7457, n7520, n7300, n7303, n6895, n6714,
    n6651, n6791, n5062, n6288, n5056, n5055, n6295, n5754, n7721, n7730,
    n7734, n7653, n7648, n7589, n7571, n7597, n7434, n7428, n5283, n6934,
    n7306, n5089, n6942, n5189, n6894, n6721, n6782, n6649, n6568, n6576,
    n6400, n7043, n6406, n6447, n6279, n5150, n7005, n6223, n6161, n6102,
    n6038, n5656, n4485, n4381, n5505, n5510, n7807, n7349, n5787, n5789,
    n7792, n7814, n7811, n7818, n7783, n7784, n4748, n6208, n6207, n5749,
    n5663, n7417, n5296, n6918, n6554, n6954, n6427, n6429, n4593, n4620,
    n6829, n4973, n4971, n6828, n4502, n6014, n6011, n6633, n7116, n5322,
    n6919, n4930, n4823, n4797, n6063, n4572, n5563, n5558, n5593, n5589,
    n5782, n6432, n6156, n6352, n6676, n6872, n7382, n7468, n7540, n7795,
    n7596, n7705, n7558, n7322, n7284, n7476, n6648, n5170, n6647, n6847,
    n6625, n6450, n5157, n6452, n5159, n6421, n6289, n7830, n5886, n5128,
    n6983, n4654, n4481, n7824, n7831, n7679, n7671, n7477, n7370, n7326,
    n7341, n6975, n6976, n6879, n6906, n6806, n6637, n6600, n6586, n6587,
    n6398, n6517, n6378, n6385, n6384, n6322, n6324, n6238, n6182, n6185,
    n6052, n5981, n5969, n5875, n5854, n5950, n5954, n5535, n7239, n4392,
    n4391, n4957, n5318, n4889, n7354, n6334, n6767, n5022, n4887, n6250,
    n7410, n7409, n7407, n6528, n6705, n6699, n6006, n5841, n7266, n6557,
    n6959, n4529, n6831, n4975, n6830, n6021, n7695, n7694, n6634, n6990,
    n6133, n6834, n6654, n5879, n6022, n5991, n4406, n6353, n6689, n6867,
    n7673, n7497, n7251, n6825, n6775, n6790, n6844, n6606, n6414, n6416,
    n6548, n6340, n6233, n6276, n6257, n5745, n5946, n5944, n7761, n5831,
    n5808, n5383, n4439, n7236, n7176, n4417, n7115, n7622, n7463, n6868,
    n4522, n6508, n6314, n4781, n5767, n5704, n5722, n5600, n5726, n5571,
    n5622, n6077, n7821, n6158, n6320, n5978, n6060, n5986, n5919, n6057,
    n5989, n5916, n7649, n4579, n4567, n7184, n4378, n4607, n7009, n7139,
    n4765, n4856, n4783, n5210, n4637, n4946, n4770, n5173, n4503, n5100,
    n4952, n5819, n7311, n4448, n7232, n4380, n4379, n4382, n4383, n4386,
    n4385, n4387, n4635, n4660, n4730, n4414, n4395, n4407, n4404, n4401,
    n4399, n4427, n4398, n4400, n4402, n4405, n5395, n4408, n4410, n4409,
    n4413, n4412, n4419, n4418, n4421, n4420, n4423, n4422, n4425, n4424,
    n4438, n4429, n4428, n4431, n4434, n4433, n4437, n4443, n4441, n4440,
    n4446, n4445, n4447, n5506, n7631, n4450, n7636, n5401, n7725, n4454,
    n4452, n4453, n4456, n4455, n4460, n4458, n4457, n4459, n4482, n4462,
    n4461, n4463, n4480, n4465, n4464, n4469, n4467, n4466, n4468, n4477,
    n4471, n4470, n4475, n4473, n4472, n4474, n4476, n4478, n4479, n5387,
    n5468, n5469, n5471, n4499, n4497, n4498, n4500, n7794, n4521, n4516,
    n4511, n6125, n5324, n4513, n4517, n4518, n5583, n7790, n4519, n6498,
    n4520, n4531, n4525, n4523, n4524, n6395, n7700, n4530, n4902, n4538,
    n4535, n6627, n5657, n5211, n7772, n7542, n4547, n4550, n4548, n4551,
    n4552, n5924, n4562, n4560, n4558, n4559, n5190, n4561, n4563, n5641,
    n4565, n4564, n4592, n4569, n4568, n4570, n4573, n4571, n5662, n4583,
    n4578, n4576, n4577, n5658, n4581, n4580, n4588, n4586, n4585, n4587,
    n4590, n5639, n5614, n4596, n4599, n4597, n4598, n4605, n4600, n4603,
    n4601, n4602, n4604, n5794, n4613, n4662, n4611, n4610, n5124, n4612,
    n4616, n4615, n5617, n5786, n4624, n4626, n4627, n4628, n5927, n4641,
    n4639, n4638, n5759, n4640, n4644, n4643, n4649, n5845, n4653, n4652,
    n4656, n4664, n4661, n4663, n5847, n5998, n4680, n4688, n4687, n6000,
    n4700, n4706, n4704, n4705, n6074, n4722, n4805, n4734, n4733, n6206,
    n4750, n4757, n4756, n6202, n6268, n4774, n6224, n4785, n4784, n6264,
    n6270, n6332, n4801, n4798, n4808, n4807, n6335, n4827, n4824, n4833,
    n4832, n6280, n4843, n6476, n4848, n4858, n4857, n6470, n4872, n4871,
    n6539, n4904, n4897, n4894, n7788, n4899, n4910, n4987, n4916, n4915,
    n6562, n4926, n4925, n4934, n4931, n4938, n4937, n6700, n6917, n4953,
    n4963, n4962, n6924, n4976, n4977, n4980, n6915, n4991, n4985, n4990,
    n6792, n5002, n5006, n7267, n5013, n5011, n5010, n6722, n5012, n5016,
    n5021, n5020, n5039, n7697, n5037, n5025, n5023, n5072, n5027, n5033,
    n5035, n5034, n5036, n5038, n5040, n5043, n7188, n5929, n7185, n7180,
    n5044, n5741, n6718, n7286, n5180, n6893, n5071, n5069, n5073, n6904,
    n5082, n5083, n5084, n6943, n7046, n5093, n5092, n7720, n7424, n5109,
    n5098, n5099, n7503, n5107, n5106, n5108, n5117, n7037, n5120, n5122,
    n5921, n5922, n5125, n5742, n5127, n5130, n5134, n5960, n5138, n6036,
    n5140, n6114, n5143, n6171, n5146, n6221, n6371, n6402, n7045, n5167,
    n6597, n6778, n5188, n7740, n5938, n6780, n6754, n5192, n5194, n5329,
    n5276, n5300, n5319, n5201, n5204, n5202, n5205, n7696, n7657, n5212,
    n5215, n5243, n6955, n6957, n7350, n7305, n7352, n7518, n5263, n5264,
    n5265, n7522, n5274, n5291, n7367, n5279, n7325, n7473, n5304, n7573,
    n5308, n5311, n5317, n7806, n7664, n5325, n5337, n5335, n5333, n5331,
    n5330, n5332, n5334, n5336, n5338, n5341, n5340, n5343, n5342, n5345,
    n5344, n5347, n5346, n5349, n5348, n5351, n5350, n5353, n5352, n5355,
    n5354, n5357, n5356, n5359, n5358, n5361, n5360, n5363, n5362, n5365,
    n5364, n5367, n5366, n5369, n5368, n5371, n5370, n5373, n5372, n5375,
    n5374, n5377, n5376, n5378, n5380, n5379, n5382, n5384, n5386, n5385,
    n5389, n5399, n5394, n5391, n5393, n5398, n5397, n7181, n6987, n5403,
    n5408, n5476, n5404, n5405, n5406, n5407, n5410, n5409, n5411, n5413,
    n5412, n5415, n5414, n5417, n5416, n5419, n5418, n5421, n5420, n5423,
    n5422, n5425, n5424, n5432, n5427, n5426, n5430, n5428, n5429, n6992,
    n5431, n5440, n5435, n5433, n5434, n5438, n5437, n5439, n5442, n5441,
    n5444, n5443, n5446, n5445, n5448, n5447, n5450, n5449, n5452, n5451,
    n5454, n5453, n5456, n5455, n5458, n5457, n5460, n5459, n5462, n5461,
    n5464, n5463, n5482, n5480, n5472, n7755, n5473, n5478, n5475, n5477,
    n5483, n5479, n5485, n5484, n5487, n5486, n5489, n5488, n5491, n5490,
    n5493, n5492, n5564, n5509, n5768, n5507, n5511, n5508, n5528, n6064,
    n7235, n5512, n5522, n5523, n5524, n5526, n5525, n5527, n5531, n7637,
    n5530, n5651, n5541, n5576, n5539, n5537, n5536, n5538, n5540, n5544,
    n5542, n5543, n5545, n5552, n5550, n5547, n5546, n5548, n5549, n5551,
    n5554, n5553, n5556, n5555, n5561, n5560, n5575, n5566, n5565, n5570,
    n5568, n5567, n5569, n5573, n5572, n5574, n5588, n5580, n5577, n5578,
    n5579, n5582, n5585, n5584, n5587, n5605, n5592, n5591, n5604, n5596,
    n5595, n5599, n5834, n5597, n5598, n5602, n5601, n5603, n5606, n5608,
    n5607, n5612, n5610, n5609, n5611, n5619, n5615, n5616, n5618, n5621,
    n5620, n5631, n5629, n5625, n5627, n5628, n5630, n5638, n5634, n5636,
    n5637, n5642, n5643, n5650, n5644, n5646, n5645, n5648, n5647, n5649,
    n5653, n5652, n5655, n5654, n5683, n5661, n5659, n5682, n5660, n5675,
    n5665, n5664, n5672, n5667, n5668, n5670, n5669, n5671, n5674, n5673,
    n5681, n5676, n5678, n5677, n5680, n5679, n5687, n5685, n5684, n5688,
    n5686, n5690, n5689, n6023, n5691, n5703, n5693, n5695, n5701, n5697,
    n5699, n5700, n5702, n5706, n5705, n5992, n5707, n5721, n5710, n5712,
    n5719, n5715, n5717, n5718, n5720, n5724, n5723, n5795, n5725, n5734,
    n5732, n5728, n5730, n5731, n5733, n5740, n5736, n5738, n5739, n5746,
    n5744, n5801, n5743, n5765, n5753, n5748, n5747, n5751, n5750, n5752,
    n5758, n5756, n5757, n5805, n5760, n5761, n5802, n5762, n5763, n5764,
    n6197, n5766, n5776, n5774, n5890, n5770, n5772, n5773, n5775, n5785,
    n5781, n5783, n5784, n5788, n5793, n5791, n5790, n5792, n5800, n5798,
    n5796, n5797, n5799, n5807, n5803, n5804, n5806, n5810, n5809, n5830,
    n5813, n5812, n5857, n5824, n5815, n5823, n5818, n5817, n5821, n5820,
    n5822, n5828, n5864, n5827, n5829, n5833, n5832, n5838, n5836, n5835,
    n5837, n5840, n5839, n5843, n5842, n5850, n5846, n5848, n5849, n5852,
    n5851, n5853, n5855, n5863, n5859, n7750, n5858, n5861, n5860, n5862,
    n5866, n5865, n5868, n5867, n5885, n5870, n5873, n5872, n5874, n5877,
    n5878, n5881, n5880, n5911, n5882, n5883, n5884, n5888, n5913, n5887,
    n6262, n5889, n5900, n5898, n5893, n5896, n6082, n5897, n5899, n5910,
    n5905, n5908, n5909, n5917, n5915, n5914, n5920, n5923, n5936, n5926,
    n5925, n5934, n5932, n5930, n5931, n5933, n5935, n5939, n5941, n5952,
    n5942, n5943, n5947, n5945, n5949, n5948, n5956, n5951, n5953, n5957,
    n5955, n5959, n5958, n5970, n5964, n5963, n5967, n5966, n5968, n5977,
    n5972, n5973, n5984, n5975, n5974, n5976, n5980, n5979, n5987, n5983,
    n5990, n5993, n6005, n5996, n5995, n6003, n5999, n6001, n6002, n6004,
    n6008, n6007, n6010, n6009, n6013, n6015, n6020, n6018, n6017, n6019,
    n6028, n6026, n6024, n6025, n6027, n6031, n6051, n6035, n6033, n6032,
    n6034, n6050, n6046, n6044, n6040, n6039, n6042, n6041, n6043, n6048,
    n6047, n6049, n6058, n6054, n6053, n6055, n6061, n6072, n6065, n6067,
    n6066, n6070, n6069, n6071, n6078, n6075, n6076, n6080, n6079, n6342,
    n6081, n6090, n6088, n6139, n6084, n6086, n6140, n6089, n6098, n6094,
    n6096, n6097, n6100, n6099, n6118, n6103, n6106, n6105, n6107, n6111,
    n6112, n6253, n6115, n6121, n6137, n6124, n6129, n6126, n6128, n6132,
    n6131, n6135, n6136, n6138, n6149, n6147, n6143, n6142, n6145, n6305,
    n6159, n6154, n6157, n6178, n6170, n6167, n6165, n6164, n6166, n6168,
    n6173, n6174, n6181, n6190, n6183, n6186, n6191, n6195, n6194, n6198,
    n6213, n6201, n6200, n6211, n6209, n6205, n6210, n6214, n6220, n6218,
    n6217, n6219, n6236, n6228, n6226, n6225, n6227, n6229, n6244, n6239,
    n6247, n6248, n6251, n6254, n6256, n6259, n6263, n6275, n6266, n6265,
    n6273, n6269, n6271, n6277, n6287, n6282, n6283, n6284, n6294, n6292,
    n6291, n6293, n6297, n6302, n6469, n6304, n6313, n6311, n6356, n6358,
    n6348, n6317, n6319, n6328, n6331, n6337, n6336, n6338, n6345, n6343,
    n6344, n6346, n6351, n6509, n6541, n6360, n6499, n6365, n6369, n6389,
    n6375, n6374, n6376, n6531, n6392, n6394, n6393, n6485, n6399, n6412,
    n6401, n6489, n6408, n6418, n6435, n6431, n6425, n6437, n6463, n6446,
    n6445, n6451, n6524, n6466, n6468, n6482, n6473, n6472, n6480, n6553,
    n6477, n6483, n6493, n6496, n6497, n6507, n6679, n6681, n6672, n6523,
    n6518, n6529, n6532, n6537, n6547, n6542, n6545, n6544, n6546, n6561,
    n6550, n6556, n6567, n6565, n6564, n6566, n6585, n6575, n6574, n6578,
    n6593, n6596, n6604, n6611, n6609, n6608, n6610, n6614, n6619, n6623,
    n6622, n6631, n6626, n6629, n6628, n6630, n6636, n6643, n6646, n6668,
    n6849, n6671, n6675, n6869, n6683, n6859, n6693, n6697, n6702, n6701,
    n6703, n6709, n6707, n6858, n6708, n6710, n6715, n6741, n6717, n6726,
    n6724, n6723, n6725, n6727, n6735, n6738, n6888, n6746, n6749, n6748,
    n6751, n6750, n6752, n6759, n6762, n6766, n6768, n6769, n6773, n6776,
    n6796, n6794, n6793, n6795, n6804, n6812, n6815, n6821, n6841, n6839,
    n6837, n6835, n7452, n6836, n6838, n6840, n6842, n6855, n6857, n7386,
    n7378, n6884, n6882, n6885, n6899, n6897, n6896, n6898, n6900, n6909,
    n6912, n6929, n7280, n6936, n6935, n6939, n6938, n6971, n6945, n7281,
    n6951, n6949, n6952, n6956, n6970, n6968, n6961, n6960, n6963, n6962,
    n6966, n6965, n6967, n6969, n6972, n6977, n6979, n6989, n7500, n7216,
    n6986, n6991, n7221, n7099, n6988, n6998, n7724, n7106, n6993, n7219,
    n6994, n7748, n6995, n7780, n7000, n7137, n7002, n7027, n7006, n7023,
    n7194, n7012, n7147, n7018, n7014, n7016, n7017, n7019, n7021, n7022,
    n7025, n7026, n7028, n7572, n7331, n7321, n7438, n7033, n7035, n7049,
    n7039, n7040, n7042, n7044, n7047, n7048, n7075, n7076, n7098, n7107,
    n7109, n7110, n7118, n7210, n7127, n7122, n7165, n7128, n7126, n7157,
    n7129, n7163, n7131, n7135, n7134, n7142, n7202, n7141, n7154, n7146,
    n7145, n7152, n7150, n7151, n7153, n7155, n7156, n7172, n7160, n7161,
    n7164, n7170, n7167, n7169, n7171, n7179, n7183, n7182, n7187, n7186,
    n7191, n7189, n7190, n7200, n7195, n7197, n7198, n7199, n7206, n7203,
    n7205, n7222, n7237, n7241, n7240, n7242, n7243, n7247, n7248, n7260,
    n7263, n7279, n7277, n7272, n7270, n7269, n7271, n7275, n7274, n7276,
    n7278, n7292, n7332, n7295, n7294, n7302, n7309, n7318, n7316, n7319,
    n7324, n7437, n7441, n7429, n7340, n7338, n7337, n7339, n7366, n7346,
    n7344, n7347, n7351, n7365, n7363, n7358, n7356, n7355, n7357, n7361,
    n7360, n7362, n7364, n7373, n7372, n7390, n7453, n7401, n7421, n7413,
    n7412, n7416, n7415, n7419, n7418, n7420, n7422, n7426, n7425, n7427,
    n7584, n7472, n7440, n7507, n7448, n7446, n7449, n7451, n7456, n7480,
    n7479, n7487, n7488, n7494, n7499, n7510, n7505, n7502, n7723, n7536,
    n7669, n7749, n7539, n7513, n7516, n7553, n7524, n7523, n7529, n7528,
    n7534, n7545, n7537, n7541, n7548, n7568, n7566, n7564, n7562, n7561,
    n7563, n7565, n7567, n7569, n7588, n7576, n7577, n7578, n7659, n7605,
    n7580, n7591, n7642, n7610, n7594, n7600, n7601, n7613, n7611, n7614,
    n7618, n7638, n7712, n7654, n7652, n7651, n7684, n7672, n7687, n7685,
    n7688, n7709, n7704, n7702, n7701, n7703, n7707, n7706, n7708, n7710,
    n7719, n7728, n7727, n7729, n7762, n7737, n7738, n7756, n7741, n7742,
    n7745, n7744, n7760, n7768, n7766, n7765, n7771, n7770, n7773, n7781,
    n7787, n7803, n7801, n7799, n7797, n7796, n7798, n7800, n7802, n7804,
    n7822, n7809, n7820, n7816, n7817, n7819, n7828, n7836;
  assign n7769 = ~n5482 | ~n5471;
  assign n7764 = ~n5482 | ~n5481;
  assign n7743 = ~n7832;
  assign n7056 = ~n5058 & ~n7159;
  assign n5826 = ~n5127 | ~n5126;
  assign n7777 = ~n5211 & ~n7542;
  assign n5209 = ~n4584 | ~n4540;
  assign n5392 = n4398 ^ IR_REG_26__SCAN_IN;
  assign n6996 = ~n6985;
  assign n6127 = ~n4511 | ~n4507;
  assign n7501 = ~n4430 ^ IR_REG_27__SCAN_IN;
  assign n4415 = ~n4411 | ~IR_REG_31__SCAN_IN;
  assign n4506 = n4444 ^ n5381;
  assign n4444 = ~n5383 | ~IR_REG_31__SCAN_IN;
  assign n4633 = ~IR_REG_2__SCAN_IN;
  assign n4948 = ~n6698 & ~n6695;
  assign n4396 = ~IR_REG_22__SCAN_IN;
  assign n6698 = ~n4926 | ~n4925;
  assign n5436 = ~n6127;
  assign n7746 = ~n5113 | ~n5465;
  assign n4584 = ~n5392 | ~n4403;
  assign n7533 = ~n5282 | ~n5281;
  assign n6832 = ~n4956 | ~n4955;
  assign n6422 = ~n4801 | ~n4800;
  assign n7767 = ~n7769;
  assign n7763 = ~n7764;
  assign n6193 = n4584 | n4406;
  assign n7595 = ~n7610 | ~n7743;
  assign n7677 = ~n7666 | ~n7665;
  assign n7666 = ~n7684 | ~n7743;
  assign n7676 = ~n7675 & ~n7674;
  assign n7683 = ~n7682 & ~n7681;
  assign n7593 = ~n7591 | ~n7590;
  assign n7609 = ~n7608 & ~n7607;
  assign n7603 = ~n7602 & ~n7601;
  assign n7450 = ~n7448 | ~n7767;
  assign n7608 = ~n7605 & ~n7678;
  assign n7602 = ~n7605 & ~n7667;
  assign n7447 = ~n7448 | ~n7763;
  assign n7320 = ~n7318 | ~n7763;
  assign n7317 = ~n7318 | ~n7767;
  assign n7483 = ~n7482 & ~n7481;
  assign n7345 = ~n7346 | ~n7763;
  assign n7348 = ~n7346 | ~n7767;
  assign n7495 = ~n7493 & ~n7492;
  assign n7444 = ~n7477 & ~n7755;
  assign n7482 = ~n7477 & ~n7476;
  assign n7256 = ~n7253 & ~n7252;
  assign n7556 = ~n7555 | ~n7554;
  assign n7376 = ~n7375 & ~n7374;
  assign n7690 = ~n5299 & ~n5298;
  assign n7314 = ~n7311 & ~n7486;
  assign n6913 = ~n6911 | ~n7767;
  assign n7330 = ~n7370 & ~n7755;
  assign n7375 = ~n7370 & ~n7476;
  assign n6910 = ~n6911 | ~n7763;
  assign n7554 = ~n7553 | ~n7552;
  assign n7253 = ~n7251 & ~n7250;
  assign n7492 = ~n7491 | ~n7490;
  assign n7519 = ~n7516 & ~n7813;
  assign n6886 = ~n6884 | ~n7763;
  assign n6883 = ~n6884 | ~n7767;
  assign n6911 = ~n7245 | ~n6908;
  assign n7304 = ~n7302 | ~n7301;
  assign n7353 = ~n7351 & ~n7813;
  assign n7498 = ~n7497 | ~n7496;
  assign n7313 = ~n7497 | ~n7312;
  assign n7423 = ~n7409 | ~n7808;
  assign n6982 = ~n6973 | ~n6972;
  assign n7732 = ~n7721 & ~n7720;
  assign n7245 = ~n6903 & ~n6902;
  assign n6907 = ~n7254 & ~n7678;
  assign n7255 = ~n7254 & ~n7667;
  assign n7484 = ~n7475 | ~n7474;
  assign n6760 = ~n6761 | ~n7763;
  assign n6903 = ~n7254 & ~n7661;
  assign n6973 = ~n6971 | ~n7743;
  assign n6763 = ~n6761 | ~n7767;
  assign n6981 = ~n6980 & ~n6979;
  assign n6881 = ~n6877 & ~n6876;
  assign n7265 = ~n7262 | ~n7808;
  assign n6739 = ~n6737 | ~n7767;
  assign n7475 = ~n7472 | ~n7743;
  assign n6736 = ~n6737 | ~n7763;
  assign n6777 = ~n6774 | ~n6773;
  assign n6947 = ~n6975 & ~n7755;
  assign n7377 = ~n7369 | ~n7368;
  assign n6761 = ~n6758 | ~n6757;
  assign n6877 = ~n5111 | ~n5110;
  assign n6811 = ~n7767 | ~n6813;
  assign n6805 = ~n7743 | ~n6803;
  assign n6958 = ~n6956 & ~n7813;
  assign n6980 = ~n6975 & ~n7476;
  assign n6814 = ~n7763 | ~n6813;
  assign n7262 = ~n7264 | ~n7263;
  assign n6774 = ~n6772 | ~n6771;
  assign n7404 = ~n7264 & ~n7263;
  assign n6758 = ~n6825 | ~n6878;
  assign n6803 = ~n6802 | ~n6810;
  assign n6737 = ~n6772 | ~n6734;
  assign n5198 = ~n5197 | ~n5196;
  assign n6941 = ~n6934 & ~n7720;
  assign n6891 = ~n6890 | ~n6889;
  assign n7369 = ~n7366 | ~n7743;
  assign n7715 = ~n7713 & ~n7712;
  assign n6813 = ~n6810 | ~n6809;
  assign n5041 = ~n5022 & ~n7813;
  assign n6802 = ~n6787 & ~n6786;
  assign n6810 = ~n6801 & ~n6800;
  assign n6930 = ~n7395 & ~n6927;
  assign n7264 = ~n7260 | ~n7259;
  assign n6772 = ~n6730 & ~n6729;
  assign n6734 = ~n6733 & ~n6732;
  assign n6827 = ~n6824 & ~n6823;
  assign n6800 = ~n6799 | ~n6798;
  assign n7112 = ~n7111 | ~n7110;
  assign n6824 = ~n6818 & ~n6817;
  assign n6730 = ~n6775 & ~n7661;
  assign n5091 = ~n5089 | ~n7046;
  assign n6927 = ~n6926 | ~n6925;
  assign n6786 = ~n6785 | ~n6784;
  assign n6933 = ~n6931 | ~n7084;
  assign n6852 = ~n6851 & ~n6850;
  assign n6743 = ~n6741 & ~n6740;
  assign n6809 = ~n6808 & ~n6807;
  assign n6667 = ~n7767 | ~n6669;
  assign n6798 = ~n6797 | ~n5472;
  assign n6843 = ~n6830 | ~n7808;
  assign n6670 = ~n7763 | ~n6669;
  assign n6926 = ~n6923 & ~n6922;
  assign n7111 = ~n7105 | ~n7104;
  assign n6931 = ~n5090 | ~n5189;
  assign n7587 = ~n7585 & ~n7584;
  assign n6642 = ~n7763 | ~n6644;
  assign n6669 = ~n6666 | ~n6849;
  assign n6922 = ~n6921 | ~n6920;
  assign n6620 = ~n7743 | ~n6618;
  assign n7291 = ~n7300 & ~n7720;
  assign n7334 = ~n7429 & ~n7333;
  assign n5090 = ~n5079 | ~n5078;
  assign n6901 = ~n6894 | ~n7647;
  assign n7105 = ~n7101 & ~n7100;
  assign n6851 = ~n6848 | ~n6847;
  assign n6645 = ~n7767 | ~n6644;
  assign n6618 = ~n6617 | ~n6641;
  assign n5079 = ~n6893 | ~n6892;
  assign n6753 = ~n6747 | ~n7647;
  assign n7101 = ~n7097 & ~n7096;
  assign n6921 = ~n6918 | ~n7808;
  assign n6848 = ~n6846 & ~n6845;
  assign n6492 = ~n7763 | ~n6494;
  assign n6854 = ~n6844 & ~n7667;
  assign n6617 = ~n6604 & ~n6603;
  assign n6661 = ~n6844 & ~n7755;
  assign n6729 = ~n6728 | ~n6727;
  assign n6711 = ~n6704 & ~n6703;
  assign n6747 = ~n6746 | ~n6745;
  assign n6495 = ~n7767 | ~n6494;
  assign n6595 = ~n7767 | ~n6594;
  assign n6584 = ~n6583 & ~n6582;
  assign n6603 = ~n6602 | ~n6601;
  assign n7290 = ~n7286 | ~n7285;
  assign n6728 = ~n6721 | ~n7647;
  assign n6592 = ~n7763 | ~n6594;
  assign n6704 = ~n6699 & ~n7813;
  assign n7095 = ~n7094 & ~n7586;
  assign n6615 = ~n6614 | ~n6613;
  assign n6745 = ~n7286 | ~n6744;
  assign n6640 = ~n6639 & ~n6638;
  assign n7094 = ~n7585 & ~n7092;
  assign n6420 = ~n6413 | ~n7743;
  assign n6491 = ~n6488 & ~n6487;
  assign n6594 = ~n6591 | ~n6590;
  assign n6526 = ~n6523 & ~n6522;
  assign n6591 = ~n6581 & ~n6580;
  assign n6657 = ~n6656 | ~n6655;
  assign n6413 = ~n6412 | ~n6486;
  assign n6720 = ~n6718 | ~n6717;
  assign n6487 = ~n6486 | ~n6485;
  assign n7092 = ~n7430 & ~n7091;
  assign n6635 = ~n6634 | ~n7808;
  assign n6419 = ~n6418 & ~n6417;
  assign n5067 = ~n6718 | ~n7121;
  assign n6522 = ~n6521 | ~n6520;
  assign n6801 = ~n6790 & ~n7720;
  assign n6521 = ~n6519 & ~n6518;
  assign n6656 = ~n6653 | ~n7647;
  assign n6590 = ~n6589 & ~n6588;
  assign n6580 = ~n6579 | ~n6578;
  assign n5168 = ~n6597;
  assign n6538 = ~n6536 | ~n7743;
  assign n6417 = ~n6416 | ~n6415;
  assign n7091 = n7090 & n7089;
  assign n6411 = n6489 & n5472;
  assign n6490 = ~n6489 | ~n7312;
  assign n6536 = ~n6535 | ~n6534;
  assign n6579 = ~n6577 & ~n6576;
  assign n6581 = ~n6586 & ~n7661;
  assign n4901 = ~n4900 | ~n4899;
  assign n6534 = ~n6533 & ~n6532;
  assign n4900 = ~n4889 | ~n7808;
  assign n6616 = ~n6606 & ~n7720;
  assign n6484 = ~n6482 & ~n6481;
  assign n7080 = ~n7078 | ~n7119;
  assign n6560 = ~n6559 & ~n6558;
  assign n6652 = ~n6651 & ~n6650;
  assign n6577 = ~n6573 & ~n7720;
  assign n6481 = ~n6480 | ~n6479;
  assign n6403 = ~n6401 | ~n7043;
  assign n6461 = ~n6460 & ~n6459;
  assign n6533 = ~n6530 | ~n6529;
  assign n6455 = ~n6454 | ~n6453;
  assign n7544 = ~n7763 | ~n7546;
  assign n7547 = ~n7767 | ~n7546;
  assign n6438 = ~n6435 & ~n6434;
  assign n6558 = ~n6557 & ~n7813;
  assign n6479 = ~n6478 | ~n6477;
  assign n7509 = ~n7763 | ~n7511;
  assign n7546 = ~n7823 | ~n7543;
  assign n6434 = ~n6433 | ~n6432;
  assign n6572 = ~n6571 | ~n7059;
  assign n7512 = ~n7767 | ~n7511;
  assign n7827 = ~n7826 | ~n7825;
  assign n6525 = ~n6524 | ~n7496;
  assign n6460 = n6524 & n7312;
  assign n6410 = ~n6409 | ~n6408;
  assign n6454 = ~n6448 & ~n6447;
  assign n6409 = ~n6406 | ~n7647;
  assign n7835 = ~n7834 | ~n7833;
  assign n7511 = ~n7829 | ~n7508;
  assign n6380 = ~n6379 | ~n6378;
  assign n6448 = ~n6444 & ~n7720;
  assign n6555 = ~n6554 & ~n6553;
  assign n5064 = ~n6570 | ~n7130;
  assign n7674 = ~n7673 | ~n7672;
  assign n7825 = ~n7824 | ~n7830;
  assign n7069 = ~n7067 & ~n7066;
  assign n6433 = ~n6431 & ~n6430;
  assign n7753 = ~n7752 & ~n7751;
  assign n6430 = ~n6429 | ~n6428;
  assign n7067 = ~n7063 & ~n7062;
  assign n6301 = ~n6300 | ~n6326;
  assign n6379 = ~n6377 & ~n6376;
  assign n7834 = ~n7831 | ~n7830;
  assign n6329 = ~n6326 | ~n6325;
  assign n7681 = ~n7680 & ~n7757;
  assign n6570 = ~n6405;
  assign n7607 = ~n7606 & ~n7757;
  assign n7481 = ~n7480 | ~n7479;
  assign n6387 = n6531 & n6386;
  assign n7471 = ~n7462 & ~n7461;
  assign n7759 = ~n7758 & ~n7757;
  assign n6443 = ~n6442 | ~n6441;
  assign n7063 = ~n7061 & ~n7060;
  assign n6300 = ~n6287 & ~n6286;
  assign n6326 = ~n6299 & ~n6298;
  assign n7751 = ~n7758 & ~n7750;
  assign n6377 = ~n6373 & ~n7720;
  assign n7374 = ~n7373 | ~n7372;
  assign n7443 = ~n7478 & ~n7757;
  assign n5061 = ~n7056 | ~n5059;
  assign n7606 = ~n7598 | ~n7669;
  assign n6234 = ~n6233 | ~n6242;
  assign n6245 = ~n6242 | ~n6241;
  assign n6192 = ~n6190 & ~n6189;
  assign n6298 = ~n6297 | ~n6296;
  assign n7461 = ~n7460 | ~n7459;
  assign n6381 = n6527 & n5472;
  assign n6347 = ~n6339 & ~n6338;
  assign n6299 = ~n6289 & ~n7720;
  assign n7490 = n7489 & n7488;
  assign n7329 = ~n7371 & ~n7757;
  assign n6325 = ~n6324 & ~n6323;
  assign n6242 = ~n6232 & ~n6231;
  assign n6278 = ~n6275 & ~n6274;
  assign n7399 = ~n7398 | ~n7397;
  assign n7459 = ~n7458 | ~n7623;
  assign n7470 = ~n7469 | ~n7617;
  assign n6426 = ~n4819 | ~n4818;
  assign n7230 = ~n7229 | ~n7228;
  assign n7469 = ~n7466 & ~n7620;
  assign n6188 = ~n6187 & ~n6186;
  assign n6231 = ~n6230 | ~n6229;
  assign n6274 = ~n6273 | ~n6272;
  assign n7458 = ~n7455 & ~n7628;
  assign n7398 = ~n7396 & ~n7395;
  assign n7400 = ~n7385 & ~n7384;
  assign n7623 = ~n7457 | ~n7456;
  assign n6179 = ~n6184 | ~n6176;
  assign n7466 = ~n7467 & ~n7468;
  assign n6875 = ~n6867 & ~n6866;
  assign n7396 = ~n7394 & ~n7393;
  assign n6215 = ~n6213 & ~n6212;
  assign n7227 = ~n7225;
  assign n6241 = ~n6240 & ~n6239;
  assign n6272 = ~n6271 | ~n6270;
  assign n7455 = ~n7456 & ~n7457;
  assign n5154 = ~n6279 | ~n5152;
  assign n5196 = ~n5195 & ~n5194;
  assign n6866 = ~n6865 | ~n6864;
  assign n7467 = ~n7465 | ~n7464;
  assign n6184 = ~n6169 & ~n6168;
  assign n5057 = ~n6222 | ~n5055;
  assign n5195 = n6876 & n6819;
  assign n6119 = ~n6252 | ~n6116;
  assign n7393 = ~n7453 | ~n7392;
  assign n7225 = ~n7223 | ~n7222;
  assign n6176 = ~n6175 & ~n6182;
  assign n7223 = ~n7220 | ~n7219;
  assign n6946 = ~n6976 & ~n7757;
  assign n7250 = ~n7249 | ~n7248;
  assign n7464 = ~n7382 | ~n7381;
  assign n6169 = ~n6161 & ~n7720;
  assign n6823 = ~n6822 | ~n6821;
  assign n6874 = ~n6873 | ~n7379;
  assign n6252 = ~n6108 & ~n6107;
  assign n6864 = ~n6863 | ~n7388;
  assign n7394 = ~n7391 & ~n7390;
  assign n6694 = ~n6692 & ~n6691;
  assign n6691 = ~n6690 | ~n6689;
  assign n6863 = ~n6861 & ~n7628;
  assign n7220 = ~n7218 | ~n7217;
  assign n7381 = ~n7380 | ~n7379;
  assign n6108 = ~n6104 | ~n6103;
  assign n6873 = ~n6871 & ~n7620;
  assign n5054 = ~n6160 & ~n7148;
  assign n6059 = ~n6056 | ~n6055;
  assign n6160 = ~n5053 | ~n6999;
  assign n7218 = ~n7214 | ~n7213;
  assign n6771 = ~n6770 & ~n6769;
  assign n6056 = ~n6046 & ~n6045;
  assign n7246 = ~n6906 & ~n7757;
  assign n6116 = ~n6253 & ~n6115;
  assign n6690 = ~n6688 & ~n6687;
  assign n5988 = ~n5985 | ~n5984;
  assign n6515 = ~n6507 & ~n6506;
  assign n6692 = ~n6678 & ~n6677;
  assign n7389 = ~n7387 | ~n7386;
  assign n7380 = ~n7387 | ~n7378;
  assign n6770 = ~n6766 & ~n6765;
  assign n6687 = ~n6686 & ~n6685;
  assign n6732 = ~n6765 & ~n6764;
  assign n4768 = ~n6206 | ~n4745;
  assign n6506 = ~n6505 | ~n6504;
  assign n5985 = ~n5983 & ~n5982;
  assign n7211 = ~n7210 & ~n7209;
  assign n6504 = ~n6503 | ~n6681;
  assign n6370 = ~n6368 & ~n6367;
  assign n6513 = ~n6511 & ~n7620;
  assign n7052 = ~n7051 & ~n7050;
  assign n6503 = ~n6501 & ~n7628;
  assign n6639 = n6600 & n6599;
  assign n6367 = ~n6366 | ~n6365;
  assign n7209 = ~n7208 & ~n7207;
  assign n7051 = ~n7032 | ~n7716;
  assign n6673 = ~REG2_REG_14__SCAN_IN | ~n6512;
  assign n6366 = ~n6541 & ~n6364;
  assign n6588 = ~n6587 & ~n7757;
  assign n6682 = ~n6680 | ~n6679;
  assign n6674 = ~n6680 | ~n6672;
  assign n6364 = ~n6363 & ~n6362;
  assign n6368 = ~n6354 & ~n6353;
  assign n6321 = ~n6313 & ~n6312;
  assign n6598 = ~n6562 | ~n6563;
  assign n6312 = ~n6311 | ~n6310;
  assign n7031 = ~n7030 | ~n7029;
  assign n6459 = ~n6517 & ~n7757;
  assign n6396 = ~n6539 | ~n6458;
  assign n6309 = ~n6307 & ~n7628;
  assign n5046 = ~n5814;
  assign n7217 = ~n7216 & ~n7215;
  assign n6349 = ~REG2_REG_12__SCAN_IN | ~n6318;
  assign n7030 = ~n6998 & ~n6997;
  assign n7104 = ~n7215;
  assign n6359 = ~n6357 | ~n6356;
  assign n6383 = ~n6280 | ~n6281;
  assign n7215 = ~n7103 | ~n7716;
  assign n6350 = ~n6357 | ~n6348;
  assign n5242 = ~n5241 & ~n5240;
  assign n5241 = ~n5237 & ~n5236;
  assign n6281 = ~n6335 & ~n6216;
  assign n7660 = ~n7641 | ~n7640;
  assign n5045 = ~n5755 | ~n5741;
  assign n7097 = ~n7102;
  assign n7555 = ~n7550 | ~n7549;
  assign n5218 = ~n7786;
  assign n5217 = ~n7785;
  assign n7655 = ~n7654 & ~n7653;
  assign n7517 = ~n7515 & ~n7551;
  assign n6216 = ~n6172 | ~n6264;
  assign n7641 = ~n7714;
  assign n7691 = ~n5316 | ~n5315;
  assign n7102 = ~n7717 & ~n7714;
  assign n7713 = ~n7640 | ~n7644;
  assign n4881 = ~n6549 | ~n6552;
  assign n5298 = ~n5297 | ~n7549;
  assign n6315 = ~n6156 | ~n6155;
  assign n5237 = ~n5235 & ~n7403;
  assign n7552 = ~n7551;
  assign n7692 = ~n5313 | ~n5314;
  assign n7776 = ~n7774 | ~n7773;
  assign n6073 = ~n6203 & ~n4744;
  assign n6204 = ~n4769 & ~n4767;
  assign n7592 = ~n7733 & ~n7649;
  assign n7436 = ~n7428 | ~n7427;
  assign n7549 = ~n5296 | ~n5295;
  assign n7785 = ~n5216 | ~n5215;
  assign n7731 = ~n7730 | ~n7729;
  assign n6172 = ~n6110 & ~n6109;
  assign n7640 = ~n7733 | ~n7780;
  assign n7257 = ~n7259 | ~n5232;
  assign n7714 = ~n7733 & ~n7780;
  assign n5844 = ~n4675 & ~n4674;
  assign n7735 = ~n7733 & ~n7792;
  assign n5613 = ~n4622 & ~n4621;
  assign n6155 = ~n6153 | ~n6152;
  assign n5235 = ~n5232 & ~n7261;
  assign n6696 = ~n4947 & ~n4946;
  assign n5184 = ~n5183 & ~n5182;
  assign n5230 = ~n5229 & ~n5236;
  assign n4909 = ~n4908 | ~n4907;
  assign n4972 = ~n4971 | ~n4970;
  assign n6552 = ~n4880 | ~n4879;
  assign n4648 = ~n4647 & ~n4646;
  assign n5214 = ~n5213 & ~n5212;
  assign n4623 = ~n4622;
  assign n4818 = ~n4817 | ~n4816;
  assign n6549 = ~n4884 | ~n4883;
  assign n4744 = ~n4743 & ~n4742;
  assign n4715 = ~n4714 & ~n6011;
  assign n6424 = ~n4839 & ~n4840;
  assign n4767 = ~n4766 & ~n4765;
  assign n6474 = ~n4878 | ~n4864;
  assign n4621 = ~n4620 & ~n4619;
  assign n7717 = ~n7789 & ~n7748;
  assign n7716 = ~n7789 | ~n7748;
  assign n4674 = ~n4673 & ~n4672;
  assign n5229 = ~n7259 | ~n5231;
  assign n7643 = ~n7791 | ~n7506;
  assign n5232 = ~n5021 | ~n5020;
  assign n7551 = ~n5293 & ~n5292;
  assign n7514 = ~n5293 | ~n5292;
  assign n7658 = ~n7791 | ~n7657;
  assign n6404 = ~n6569 | ~n7059;
  assign n7289 = ~n7288 & ~n7287;
  assign n5176 = ~n6714 & ~n5175;
  assign n5183 = ~n5179 & ~n5178;
  assign n7733 = ~n7778;
  assign n5001 = ~n5000 | ~n4999;
  assign n7575 = ~n7574 | ~n7573;
  assign n5260 = ~n5259 | ~n5258;
  assign n5310 = ~n5309 | ~n5308;
  assign n6372 = ~n6440 | ~n6441;
  assign n7778 = ~n5328 | ~n5327;
  assign n4675 = ~n4670 & ~n4671;
  assign n4696 = ~n4695 | ~n4694;
  assign n5314 = ~n5312 | ~n5311;
  assign n5252 = ~n5251 | ~n5250;
  assign n4906 = ~n4546 & ~n4545;
  assign n4816 = ~n4815;
  assign n4712 = ~n6012 & ~n4713;
  assign n7586 = ~n7093;
  assign n4793 = ~n4792 | ~n4791;
  assign n5063 = ~n5164 & ~n7059;
  assign n5060 = ~n7158 | ~n5158;
  assign n7582 = ~n7581 | ~n7580;
  assign n4769 = ~n4763 & ~n4764;
  assign n7791 = ~n7696;
  assign n6799 = ~n6796 & ~n6795;
  assign n7034 = ~n7065 | ~n7124;
  assign n5289 = ~n5295;
  assign n7003 = ~n7132 & ~n7149;
  assign n5240 = ~n5239 & ~n7405;
  assign n6141 = ~n6151 | ~n6139;
  assign n6153 = ~n6151 | ~n6150;
  assign n5175 = ~n5174 | ~n6887;
  assign n4622 = ~n4618 & ~n4617;
  assign n4945 = ~n4943 & ~n4942;
  assign n7525 = ~n7524 & ~n7523;
  assign n7789 = ~n6134 & ~n6133;
  assign n4647 = ~n4645;
  assign n7288 = ~n7168 & ~n7087;
  assign n7261 = ~n5231;
  assign n5179 = ~n6740 & ~n5177;
  assign n4591 = ~n5534 & ~n5533;
  assign n7020 = ~n6647 | ~n7120;
  assign n6203 = ~n4741 & ~n4740;
  assign n5000 = ~n4997;
  assign n5295 = ~n5288 | ~n5287;
  assign n5286 = ~n5285 | ~n5284;
  assign n7068 = ~n7124 | ~n7120;
  assign n4919 = ~n4918 | ~n4917;
  assign n4966 = ~n4965 | ~n4964;
  assign n5273 = ~n5271 | ~n5270;
  assign n4943 = ~n6649 & ~n5015;
  assign n7333 = ~n7054;
  assign n5292 = n5275 & n5274;
  assign n4546 = ~n6540 & ~n5015;
  assign n6719 = ~n7074 & ~n7072;
  assign n5148 = ~n6290 | ~n5147;
  assign n4970 = ~n4968 | ~n4967;
  assign n4544 = ~n4542 | ~n4541;
  assign n4883 = ~n4877 | ~n4876;
  assign n7430 = ~n7055 | ~n7054;
  assign n7168 = ~n7086 & ~n7085;
  assign n7574 = ~n7579;
  assign n7439 = ~n7698 | ~n7559;
  assign n4875 = ~n4874 | ~n4873;
  assign n4999 = ~n4998;
  assign n5251 = ~n5249;
  assign n4879 = ~n4863 | ~n4862;
  assign n5825 = ~n7007 | ~n7196;
  assign n4861 = ~n4860 | ~n4859;
  assign n5239 = ~n7406;
  assign n5236 = ~n7406 & ~n5238;
  assign n7431 = ~n7698 | ~n7325;
  assign n4840 = ~n4838 | ~n4837;
  assign n5160 = ~n6471 | ~n6539;
  assign n4836 = ~n4835 | ~n4834;
  assign n5231 = ~n5234 | ~n5233;
  assign n4815 = ~n4813 | ~n4812;
  assign n4791 = ~n4790 | ~n4789;
  assign n7403 = ~n5234 & ~n5233;
  assign n7530 = ~n7529 | ~n7528;
  assign n4811 = ~n4810 | ~n4809;
  assign n5164 = ~n6607 & ~n6621;
  assign n5110 = ~n5109 & ~n5108;
  assign n6150 = ~n6093 | ~n6092;
  assign n5163 = ~n6540 | ~n5162;
  assign n5158 = ~n6471 | ~n6457;
  assign n5152 = ~n5151 | ~n6280;
  assign n4941 = ~n4940 | ~n4939;
  assign n6632 = ~n4921 | ~n4920;
  assign n7496 = ~n7667;
  assign n4694 = ~n4693 | ~n4692;
  assign n4566 = ~n5640;
  assign n5171 = ~n6791 | ~n6663;
  assign n6134 = ~n7747 & ~n6123;
  assign n5155 = ~n6439 | ~n6470;
  assign n4691 = ~n4690 & ~n4689;
  assign n7166 = ~n6928 & ~n5065;
  assign n7747 = ~n6122 | ~REG3_REG_28__SCAN_IN;
  assign n7667 = ~n7743 | ~n6779;
  assign n6713 = ~n6654 | ~n6792;
  assign n7201 = ~n6022 | ~n5994;
  assign n6290 = ~n6422;
  assign n7336 = ~n7560;
  assign n5153 = ~n6467 | ~n6436;
  assign n5169 = ~n6928 | ~n6700;
  assign n7057 = ~n6407 | ~n6539;
  assign n5145 = ~n6341 | ~n6163;
  assign n5123 = ~n5120 & ~n5656;
  assign n6471 = ~n6407;
  assign n4671 = ~n4669 & ~n4668;
  assign n4619 = ~n4616 | ~n4615;
  assign n6092 = ~n5907 | ~n5906;
  assign n7138 = ~n5879 | ~n5135;
  assign n6441 = ~n6543 | ~n6470;
  assign n7120 = ~n6832 | ~n6663;
  assign n7793 = ~n7700;
  assign n4667 = ~n4666 & ~n4665;
  assign n5137 = ~n5879 | ~n6016;
  assign n6439 = ~n6543;
  assign n6607 = ~n6706;
  assign n4646 = ~n4644 | ~n4643;
  assign n4642 = ~n4641 | ~n4640;
  assign n7521 = ~n7794;
  assign n4760 = ~n4759 & ~n4758;
  assign n5142 = ~n6261 | ~n6109;
  assign n7007 = ~n5991 | ~n5841;
  assign n4998 = ~n4996 & ~n4995;
  assign n4764 = ~n4762 & ~n4761;
  assign n5014 = ~n5013 & ~n5012;
  assign n5126 = ~n5819 | ~n5759;
  assign n4994 = ~n4993 & ~n4992;
  assign n7008 = ~n5819 & ~n5789;
  assign n4742 = ~n4739 | ~n4738;
  assign n7698 = ~n7533;
  assign n7252 = ~n7743 & ~REG2_REG_21__SCAN_IN;
  assign n7823 = ~n7537 & ~n7536;
  assign n4788 = ~n4787 & ~n4786;
  assign n5019 = ~n5017 & ~n5016;
  assign n4737 = ~n4736 | ~n4735;
  assign n7087 = ~n7117 | ~n7178;
  assign n7121 = ~n6716 & ~n7072;
  assign n5151 = ~n6467;
  assign n5149 = ~n6422 | ~n6335;
  assign n4709 = ~n4708 & ~n4707;
  assign n5156 = ~n6543 | ~n6382;
  assign n5118 = ~n7743 & ~REG2_REG_22__SCAN_IN;
  assign n7283 = ~n7282 | ~n7305;
  assign n5208 = ~n7596 & ~n6123;
  assign n4713 = ~n4711 & ~n4710;
  assign n5876 = ~n5811 & ~n5816;
  assign n7829 = ~n7505 & ~n7536;
  assign n6540 = ~n6627;
  assign n7072 = ~n7267 & ~n6722;
  assign n5139 = ~n6196 | ~n6068;
  assign n5894 = ~n5892 | ~n5891;
  assign n6341 = ~n6224;
  assign n7010 = ~n6162 | ~n6109;
  assign n6543 = ~n4851 | ~n4850;
  assign n7140 = ~n5965 | ~n5132;
  assign n6706 = ~n4897 | ~n4896;
  assign n6261 = ~n6162;
  assign n6944 = ~n7414 | ~n6943;
  assign n7628 = ~n7392;
  assign n6974 = ~n7832 & ~n7740;
  assign n5136 = ~n6063 | ~n5135;
  assign n7532 = ~n7788;
  assign n6819 = ~n7832 & ~n7636;
  assign n5906 = ~n5904 | ~n5903;
  assign n6467 = ~n4827 | ~n4826;
  assign n7143 = ~n6063 | ~n6016;
  assign n7177 = ~n5662 & ~n5658;
  assign n7123 = ~n7081 | ~n7079;
  assign n5811 = ~n5940 | ~n5759;
  assign n7013 = ~n5927 & ~n5759;
  assign n4996 = ~n6915 & ~n5015;
  assign n5078 = ~n7085;
  assign n6740 = ~n7267 & ~n6731;
  assign n5221 = ~n5220 | ~n5219;
  assign n5068 = ~n7082;
  assign n5233 = n5223 & n5222;
  assign n7084 = ~n7414 | ~n6964;
  assign n7196 = ~n5871 | ~n5816;
  assign n6928 = ~n4934 | ~n4933;
  assign n5187 = ~n5186 | ~n6904;
  assign n5226 = ~n5225 | ~n5224;
  assign n7808 = ~n7813;
  assign n6407 = ~n4516 | ~n4515;
  assign n5182 = ~n6889 | ~n5181;
  assign n5246 = ~n5245 | ~n5244;
  assign n7073 = ~n6915 | ~n6792;
  assign n5238 = ~n5228 | ~n5227;
  assign n4850 = ~n4849 & ~n4848;
  assign n7178 = ~n6937 | ~n6943;
  assign n5532 = n4501 & n4500;
  assign n7085 = ~n7268 & ~n6904;
  assign n7414 = ~n6937;
  assign n7620 = ~n7383;
  assign n7462 = ~n7452 | ~n7451;
  assign n5269 = ~n5263 & ~n5262;
  assign n7081 = ~n7268 | ~n6904;
  assign n7504 = ~n5430 & ~n5429;
  assign n7527 = ~n5104 | ~n5103;
  assign n4800 = ~n4799 & ~n4798;
  assign n7082 = ~n7411 & ~n5180;
  assign n5940 = ~n5938 & ~n5937;
  assign n7079 = ~n7411 | ~n5180;
  assign n6889 = ~n7411 | ~n7273;
  assign n5327 = ~n5326 & ~n5325;
  assign n6162 = ~n4753 & ~n4752;
  assign n7392 = n5507 & n5511;
  assign n6196 = ~n4728 | ~n4727;
  assign n5994 = ~n5132;
  assign n6937 = ~n5088 | ~n5087;
  assign n5009 = ~n5004 | ~n5003;
  assign n7397 = ~n7631 | ~ADDR_REG_17__SCAN_IN;
  assign n7411 = ~n5031 | ~n5030;
  assign n6199 = ~n6109;
  assign n4683 = ~n4678 | ~n4677;
  assign n4895 = ~n4892 | ~n4891;
  assign n4728 = ~n4722 & ~n4721;
  assign n4932 = ~n4929 | ~n4928;
  assign n5892 = ~n5902 | ~n5890;
  assign n4954 = ~n4951 | ~n4950;
  assign n4659 = ~n4651 | ~n4650;
  assign n7632 = ~n7631 | ~ADDR_REG_19__SCAN_IN;
  assign n5904 = ~n5902 | ~n5901;
  assign n7268 = ~n5077 | ~n5076;
  assign n4753 = ~n4747 | ~n4746;
  assign n4799 = ~n4796 | ~n4795;
  assign n4777 = ~n4773 | ~n4772;
  assign n4703 = ~n4698 | ~n4697;
  assign n6731 = ~n6722;
  assign n6068 = ~n6029;
  assign n6663 = ~n6924;
  assign n4776 = ~n4775 | ~n4774;
  assign n6621 = ~n6562;
  assign n4982 = ~n4981 | ~n4980;
  assign n4888 = ~n4526 & ~n5388;
  assign n5262 = ~n6123 & ~n7520;
  assign n5326 = ~n5323 | ~n5322;
  assign n5280 = ~n5278 | ~n5277;
  assign n4825 = ~n4822 | ~n4821;
  assign n4556 = ~n4550 & ~n4549;
  assign n6436 = ~n6280;
  assign n5104 = ~n5098 & ~n5097;
  assign n4501 = ~n4496 | ~n4526;
  assign n6382 = ~n6470;
  assign n5305 = ~n5303 | ~n5302;
  assign n4514 = ~n4509 | ~n4508;
  assign n4575 = ~n4569 & ~n4568;
  assign n5937 = ~n5124;
  assign n4849 = ~n4846 | ~n4845;
  assign n4632 = ~n4626 & ~n4625;
  assign n4898 = ~n4526 & ~n4517;
  assign n4536 = ~n4533 | ~n4532;
  assign n5207 = ~n5206 | ~n5205;
  assign n4532 = ~n5436 | ~REG0_REG_14__SCAN_IN;
  assign n4929 = ~n5321 | ~REG1_REG_16__SCAN_IN;
  assign n4574 = ~n4573 & ~n4572;
  assign n4891 = ~n5436 | ~REG0_REG_15__SCAN_IN;
  assign n7506 = ~n7657;
  assign n4508 = ~n5436 | ~REG0_REG_13__SCAN_IN;
  assign n4892 = ~n5321 | ~REG1_REG_15__SCAN_IN;
  assign n6029 = ~n4734 & ~n4733;
  assign n5253 = ~n7359 | ~n7772;
  assign n4533 = ~n5321 | ~REG1_REG_14__SCAN_IN;
  assign n4752 = ~n4751 | ~n4750;
  assign n5087 = ~n5086 & ~n5085;
  assign n4845 = ~n5436 | ~REG0_REG_12__SCAN_IN;
  assign n6016 = ~n4706 | ~n4705;
  assign n5206 = ~n5204 & ~n5203;
  assign n4631 = ~n4630 & ~n4629;
  assign n4702 = ~n4701 | ~n4700;
  assign n4981 = ~n4979 & ~n4978;
  assign n4928 = ~n5436 | ~REG0_REG_16__SCAN_IN;
  assign n4727 = ~n4726 & ~n4725;
  assign n5115 = ~n5481 | ~n5469;
  assign n5277 = ~n5436 | ~REG0_REG_25__SCAN_IN;
  assign n5278 = ~n5321 | ~REG1_REG_25__SCAN_IN;
  assign n5077 = ~n5071 & ~n5070;
  assign n4951 = ~n5321 | ~REG1_REG_17__SCAN_IN;
  assign n5031 = ~n5025 & ~n5024;
  assign n4775 = ~n5436 | ~REG0_REG_9__SCAN_IN;
  assign n4821 = ~n5436 | ~REG0_REG_11__SCAN_IN;
  assign n7559 = ~n7325;
  assign n5097 = ~n6123 & ~n7354;
  assign n4658 = ~n4657 | ~n4656;
  assign n4651 = ~n5321 | ~REG1_REG_4__SCAN_IN;
  assign n4555 = ~n4554 & ~n4553;
  assign n5901 = ~n5780 & ~n5779;
  assign n5003 = ~n5436 | ~REG0_REG_19__SCAN_IN;
  assign n5302 = ~n5436 | ~REG0_REG_26__SCAN_IN;
  assign n4950 = ~n5436 | ~REG0_REG_17__SCAN_IN;
  assign n5004 = ~n5321 | ~REG1_REG_19__SCAN_IN;
  assign n4682 = ~n4681 | ~n4680;
  assign n5303 = ~n5321 | ~REG1_REG_26__SCAN_IN;
  assign n7726 = ~n7748;
  assign n6109 = ~n4757 | ~n4756;
  assign n5400 = ~n5399;
  assign n4657 = ~n5320 | ~n4655;
  assign n4553 = ~n6125 & ~n4552;
  assign n4851 = ~n6528 | ~n5320;
  assign n5481 = ~n5471;
  assign n4549 = ~n6127 & ~n4548;
  assign n4629 = ~n6127 & ~n4628;
  assign n4630 = ~n6125 & ~n4627;
  assign n5470 = ~n5468 | ~n5467;
  assign n7699 = ~n7573;
  assign n7308 = ~n7522;
  assign n5028 = ~n6127 & ~n5027;
  assign n5261 = n5200 & REG3_REG_23__SCAN_IN;
  assign n5267 = ~n6125 & ~n5264;
  assign n5266 = ~n6127 & ~n5265;
  assign n7538 = ~n7500;
  assign n5024 = ~n6125 & ~n5023;
  assign n5102 = ~n6125 & ~n5099;
  assign n7273 = ~n5180;
  assign n4956 = ~n6919 | ~n5320;
  assign n5101 = ~n6127 & ~n5100;
  assign n5070 = ~n6125 & ~n5069;
  assign n5074 = ~n6127 & ~n5073;
  assign n6964 = ~n6943;
  assign n5116 = ~n5468 | ~n5114;
  assign n5086 = ~n6125 & ~n5083;
  assign n5085 = ~n6127 & ~n5084;
  assign n5081 = ~n6123 & ~n6959;
  assign n5467 = ~n5466 & ~n5465;
  assign n4625 = ~n6123 & ~REG3_REG_3__SCAN_IN;
  assign n4983 = ~n6831 & ~n6123;
  assign n4496 = ~n4454 | ~n4886;
  assign n5503 = ~n5502 | ~n5694;
  assign n7668 = ~n7746;
  assign n5114 = ~n5466;
  assign n5200 = n5096 & REG3_REG_22__SCAN_IN;
  assign n5466 = ~n5113 | ~n5112;
  assign n5694 = ~REG1_REG_6__SCAN_IN | ~n5692;
  assign n4491 = ~n5387 & ~D_REG_1__SCAN_IN;
  assign n5015 = ~n7777;
  assign n5096 = n5080 & REG3_REG_21__SCAN_IN;
  assign n7234 = ~n5388 & ~n5402;
  assign n5080 = n5072 & REG3_REG_20__SCAN_IN;
  assign n5113 = ~n5388;
  assign n5502 = ~n5704 | ~n5501;
  assign n7661 = ~n5472;
  assign n5521 = ~n5704 | ~n5520;
  assign n7779 = ~n5209;
  assign n4510 = n4439 ^ IR_REG_29__SCAN_IN;
  assign n7650 = ~n7725;
  assign n4886 = ~n4453 | ~n7725;
  assign n5388 = ~n4584 | ~n5395;
  assign n5501 = ~n5500 | ~n5711;
  assign n7757 = ~n7542;
  assign n5026 = ~n5005 | ~REG3_REG_18__SCAN_IN;
  assign n5396 = ~n5392 & ~n4490;
  assign n5711 = ~n5708 | ~n5709;
  assign n5465 = ~n7678 & ~n7176;
  assign n5112 = ~n5095 | ~n7224;
  assign n6500 = ~REG1_REG_13__SCAN_IN | ~n6508;
  assign n5005 = ~n4974 & ~n6914;
  assign n7647 = ~n7720;
  assign n5474 = ~n5401;
  assign n4430 = ~n4438 | ~IR_REG_31__SCAN_IN;
  assign n4490 = ~n4483;
  assign n5272 = ~n7775;
  assign n4492 = ~n5390;
  assign n4974 = ~n4949 | ~REG3_REG_16__SCAN_IN;
  assign n7775 = ~n5657 | ~n4543;
  assign n4486 = ~n5390 | ~n4485;
  assign n5095 = ~n5105;
  assign n6779 = ~n5657 & ~n7485;
  assign n4451 = ~n7224;
  assign n6083 = ~REG1_REG_9__SCAN_IN | ~n6091;
  assign n5105 = ~n7176 | ~n7238;
  assign n5518 = ~n5600 | ~n5517;
  assign n4949 = ~n4927 & ~n6624;
  assign n4528 = ~n7226;
  assign n6093 = ~REG2_REG_9__SCAN_IN | ~n6091;
  assign n5499 = ~n5600 | ~n5498;
  assign n6357 = n4867 ^ n4866;
  assign n4527 = ~n7238;
  assign n5517 = ~n5516 | ~n5737;
  assign n4868 = ~n4867 | ~n4866;
  assign n7224 = ~n4539 | ~n7485;
  assign n7226 = ~n4539 | ~n7636;
  assign n4927 = ~n4890 | ~REG3_REG_14__SCAN_IN;
  assign n6091 = n4782 ^ n4781;
  assign n4961 = ~n4959 | ~IR_REG_31__SCAN_IN;
  assign n6316 = ~REG2_REG_11__SCAN_IN | ~n6314;
  assign n4539 = ~n7115;
  assign n4890 = ~n4505 & ~n6355;
  assign n6306 = ~REG1_REG_11__SCAN_IN | ~n6314;
  assign n5902 = n4779 ^ n4778;
  assign n4959 = ~n4958 | ~n4957;
  assign n7485 = ~n7636;
  assign n4505 = ~n4844 | ~REG3_REG_12__SCAN_IN;
  assign n5500 = ~REG1_REG_5__SCAN_IN | ~n5722;
  assign n7387 = n4958 ^ n4957;
  assign n4855 = ~n4854 | ~n4853;
  assign n5519 = ~REG2_REG_5__SCAN_IN | ~n5722;
  assign n4780 = ~n4779 | ~n4778;
  assign n5779 = ~REG2_REG_7__SCAN_IN & ~n5767;
  assign n5778 = REG2_REG_7__SCAN_IN & n5767;
  assign n4489 = ~n4482 & ~n4481;
  assign n5515 = ~n5514 | ~n5559;
  assign n5769 = ~REG1_REG_7__SCAN_IN | ~n5767;
  assign n4989 = ~n4988 | ~IR_REG_31__SCAN_IN;
  assign n6151 = n4806 ^ IR_REG_10__SCAN_IN;
  assign n4936 = ~n4987 | ~n4935;
  assign n6680 = n4523 ^ n4522;
  assign n4988 = ~n4987 | ~n4986;
  assign n4755 = ~n4754 | ~n4802;
  assign n5514 = ~REG2_REG_2__SCAN_IN | ~n5571;
  assign n6062 = ~n4720 | ~n4749;
  assign n4685 = ~n4684 & ~IR_REG_4__SCAN_IN;
  assign n5557 = ~n5513 | ~n5626;
  assign n4794 = n4771 & REG3_REG_9__SCAN_IN;
  assign n5562 = ~n5494 | ~n5635;
  assign n5495 = ~REG1_REG_2__SCAN_IN | ~n5571;
  assign n4636 = ~n4634 | ~IR_REG_31__SCAN_IN;
  assign n4731 = ~n4805 | ~IR_REG_31__SCAN_IN;
  assign n4771 = ~n4749 & ~n4748;
  assign n5626 = ~n5624 | ~n5623;
  assign n4699 = ~n6021;
  assign n5635 = ~n5633 | ~n5632;
  assign n5856 = ~n4654 | ~n4679;
  assign n4986 = ~n4985 & ~IR_REG_17__SCAN_IN;
  assign n4388 = ~n4384 & ~n4383;
  assign n4718 = ~n4679 & ~n4502;
  assign n5632 = ~n4607 & ~n4579;
  assign n7395 = ~STATE_REG_SCAN_IN & ~n6914;
  assign n4504 = ~n5510 & ~n4503;
  assign n5623 = ~n4607 & ~n4567;
  assign n4804 = ~n4803 | ~n4802;
  assign n4442 = ~IR_REG_29__SCAN_IN;
  assign n4866 = ~IR_REG_12__SCAN_IN;
  assign n6355 = ~REG3_REG_13__SCAN_IN;
  assign n4436 = ~IR_REG_28__SCAN_IN;
  assign n5381 = ~IR_REG_30__SCAN_IN;
  assign n4435 = ~IR_REG_27__SCAN_IN;
  assign n4802 = ~IR_REG_7__SCAN_IN;
  assign n4512 = ~REG2_REG_13__SCAN_IN;
  assign n5301 = ~REG3_REG_26__SCAN_IN;
  assign n4847 = ~REG2_REG_12__SCAN_IN;
  assign n4679 = ~REG3_REG_3__SCAN_IN | ~REG3_REG_4__SCAN_IN;
  assign n4778 = ~IR_REG_8__SCAN_IN;
  assign n4426 = ~IR_REG_26__SCAN_IN;
  assign n4935 = ~IR_REG_15__SCAN_IN;
  assign n4853 = ~IR_REG_11__SCAN_IN;
  assign n4960 = ~IR_REG_17__SCAN_IN;
  assign n6914 = ~REG3_REG_17__SCAN_IN;
  assign n4914 = ~DATAI_15_;
  assign n6624 = ~REG3_REG_15__SCAN_IN;
  assign n4803 = ~IR_REG_8__SCAN_IN & ~IR_REG_9__SCAN_IN;
  assign n4893 = ~REG2_REG_15__SCAN_IN;
  assign n5032 = ~REG3_REG_19__SCAN_IN;
  assign n4394 = ~IR_REG_21__SCAN_IN;
  assign n4912 = ~IR_REG_31__SCAN_IN;
  assign n4389 = ~IR_REG_18__SCAN_IN;
  assign n4534 = ~REG2_REG_14__SCAN_IN;
  assign n4397 = ~IR_REG_24__SCAN_IN;
  assign n7754 = ~n7745 | ~n7744;
  assign n7615 = ~n7613 | ~n7767;
  assign n7612 = ~n7613 | ~n7763;
  assign n7604 = ~n7595 | ~n7594;
  assign n7689 = ~n7687 | ~n7763;
  assign n7686 = ~n7687 | ~n7767;
  assign n7662 = ~n7679 & ~n7661;
  assign n7675 = ~n7679 & ~n7667;
  assign n7682 = ~n7679 & ~n7678;
  assign n5339 = ~n5318 & ~n7813;
  assign n7583 = ~n7605 & ~n7661;
  assign n7711 = ~n7695 | ~n7808;
  assign n7445 = ~n7444 & ~n7443;
  assign n7570 = ~n7557 | ~n7808;
  assign n7535 = ~n7531 & ~n7530;
  assign n7315 = ~n7314 | ~n7313;
  assign n7557 = ~n4378 | ~n7556;
  assign n7531 = ~n7526 | ~n7525;
  assign n7343 = ~n7330 & ~n7329;
  assign n7493 = ~n7299 | ~n7298;
  assign n7526 = ~n7519 | ~n7553;
  assign n7298 = ~n7297 & ~n7296;
  assign n5299 = ~n5291 & ~n5290;
  assign n7297 = ~n7293 & ~n7303;
  assign n6953 = ~n6951 | ~n7767;
  assign n7491 = ~n7304 | ~n7303;
  assign n6950 = ~n6951 | ~n7763;
  assign n7293 = ~n7292 & ~n7291;
  assign n5199 = ~n5119 & ~n5118;
  assign n6908 = ~n6907 & ~n7246;
  assign n7244 = ~n7233 | ~n7232;
  assign n7663 = ~n7656 | ~n7655;
  assign n7656 = ~n7648 | ~n7647;
  assign n6948 = ~n6947 & ~n6946;
  assign n7233 = ~n7231 | ~n7230;
  assign n5119 = ~n6877 & ~n7832;
  assign n7231 = ~n7116 | ~n7115;
  assign n7254 = ~n6891 ^ n7001;
  assign n7408 = ~n7404 & ~n7403;
  assign n6826 = ~n6825 | ~n6974;
  assign n7646 = ~n7712 & ~n7645;
  assign n5111 = ~n5094 | ~n7647;
  assign n7590 = ~n7589 | ~n7647;
  assign n5197 = ~n6879 | ~n6974;
  assign n7114 = ~n7113 | ~n7112;
  assign n7435 = ~n7434 & ~n7720;
  assign n5094 = ~n5091 | ~n6931;
  assign n6880 = ~n6879 | ~n6878;
  assign n6890 = ~n6888 | ~n6887;
  assign n6856 = ~n6854 & ~n6853;
  assign n7342 = ~n7335 & ~n7720;
  assign n6733 = ~n6775 & ~n7678;
  assign n6853 = ~n7832 & ~n6852;
  assign n6757 = ~n6816 & ~n6820;
  assign n6785 = ~n6797 | ~n6779;
  assign n6818 = ~n6816 & ~n7832;
  assign n7433 = ~n7584 & ~n7432;
  assign n7258 = ~n5002 | ~n5001;
  assign n6902 = ~n6901 | ~n6900;
  assign n6816 = ~n6753 | ~n6752;
  assign n6807 = ~n6806 & ~n7678;
  assign n7301 = ~n7300 | ~n7647;
  assign n6666 = ~n6661 & ~n6845;
  assign n5185 = ~n6778 | ~n5176;
  assign n6644 = ~n6641 | ~n6640;
  assign n6641 = ~n6616 & ~n6615;
  assign n6846 = ~n6844 & ~n7661;
  assign n7096 = ~n7643 | ~n7095;
  assign n6494 = ~n6491 | ~n6490;
  assign n6845 = ~n6660 | ~n6659;
  assign n6613 = ~n6612 | ~n5472;
  assign n6602 = ~n6612 | ~n6779;
  assign n6583 = ~n7832 & ~n6591;
  assign n6660 = ~n6658 & ~n6657;
  assign n6638 = ~n6637 & ~n7678;
  assign n6462 = ~n7767 | ~n6464;
  assign n6486 = ~n6411 & ~n6410;
  assign n6465 = ~n7763 | ~n6464;
  assign n6464 = ~n6516 | ~n6461;
  assign n6789 = ~n5066 & ~n7071;
  assign n6519 = ~n7832 & ~n6516;
  assign n6415 = ~n6489 | ~n7496;
  assign n6589 = ~n6586 & ~n7678;
  assign n7090 = ~n7080 | ~n7285;
  assign n6582 = ~n6586 & ~n7667;
  assign n6391 = ~n7763 | ~n6390;
  assign n6516 = ~n6456 & ~n6455;
  assign n6388 = ~n7767 | ~n6390;
  assign n7078 = ~n7070 | ~n7121;
  assign n6390 = ~n6530 | ~n6387;
  assign n7070 = ~n7069 & ~n7068;
  assign n6530 = ~n6381 & ~n6380;
  assign n6605 = ~n5064 | ~n7125;
  assign n6453 = ~n6524 | ~n5472;
  assign n6327 = ~n7767 | ~n6329;
  assign n6303 = ~n7743 | ~n6301;
  assign n7543 = ~n7824 | ~n7542;
  assign n4885 = ~n4882 & ~n4881;
  assign n7639 = ~n7635 & ~n7634;
  assign n6330 = ~n7763 | ~n6329;
  assign n6571 = ~n6570 | ~n6569;
  assign n6478 = ~n6553 & ~n7813;
  assign n4882 = ~n6476 & ~n4865;
  assign n7508 = ~n7831 | ~n7542;
  assign n7634 = ~n7633 | ~n7632;
  assign n6428 = ~n6427 | ~n7808;
  assign n6246 = ~n7763 | ~n6245;
  assign n6235 = ~n6234 | ~n7743;
  assign n7633 = ~n7630 & ~n7629;
  assign n7680 = ~n7671 | ~n7670;
  assign n6243 = ~n7767 | ~n6245;
  assign n6405 = ~n5061 | ~n5060;
  assign n7599 = ~n7606 & ~n7750;
  assign n7635 = ~n7621 & ~n7620;
  assign n6442 = ~n7056 | ~n6440;
  assign n6386 = ~n6527 | ~n7312;
  assign n7402 = ~n7400 & ~n7399;
  assign n6286 = ~n6285 | ~n6284;
  assign n7061 = ~n7056 & ~n7158;
  assign n7630 = ~n7628 & ~n7627;
  assign n6535 = ~n6527 | ~n6779;
  assign n6296 = ~n6295 | ~n5472;
  assign n7598 = ~n7597 | ~n7657;
  assign n6189 = ~n7832 & ~n6188;
  assign n6285 = ~n6295 | ~n6779;
  assign n7670 = ~n7669 | ~n7780;
  assign n7478 = ~n7597 | ~n7442;
  assign n6260 = ~n6258 | ~n7743;
  assign n7228 = ~n7227 | ~n7226;
  assign n5058 = ~n6288 & ~n7133;
  assign n6258 = ~n6257 | ~n6256;
  assign n7489 = ~n7486 | ~n7485;
  assign n7626 = ~n7624 | ~n7623;
  assign n4819 = ~n4814 | ~n6333;
  assign n6177 = ~n7767 | ~n6179;
  assign n7371 = ~n7328 | ~n7441;
  assign n7229 = ~n7225 | ~n7224;
  assign n6339 = ~n6334 & ~n7813;
  assign n6323 = ~n6322 & ~n7678;
  assign n6180 = ~n7763 | ~n6179;
  assign n7619 = ~n7617 | ~n7616;
  assign n7328 = ~n7326 | ~n7325;
  assign n6120 = ~n7763 | ~n6119;
  assign n7617 = ~n7468 | ~n7467;
  assign n6187 = ~n6184 | ~n6183;
  assign n6117 = ~n7767 | ~n6119;
  assign n7442 = ~n7441 | ~n7699;
  assign n6230 = ~n6223 | ~n7647;
  assign n7486 = ~n7310 & ~n7327;
  assign n6212 = ~n6211 | ~n6210;
  assign n7310 = ~n7307 | ~n7542;
  assign n6240 = n6237 & n7312;
  assign n7384 = ~n7383 | ~n7464;
  assign n6232 = n6237 & n5472;
  assign n6255 = ~n6252 | ~n6251;
  assign n7307 = ~n7309 | ~n7308;
  assign n6978 = ~n6976 & ~n7750;
  assign n6222 = ~n5054 & ~n7011;
  assign n7385 = ~n7382 & ~n7381;
  assign n6876 = ~n5193 & ~n7306;
  assign n7249 = ~n7246 | ~n7485;
  assign n6822 = ~n6820 | ~n6819;
  assign n6175 = ~n6185 & ~n7755;
  assign n5193 = ~n5191 | ~n7542;
  assign n6820 = ~n6756 & ~n6905;
  assign n5191 = ~n5192 | ~n6964;
  assign n7214 = ~n7586 & ~n7212;
  assign n6104 = ~n6102 | ~n7647;
  assign n6871 = ~REG2_REG_16__SCAN_IN & ~n6872;
  assign n7379 = ~REG2_REG_16__SCAN_IN | ~n6872;
  assign n7388 = ~REG1_REG_16__SCAN_IN | ~n6862;
  assign n6861 = ~REG1_REG_16__SCAN_IN & ~n6862;
  assign n6756 = ~n6755 | ~n7542;
  assign n6045 = ~n6044 | ~n6043;
  assign n6784 = ~n6808 | ~n7485;
  assign n5053 = ~n6101 | ~n7010;
  assign n7212 = ~n7585 & ~n7211;
  assign n6850 = ~n6849 & ~n7636;
  assign n6677 = ~n7383 | ~n6869;
  assign n6685 = ~n6859 | ~n7392;
  assign n6101 = ~n5052 & ~n5051;
  assign n6808 = ~n6783 & ~n6782;
  assign n6755 = ~n6754 | ~n7273;
  assign n6765 = ~n6754 | ~n7542;
  assign n7113 = ~n7052 | ~n7108;
  assign n5982 = ~n5969 | ~n5968;
  assign n6783 = ~n6781 | ~n7542;
  assign n6686 = ~n6684 & ~n6683;
  assign n6601 = ~n6639 | ~n7485;
  assign n6514 = ~n6513 | ~n6673;
  assign n6678 = ~n6676 & ~n6675;
  assign n5918 = ~n5915 | ~n5914;
  assign n5052 = ~n6037 & ~n7036;
  assign n6764 = ~n6782 & ~n6731;
  assign n6037 = ~n5049 | ~n7138;
  assign n6664 = ~n7542 | ~n6780;
  assign n6781 = ~n6792 | ~n6780;
  assign n7032 = ~n7031 & ~n7572;
  assign n5912 = ~n5875 | ~n5874;
  assign n6665 = ~n6663 & ~n6662;
  assign n6599 = ~n7757 & ~n6662;
  assign n5049 = ~n5961 | ~n7143;
  assign n6501 = ~REG1_REG_14__SCAN_IN & ~n6502;
  assign n6511 = ~REG2_REG_14__SCAN_IN & ~n6512;
  assign n5961 = ~n5048 | ~n7201;
  assign n6362 = ~n6499 | ~n7392;
  assign n5048 = ~n5869 | ~n7140;
  assign n6354 = ~n6352 & ~n6351;
  assign n6310 = ~n6309 | ~n6358;
  assign n6363 = ~n6361 & ~n6360;
  assign n5869 = ~n5047 | ~n7007;
  assign n6397 = ~n6396 | ~n6395;
  assign n5047 = ~n5046 | ~n7196;
  assign n6307 = ~REG1_REG_12__SCAN_IN & ~n6308;
  assign n7815 = ~n7814 & ~n7813;
  assign n7810 = ~n7818;
  assign n5814 = ~n5045 | ~n7193;
  assign n7693 = ~n7692 | ~n7691;
  assign n6475 = ~n6474 | ~n6552;
  assign n7103 = ~n7102 | ~n7713;
  assign n7213 = n7643 & n7102;
  assign n7812 = ~n7786 | ~n7785;
  assign n6423 = ~n4842 & ~n4841;
  assign n7060 = ~n7059 | ~n7162;
  assign n5297 = ~n7550 | ~n7551;
  assign n5755 = ~n5044 | ~n7192;
  assign n7739 = ~n7718 & ~n7717;
  assign n7125 = ~n5063 & ~n5062;
  assign n6695 = ~n4944 & ~n4945;
  assign n7162 = ~n7058 | ~n7057;
  assign n6551 = ~n4884 & ~n4883;
  assign n6449 = ~n7041;
  assign n4595 = ~n4592 & ~n5639;
  assign n5316 = ~n5313;
  assign n7062 = ~n7130;
  assign n7718 = ~n7716;
  assign n7550 = ~n5294 | ~n5289;
  assign n5997 = n4695 ^ n4694;
  assign n5216 = ~n7791 | ~n7777;
  assign n7119 = n7077 & n7076;
  assign n7585 = ~n7053 | ~n7431;
  assign n7089 = ~n7288 & ~n7088;
  assign n7066 = ~n7065 | ~n7064;
  assign n7645 = ~n7644;
  assign n6110 = ~n6030 | ~n6029;
  assign n4594 = ~n4593 & ~n5640;
  assign n7736 = ~n7778 & ~n7780;
  assign n6152 = ~REG2_REG_10__SCAN_IN | ~n6095;
  assign n7259 = ~n5018 | ~n5019;
  assign n5928 = ~n5666 | ~n5042;
  assign n4673 = ~n4670;
  assign n7432 = ~n7431;
  assign n7058 = ~n5158 | ~n6440;
  assign n6940 = ~n6939 | ~n6938;
  assign n7041 = ~n5158 | ~n7057;
  assign n7130 = ~n5164 & ~n5161;
  assign n7133 = ~n5151 & ~n6436;
  assign n7053 = ~n7574 | ~n7699;
  assign n6658 = ~n6649 & ~n7424;
  assign n5213 = ~n7696 & ~n5209;
  assign n4695 = n4691 ^ n7775;
  assign n6984 = ~n7138 | ~n7143;
  assign n5161 = ~n6540 & ~n6395;
  assign n7059 = ~n6540 | ~n6395;
  assign n6456 = ~n6439 & ~n7424;
  assign n4670 = n4667 ^ n5272;
  assign n7064 = ~n6607 | ~n6621;
  assign n4672 = ~n4671;
  assign n6488 = ~n6394 | ~n6393;
  assign n5177 = ~n6713 & ~n6742;
  assign n6440 = ~n6439 | ~n6382;
  assign n7644 = ~n7696 | ~n7657;
  assign n6113 = ~n6999 | ~n7010;
  assign n7158 = ~n7057 | ~n6441;
  assign n5666 = ~n7038 | ~n7177;
  assign n5166 = ~n6607 | ~n6562;
  assign n6030 = ~n5971 & ~n6016;
  assign n6012 = ~n4709 ^ n7775;
  assign n7132 = ~n6290 & ~n6335;
  assign n4940 = ~n6928 | ~n7779;
  assign n7071 = ~n6832 & ~n6663;
  assign n7074 = ~n7015;
  assign n5133 = ~n6022 | ~n5132;
  assign n7323 = ~n7336 & ~n7522;
  assign n7055 = ~n7533 | ~n7559;
  assign n4968 = ~n6832 | ~n7777;
  assign n7174 = ~n7331 & ~n7287;
  assign n7036 = ~n7136 | ~n7144;
  assign n4965 = ~n6832 | ~n7779;
  assign n7149 = ~n6422 & ~n5147;
  assign n7093 = ~n7579 | ~n7573;
  assign n4693 = ~n6022 | ~n7777;
  assign n5534 = ~n4589;
  assign n4860 = ~n6543 | ~n7779;
  assign n6788 = ~n6713 | ~n6712;
  assign n5309 = ~n7579 | ~n7779;
  assign n5288 = ~n7533 | ~n7777;
  assign n4863 = ~n6543 | ~n7777;
  assign n4810 = ~n6422 | ~n7779;
  assign n7124 = ~n6928 | ~n5065;
  assign n7011 = ~n6341 & ~n6264;
  assign n5312 = ~n7579 | ~n7777;
  assign n5172 = ~n6832 | ~n6924;
  assign n4874 = ~n6407 | ~n7779;
  assign n5285 = ~n7533 | ~n7779;
  assign n6999 = ~n6261 | ~n6199;
  assign n6742 = ~n6834 & ~n6722;
  assign n4618 = n4614 ^ n7775;
  assign n4877 = ~n6407 | ~n7777;
  assign n6559 = ~n7521 & ~n6548;
  assign n4838 = ~n6467 | ~n7777;
  assign n4542 = ~n6627 | ~n7779;
  assign n4835 = ~n6467 | ~n7779;
  assign n5971 = ~n5876 | ~n5994;
  assign n7285 = ~n7123 & ~n7087;
  assign n4790 = ~n6341 | ~n7777;
  assign n7038 = ~n7185 & ~n7180;
  assign n4921 = ~n6706 | ~n7777;
  assign n7159 = ~n6467 & ~n6280;
  assign n5328 = ~n7795 | ~n5320;
  assign n4813 = ~n6422 | ~n7777;
  assign n5129 = ~n5991 | ~n5816;
  assign n7752 = ~n7747 & ~n7746;
  assign n7299 = ~n7533 | ~n7503;
  assign n4918 = ~n6706 | ~n7779;
  assign n5275 = ~n7560 | ~n7777;
  assign n4614 = ~n4613 | ~n4612;
  assign n5131 = ~n5965 | ~n5994;
  assign n5255 = ~n5254 | ~n5253;
  assign n7144 = ~n5050 | ~n6068;
  assign n5258 = ~n5257 | ~n5256;
  assign n4690 = ~n5965 & ~n5209;
  assign n4666 = ~n5871 & ~n5209;
  assign n5640 = ~n4565 | ~n4564;
  assign n7296 = ~n7295 | ~n7294;
  assign n4669 = ~n5871 & ~n5015;
  assign n5271 = ~n7560 | ~n7779;
  assign n7024 = ~n5068 | ~n7079;
  assign n7148 = ~n6224 & ~n6163;
  assign n7086 = ~n7084 | ~n7083;
  assign n6817 = ~n7743 & ~REG2_REG_20__SCAN_IN;
  assign n7001 = ~n5078 | ~n7081;
  assign n7054 = ~n7560 | ~n7522;
  assign n5017 = ~n7267 & ~n5015;
  assign n5144 = ~n6224 | ~n6264;
  assign n6920 = ~n7794 | ~n6919;
  assign n6925 = ~n7700 | ~n6924;
  assign n4711 = ~n6063 & ~n5015;
  assign n4708 = ~n6063 & ~n5209;
  assign n7579 = ~n5307 | ~n5306;
  assign n7015 = ~n7267 | ~n6722;
  assign n4589 = ~n4583 | ~n4582;
  assign n4759 = ~n6162 & ~n5209;
  assign n5141 = ~n6162 | ~n6199;
  assign n4787 = ~n6224 & ~n5209;
  assign n4762 = ~n6162 & ~n5015;
  assign n4993 = ~n6915 & ~n5209;
  assign n4955 = ~n4954 & ~n4953;
  assign n6923 = ~n6915 & ~n7788;
  assign n5281 = ~n5280 & ~n5279;
  assign n5871 = ~n4659 & ~n4658;
  assign n7826 = ~n7832 | ~REG2_REG_31__SCAN_IN;
  assign n5965 = ~n4683 & ~n4682;
  assign n7833 = ~n7832 | ~REG2_REG_30__SCAN_IN;
  assign n5307 = ~n7705 | ~n5320;
  assign n7136 = ~n6196 | ~n6029;
  assign n6122 = n5319 & REG3_REG_27__SCAN_IN;
  assign n6712 = ~n6915 | ~n6833;
  assign n4896 = ~n4895 & ~n4894;
  assign n4515 = ~n4514 & ~n4513;
  assign n7665 = ~n7832 | ~n7664;
  assign n5306 = ~n5305 & ~n5304;
  assign n4736 = ~n6196 | ~n7779;
  assign n6520 = ~REG2_REG_13__SCAN_IN | ~n7832;
  assign n6887 = ~n6895 | ~n5180;
  assign n4826 = ~n4825 & ~n4824;
  assign n5250 = ~n5248 | ~n5247;
  assign n6716 = ~n6915 & ~n6792;
  assign n7117 = ~n7527 | ~n7305;
  assign n5257 = ~n7527 | ~n7777;
  assign n7287 = ~n7527 & ~n7305;
  assign n4933 = ~n4932 & ~n4931;
  assign n4739 = ~n6196 | ~n7777;
  assign n7560 = ~n5269 | ~n5268;
  assign n4537 = ~n4536 & ~n4535;
  assign n7474 = ~n7832 | ~n7473;
  assign n5121 = ~n5924;
  assign n7368 = ~n7832 | ~n7367;
  assign n5254 = ~n7527 | ~n7779;
  assign n5282 = ~n7558 | ~n5320;
  assign n5220 = ~n7411 | ~n7779;
  assign n5181 = ~n7268 | ~n7417;
  assign n4789 = ~n6163 | ~n7779;
  assign n4834 = ~n6436 | ~n7772;
  assign n4995 = ~n6833 & ~n5209;
  assign n4837 = ~n6436 | ~n7779;
  assign n5891 = ~REG1_REG_8__SCAN_IN | ~n5771;
  assign n4859 = ~n6382 | ~n7772;
  assign n5245 = ~n6937 | ~n7779;
  assign n4862 = ~n6382 | ~n7779;
  assign n4873 = ~n6457 | ~n7772;
  assign n5228 = ~n7268 | ~n7777;
  assign n4992 = ~n6833 & ~n5211;
  assign n7813 = ~n4888 | ~n4887;
  assign n4876 = ~n6457 | ~n7779;
  assign n5225 = ~n7268 | ~n7779;
  assign n4545 = ~n5162 & ~n5209;
  assign n4917 = ~n6621 | ~n7772;
  assign n4920 = ~n6621 | ~n7779;
  assign n4942 = ~n5065 & ~n5209;
  assign n7460 = ~n7637 | ~n7622;
  assign n7832 = ~n5117 & ~n7668;
  assign n6865 = ~n7637 | ~n7387;
  assign n4665 = ~n5841 & ~n5211;
  assign n4668 = ~n5841 & ~n5209;
  assign n5903 = ~REG2_REG_8__SCAN_IN | ~n5782;
  assign n4689 = ~n5994 & ~n5211;
  assign n4707 = ~n5135 & ~n5211;
  assign n5248 = ~n6937 | ~n7777;
  assign n4710 = ~n5135 & ~n5209;
  assign n4735 = ~n6068 | ~n7772;
  assign n4738 = ~n6068 | ~n7779;
  assign n4761 = ~n6199 & ~n5209;
  assign n4758 = ~n6199 & ~n5211;
  assign n4692 = ~n5132 | ~n7779;
  assign n6659 = ~n6924 | ~n7650;
  assign n6833 = ~n6792;
  assign n4509 = ~n5321 | ~REG1_REG_13__SCAN_IN;
  assign n4678 = ~n5321 | ~REG1_REG_5__SCAN_IN;
  assign n4822 = ~n5321 | ~REG1_REG_11__SCAN_IN;
  assign n4846 = ~n5321 | ~REG1_REG_12__SCAN_IN;
  assign n4796 = ~n5321 | ~REG1_REG_10__SCAN_IN;
  assign n6457 = ~n6539;
  assign n5323 = ~n5321 | ~REG1_REG_28__SCAN_IN;
  assign n4698 = ~n5321 | ~REG1_REG_6__SCAN_IN;
  assign n5065 = ~n6700;
  assign n4541 = ~n6395 | ~n7772;
  assign n4812 = ~n6335 | ~n7779;
  assign n4964 = ~n6924 | ~n7772;
  assign n4786 = ~n6264 & ~n5211;
  assign n4939 = ~n6700 | ~n7772;
  assign n4747 = ~n5321 | ~REG1_REG_8__SCAN_IN;
  assign n4772 = ~n5321 | ~REG1_REG_9__SCAN_IN;
  assign n7383 = ~n5529 & ~n5512;
  assign n4809 = ~n6335 | ~n7772;
  assign n4967 = ~n6924 | ~n7779;
  assign n4677 = ~n5436 | ~REG0_REG_5__SCAN_IN;
  assign n4795 = ~n5436 | ~REG0_REG_10__SCAN_IN;
  assign n5816 = ~n4664 | ~n4663;
  assign n5132 = ~n4688 | ~n4687;
  assign n4697 = ~n5436 | ~REG0_REG_6__SCAN_IN;
  assign n5529 = ~n5506 | ~n5505;
  assign n4746 = ~n5436 | ~REG0_REG_8__SCAN_IN;
  assign n5227 = ~n7417 | ~n7779;
  assign n5008 = ~n5007 | ~n5006;
  assign n4650 = ~n5436 | ~REG0_REG_4__SCAN_IN;
  assign n5244 = ~n6964 | ~n7772;
  assign n5224 = ~n7417 | ~n7772;
  assign n5268 = ~n5267 & ~n5266;
  assign n5076 = ~n5075 & ~n5074;
  assign n5103 = ~n5102 & ~n5101;
  assign n4526 = ~n5468 | ~n4495;
  assign n5247 = ~n6964 | ~n7779;
  assign n5088 = ~n5082 & ~n5081;
  assign n5030 = ~n5029 & ~n5028;
  assign n5321 = ~n6125;
  assign n4681 = ~n5320 | ~n6006;
  assign n4751 = ~n5320 | ~n6250;
  assign n4726 = ~n6125 & ~n4723;
  assign n4725 = ~n6127 & ~n4724;
  assign n4773 = ~n5320 | ~n6276;
  assign n4701 = ~n5320 | ~n4699;
  assign n5007 = ~n5320 | ~n6767;
  assign n5780 = ~n5778 & ~n5777;
  assign n4979 = ~n6125 & ~n4976;
  assign n4978 = ~n6127 & ~n4977;
  assign n7359 = ~n7305;
  assign n5203 = ~n6127 & ~n5202;
  assign n7722 = ~n7424;
  assign n4721 = ~n6123 & ~n6062;
  assign n5029 = ~n6123 & ~n7266;
  assign n5075 = ~n6123 & ~n7410;
  assign n6787 = ~n6831 & ~n7746;
  assign n4554 = ~n6123 & ~n4551;
  assign n5777 = ~n5521 | ~n5698;
  assign n6878 = ~n7755;
  assign n5698 = ~REG2_REG_6__SCAN_IN | ~n5696;
  assign n4494 = ~n5387 & ~D_REG_0__SCAN_IN;
  assign n4507 = ~n4510;
  assign n4488 = ~n4487 | ~n4486;
  assign n5520 = ~n5519 | ~n5716;
  assign n4493 = ~n5392 & ~n4492;
  assign n5716 = ~n5713 | ~n5714;
  assign n4487 = ~n4484 | ~B_REG_SCAN_IN;
  assign n5714 = ~n5518 | ~n5594;
  assign n6510 = ~REG2_REG_13__SCAN_IN | ~n6508;
  assign n7312 = ~n7678;
  assign n4484 = ~n4483 | ~n5390;
  assign n5402 = ~n5095 | ~n4451;
  assign n5709 = ~n5499 | ~n5590;
  assign n4403 = ~n4483 & ~n5390;
  assign n5590 = ~REG1_REG_4__SCAN_IN | ~n5589;
  assign n7678 = ~n4528 | ~n4527;
  assign n4540 = ~n5657;
  assign n4483 = n4400 ^ IR_REG_25__SCAN_IN;
  assign n5594 = ~REG2_REG_4__SCAN_IN | ~n5593;
  assign n5390 = ~n4402 ^ IR_REG_24__SCAN_IN;
  assign n7465 = ~REG2_REG_17__SCAN_IN | ~n7463;
  assign n4869 = ~n4868 | ~IR_REG_31__SCAN_IN;
  assign n7454 = ~REG1_REG_17__SCAN_IN | ~n7463;
  assign n4543 = ~n7238 | ~n7485;
  assign n5498 = ~n5497 | ~n5729;
  assign n7238 = n4408 ^ IR_REG_22__SCAN_IN;
  assign n7616 = ~n7622 | ~REG2_REG_18__SCAN_IN;
  assign n4782 = ~n4780 | ~IR_REG_31__SCAN_IN;
  assign n5737 = ~REG2_REG_3__SCAN_IN | ~n5735;
  assign n5729 = ~REG1_REG_3__SCAN_IN | ~n5727;
  assign n4867 = ~n4855 | ~IR_REG_31__SCAN_IN;
  assign n7624 = ~n7622 | ~REG1_REG_18__SCAN_IN;
  assign n4416 = ~n4415 | ~n4414;
  assign n5497 = ~n5726 | ~n5496;
  assign n5516 = ~n5726 | ~n5515;
  assign n6860 = ~REG1_REG_15__SCAN_IN | ~n6868;
  assign n6870 = ~REG2_REG_15__SCAN_IN | ~n6868;
  assign n4958 = ~n4936 | ~IR_REG_31__SCAN_IN;
  assign n5496 = ~n5495 | ~n5564;
  assign n4844 = n4820 & REG3_REG_11__SCAN_IN;
  assign n4779 = ~n4755 | ~IR_REG_31__SCAN_IN;
  assign n4830 = ~n4852 | ~IR_REG_31__SCAN_IN;
  assign n4913 = ~n4987 & ~n4912;
  assign n4686 = ~n4685 & ~n4912;
  assign n4820 = n4794 & REG3_REG_10__SCAN_IN;
  assign n4806 = ~n4829 & ~n4912;
  assign n5559 = ~n5558 | ~n5557;
  assign n4852 = ~n4829 | ~n4828;
  assign n4829 = ~n4805 & ~n4804;
  assign n4720 = ~n4719 | ~n5510;
  assign n4634 = ~n4662 | ~n4633;
  assign n4684 = ~n4662 | ~n4661;
  assign n5513 = ~REG2_REG_1__SCAN_IN | ~n5622;
  assign n4749 = ~n4718 | ~n4504;
  assign n5494 = ~REG1_REG_1__SCAN_IN | ~n5622;
  assign n6688 = ~STATE_REG_SCAN_IN & ~n6624;
  assign n7629 = ~n5032 & ~STATE_REG_SCAN_IN;
  assign n4390 = ~n4389 | ~n4960;
  assign n4384 = ~n4380 | ~n4379;
  assign n4608 = ~n4607 | ~n4606;
  assign U3149 = ~STATE_REG_SCAN_IN;
  assign n4393 = ~IR_REG_19__SCAN_IN;
  assign n4984 = ~IR_REG_15__SCAN_IN & ~IR_REG_16__SCAN_IN;
  assign n4557 = ~IR_REG_31__SCAN_IN | ~IR_REG_0__SCAN_IN;
  assign n4411 = ~n4449 | ~n4393;
  assign n4449 = ~n4911 & ~n4392;
  assign n5581 = n4432 ^ n4436;
  assign n4432 = ~n4431 | ~IR_REG_31__SCAN_IN;
  assign n6123 = ~n4506 | ~n4510;
  assign n6130 = ~n4511 & ~n4510;
  assign n6985 = n5581 | n7501;
  assign n4741 = n4737 ^ n7775;
  assign n4763 = n4760 ^ n5272;
  assign n4839 = ~n4836 ^ n7775;
  assign n4908 = ~n4905;
  assign n6573 = ~n6572 ^ n7045;
  assign n5051 = ~n7144;
  assign n4740 = ~n4742;
  assign n6085 = n6151 ^ n6139;
  assign n6502 = n6680 ^ n6679;
  assign n4716 = ~n6014 & ~n4712;
  assign n4714 = ~n6012;
  assign n4854 = ~n4852;
  assign n4754 = ~n4805;
  assign n7175 = ~n7173 | ~n7178;
  assign n7173 = ~n7172 | ~n7171;
  assign n6997 = ~n7219 | ~n7213;
  assign n6569 = ~n5161;
  assign n5018 = ~n5014 ^ n7775;
  assign n4864 = ~n4879;
  assign n5178 = ~n6887;
  assign n5174 = ~n6742;
  assign n5162 = ~n6395;
  assign n5059 = ~n7058;
  assign n6444 = ~n6443 ^ n6449;
  assign n5147 = ~n6335;
  assign n5050 = ~n6196;
  assign n4905 = n4544 ^ n7775;
  assign n4792 = n4788 ^ n7775;
  assign n4817 = n4811 ^ n7775;
  assign n7786 = n5214 ^ n7775;
  assign n7774 = ~n7778 | ~n7779;
  assign n7782 = ~n7778 | ~n7777;
  assign n4766 = ~n4763;
  assign n5287 = ~n7325 | ~n7779;
  assign n5294 = n5286 ^ n7775;
  assign n5284 = ~n7325 | ~n7772;
  assign n4676 = ~n4675;
  assign n4880 = ~n4878;
  assign n4884 = ~n4875 ^ n7775;
  assign n4841 = ~n4840;
  assign n4842 = ~n4839;
  assign n4617 = ~n4619;
  assign n4969 = n4966 ^ n7775;
  assign n6916 = ~n4969 ^ n4970;
  assign n4997 = ~n4994 ^ n7775;
  assign n7100 = ~n7099 | ~n7098;
  assign n7050 = ~n7049 | ~n7048;
  assign n7108 = ~n7176;
  assign n4655 = ~n5856;
  assign n5624 = REG2_REG_1__SCAN_IN ^ n5622;
  assign n5727 = n5726 ^ n5496;
  assign n5708 = REG1_REG_5__SCAN_IN ^ n5722;
  assign n5713 = REG2_REG_5__SCAN_IN ^ n5722;
  assign n5692 = n5704 ^ n5501;
  assign n5696 = n5704 ^ n5520;
  assign n5895 = REG1_REG_9__SCAN_IN ^ n6091;
  assign n7282 = ~n7527;
  assign n6797 = ~n6806;
  assign n7065 = ~n7166;
  assign n6612 = ~n6637;
  assign n7335 = ~n7438 ^ n7334;
  assign n7327 = ~n7309 & ~n7308;
  assign n6932 = ~n7287;
  assign n5186 = ~n7268;
  assign n6905 = ~n6754 & ~n7273;
  assign n6655 = ~n6654 | ~n7503;
  assign n6653 = n6652 ^ n7020;
  assign n6662 = ~n6700 & ~n6598;
  assign n5165 = ~n5164;
  assign n6563 = ~n6395 & ~n6396;
  assign n6458 = ~n6383 & ~n6382;
  assign n4732 = ~DATAI_7_;
  assign n5962 = ~n5961 ^ n6984;
  assign n4743 = ~n4741;
  assign n4903 = n4905 ^ n4906;
  assign n6333 = ~n4817 ^ n4815;
  assign n7406 = ~n5226 ^ n7775;
  assign n7405 = ~n5238;
  assign n4923 = ~n4922;
  assign n4947 = ~n4944;
  assign n4831 = ~DATAI_11_;
  assign n5315 = ~n5314;
  assign n5320 = ~n6123;
  assign n4723 = ~REG1_REG_7__SCAN_IN;
  assign n4717 = ~REG2_REG_7__SCAN_IN;
  assign n4724 = ~REG0_REG_7__SCAN_IN;
  assign n5633 = REG1_REG_1__SCAN_IN ^ n5622;
  assign n5735 = n5726 ^ n5515;
  assign n5504 = REG1_REG_7__SCAN_IN ^ n5767;
  assign n5907 = REG2_REG_9__SCAN_IN ^ n6091;
  assign n6095 = n6151 ^ n6150;
  assign n6318 = n6357 ^ n6348;
  assign n6512 = n6680 ^ n6672;
  assign n7627 = n7626 ^ n7625;
  assign n7625 = ~n7636 ^ REG1_REG_19__SCAN_IN;
  assign n5066 = ~n6651 & ~n7068;
  assign n7758 = n7749 ^ n7748;
  assign n6527 = n6371 ^ n6372;
  assign n6237 = ~n6221 ^ n7003;
  assign n6249 = n6114 ^ n6113;
  assign n4911 = ~n4388 | ~n4730;
  assign n4828 = ~IR_REG_10__SCAN_IN;
  assign n4729 = ~IR_REG_6__SCAN_IN;
  assign n4606 = ~IR_REG_1__SCAN_IN;
  assign n4719 = ~n4718 | ~REG3_REG_6__SCAN_IN;
  assign n7805 = ~n7818 | ~n7787;
  assign n4870 = ~DATAI_13_;
  assign n6087 = ~n6086 | ~n6140;
  assign n6148 = ~n6147 | ~n6146;
  assign n6146 = ~n6145 | ~n6305;
  assign n6505 = ~n7637 | ~n6680;
  assign n7621 = n7619 ^ n7618;
  assign n7077 = ~n7121 | ~n7071;
  assign n7204 = ~n7135 | ~n7134;
  assign n7088 = ~n7174;
  assign n7083 = ~n7082 | ~n7081;
  assign n7004 = ~n6372;
  assign n7193 = ~n7013;
  assign n4878 = n4861 ^ n7775;
  assign n4814 = ~n6332;
  assign n5293 = ~n5273 ^ n5272;
  assign n5270 = ~n7308 | ~n7772;
  assign n7207 = ~n7206 & ~n7205;
  assign n7208 = ~n7175 | ~n7174;
  assign n7029 = ~n7028 & ~n7713;
  assign n7192 = ~n5043;
  assign n7581 = ~n7579 | ~n7722;
  assign n6892 = ~n7001;
  assign n6744 = ~n7024;
  assign n6650 = ~n7124;
  assign n6373 = ~n7056 ^ n7004;
  assign n6163 = ~n6264;
  assign n5042 = ~n7185;
  assign n4865 = ~n6474;
  assign n5259 = ~n5255 ^ n7775;
  assign n5256 = ~n7359 | ~n7779;
  assign n4745 = ~n6203;
  assign n4582 = ~n4581 & ~n4580;
  assign n5234 = ~n5221 ^ n5272;
  assign n5219 = ~n7273 | ~n7772;
  assign n5222 = ~n7273 | ~n7779;
  assign n5223 = ~n7411 | ~n7777;
  assign n4944 = n4941 ^ n7775;
  assign n7515 = ~n7514;
  assign n4645 = n4642 ^ n7775;
  assign n6267 = n4792 ^ n4791;
  assign n5533 = ~n4588 | ~n4587;
  assign n5249 = n5246 ^ n7775;
  assign n4609 = ~DATAI_2_;
  assign n5135 = ~n6016;
  assign n4495 = n5469 & n5471;
  assign n5290 = ~n7550;
  assign n5313 = ~n5310 ^ n7775;
  assign n4922 = ~n4919 ^ n5272;
  assign n4924 = ~n4910 | ~n4909;
  assign n4907 = ~n4906;
  assign n5771 = n5902 ^ n5890;
  assign n6144 = REG1_REG_11__SCAN_IN ^ n6314;
  assign n6308 = n6357 ^ n6356;
  assign n6361 = REG1_REG_13__SCAN_IN ^ n6508;
  assign n6684 = REG1_REG_15__SCAN_IN ^ n6868;
  assign n6862 = n7387 ^ n7386;
  assign n7391 = REG1_REG_17__SCAN_IN ^ n7463;
  assign n7457 = n7622 ^ REG1_REG_18__SCAN_IN;
  assign n7520 = ~REG3_REG_24__SCAN_IN ^ n5261;
  assign n7300 = ~n7332;
  assign n7303 = ~n7321;
  assign n6895 = ~n7411;
  assign n6714 = ~n6712;
  assign n6651 = ~n6605 & ~n7166;
  assign n6791 = ~n6832;
  assign n5062 = ~n7064;
  assign n6288 = ~n5057 | ~n5056;
  assign n5056 = ~n7132;
  assign n5055 = ~n7149;
  assign n6295 = ~n6322;
  assign n5754 = ~n5741;
  assign n7721 = n7719 ^ n7739;
  assign n7730 = ~n7778 | ~n7722;
  assign n7734 = ~n7659 | ~n7658;
  assign n7653 = ~n7652 | ~n7651;
  assign n7648 = ~n7660 ^ n7646;
  assign n7589 = n7588 ^ n7642;
  assign n7571 = ~n7440 | ~n7439;
  assign n7597 = ~n7507;
  assign n7434 = n7572 ^ n7433;
  assign n7428 = ~n7791 | ~n7503;
  assign n5283 = ~DATAI_25_;
  assign n6934 = ~n6933 ^ n7280;
  assign n7306 = ~n5192 & ~n6964;
  assign n5089 = ~n5090;
  assign n6942 = ~n5188 | ~n5187;
  assign n5189 = ~n7046;
  assign n6894 = ~n6893 ^ n6892;
  assign n6721 = n6720 ^ n6719;
  assign n6782 = ~n6792 & ~n6780;
  assign n6649 = ~n6928;
  assign n6568 = ~n6402 | ~n5163;
  assign n6576 = ~n6575 | ~n6574;
  assign n6400 = ~n6452 | ~n5160;
  assign n7043 = ~n6404;
  assign n6406 = ~n6405 ^ n6404;
  assign n6447 = ~n6446 | ~n6445;
  assign n6279 = ~n5150 | ~n5149;
  assign n5150 = ~n6221 | ~n5148;
  assign n7005 = ~n6467 ^ n6280;
  assign n6223 = n6222 ^ n7003;
  assign n6161 = ~n6160 ^ n6170;
  assign n6102 = ~n6101 ^ n6113;
  assign n6038 = ~n6037 ^ n7036;
  assign n5656 = ~n5662 | ~n5535;
  assign n4485 = ~B_REG_SCAN_IN;
  assign n4381 = ~IR_REG_6__SCAN_IN & ~IR_REG_13__SCAN_IN;
  assign n5505 = ~n5388 | ~n7236;
  assign n5510 = ~REG3_REG_7__SCAN_IN;
  assign n7807 = ~n5218 ^ n5217;
  assign n7349 = n5259 ^ n5258;
  assign n5787 = n4645 ^ n4646;
  assign n5789 = ~n5759;
  assign n7792 = ~n7780;
  assign n7814 = ~n7812;
  assign n7811 = ~n7807 & ~n7806;
  assign n7818 = ~n7784 ^ n7783;
  assign n7783 = ~n7782 | ~n7781;
  assign n7784 = ~n7776 ^ n7775;
  assign n4748 = ~REG3_REG_8__SCAN_IN;
  assign n6208 = ~n6207 | ~n7808;
  assign n6207 = ~n6206 | ~n6205;
  assign n5749 = ~n5794;
  assign n5663 = ~n5190;
  assign n7417 = ~n6904;
  assign n5296 = ~n5294;
  assign n6918 = n6917 ^ n6916;
  assign n6554 = ~n6552;
  assign n6954 = ~n5249 ^ n5250;
  assign n6427 = ~n6426 ^ n6425;
  assign n6429 = ~n6422 | ~n7790;
  assign n4593 = ~n5641;
  assign n4620 = ~n4618;
  assign n6829 = ~n4973 | ~n4972;
  assign n4973 = ~n6917 | ~n6916;
  assign n4971 = ~n4969;
  assign n6828 = n4997 ^ n4998;
  assign n4502 = ~REG3_REG_5__SCAN_IN;
  assign n6014 = ~n6000 | ~n4696;
  assign n6011 = ~n4713;
  assign n6633 = ~n4924 ^ n4922;
  assign n7116 = n7114 ^ n7636;
  assign n5322 = ~n5436 | ~REG0_REG_28__SCAN_IN;
  assign n6919 = n6914 ^ n4974;
  assign n4930 = ~REG2_REG_16__SCAN_IN;
  assign n4823 = ~REG2_REG_11__SCAN_IN;
  assign n4797 = ~REG2_REG_10__SCAN_IN;
  assign n6063 = ~n4703 & ~n4702;
  assign n4572 = ~n6127 & ~n4571;
  assign n5563 = REG1_REG_2__SCAN_IN ^ n5571;
  assign n5558 = n5571 ^ REG2_REG_2__SCAN_IN;
  assign n5593 = n5600 ^ n5517;
  assign n5589 = n5600 ^ n5498;
  assign n5782 = n5902 ^ n5901;
  assign n6432 = ~REG3_REG_11__SCAN_IN | ~U3149;
  assign n6156 = REG2_REG_11__SCAN_IN ^ n6314;
  assign n6352 = REG2_REG_13__SCAN_IN ^ n6508;
  assign n6676 = REG2_REG_15__SCAN_IN ^ n6868;
  assign n6872 = n7387 ^ n7378;
  assign n7382 = REG2_REG_17__SCAN_IN ^ n7463;
  assign n7468 = n7622 ^ REG2_REG_18__SCAN_IN;
  assign n7540 = ~n6991;
  assign n7795 = REG3_REG_28__SCAN_IN ^ n6122;
  assign n7596 = n5329 ^ n5319;
  assign n7705 = n5301 ^ n5300;
  assign n7558 = REG3_REG_25__SCAN_IN ^ n5276;
  assign n7322 = ~n7284 | ~n7283;
  assign n7284 = ~n7281 | ~n7280;
  assign n7476 = ~n6974;
  assign n6648 = ~n5170 | ~n5169;
  assign n5170 = ~n5168 | ~n7034;
  assign n6647 = ~n7071;
  assign n6847 = ~n7668 | ~n6919;
  assign n6625 = ~n6624 ^ n4927;
  assign n6450 = ~n5157 | ~n5156;
  assign n5157 = ~n6371 | ~n5155;
  assign n6452 = ~n5159 | ~n7041;
  assign n5159 = ~n6450;
  assign n6421 = ~REG3_REG_11__SCAN_IN ^ n4820;
  assign n6289 = n6288 ^ n7005;
  assign n7830 = ~n7750;
  assign n5886 = ~n5130 | ~n5129;
  assign n5128 = ~n5826;
  assign n6983 = ~n7201 | ~n7140;
  assign n4654 = ~n4653 | ~n4652;
  assign n4481 = ~n4480 | ~n4479;
  assign n7824 = n7541 ^ n7540;
  assign n7831 = n7539 ^ n7538;
  assign n7679 = ~n7660 ^ n7734;
  assign n7671 = ~n7749;
  assign n7477 = n7572 ^ n7571;
  assign n7370 = n7438 ^ n7437;
  assign n7326 = ~n7327;
  assign n7341 = ~n7340 | ~n7339;
  assign n6975 = n7281 ^ n7280;
  assign n6976 = ~n7306 ^ n7305;
  assign n6879 = n6942 ^ n5189;
  assign n6906 = ~n6905 ^ n6904;
  assign n6806 = n6778 ^ n6788;
  assign n6637 = n6597 ^ n7034;
  assign n6600 = ~n6700 | ~n6598;
  assign n6586 = n6568 ^ n7045;
  assign n6587 = ~n6563 ^ n6562;
  assign n6398 = ~n7542 | ~n6397;
  assign n6517 = n6458 ^ n6457;
  assign n6378 = ~n6467 | ~n7722;
  assign n6385 = ~n7542 | ~n6384;
  assign n6384 = ~n6383 | ~n6382;
  assign n6322 = ~n6279 ^ n7005;
  assign n6324 = n6383 & n6283;
  assign n6238 = n6216 ^ n6335;
  assign n6182 = n6174 & n6216;
  assign n6185 = n6171 ^ n6170;
  assign n6052 = ~n6036 ^ n7036;
  assign n5981 = ~n5960 ^ n6984;
  assign n5969 = ~n5962 | ~n7647;
  assign n5875 = ~n5870 | ~n7647;
  assign n5854 = ~n5823 | ~n5822;
  assign n5950 = ~n5923 | ~n5922;
  assign n5954 = ~n5936 | ~n5935;
  assign n5535 = ~n5658;
  assign n7239 = ~n4405 ^ IR_REG_23__SCAN_IN;
  assign n4392 = ~n4391 | ~n4984;
  assign n4391 = ~n4390 & ~IR_REG_14__SCAN_IN;
  assign n4957 = ~IR_REG_16__SCAN_IN;
  assign n5318 = ~n7807 ^ n7806;
  assign n4889 = n4903 ^ n4904;
  assign n7354 = ~REG3_REG_23__SCAN_IN ^ n5200;
  assign n6334 = ~n6333 ^ n6332;
  assign n6767 = ~REG3_REG_19__SCAN_IN ^ n5026;
  assign n5022 = n7258 ^ n7257;
  assign n4887 = ~n4886;
  assign n6250 = n4749 ^ n4748;
  assign n7410 = ~REG3_REG_21__SCAN_IN ^ n5080;
  assign n7409 = ~n7408 ^ n7407;
  assign n7407 = ~n7406 ^ n7405;
  assign n6528 = REG3_REG_12__SCAN_IN ^ n4844;
  assign n6705 = ~REG3_REG_16__SCAN_IN ^ n4949;
  assign n6699 = ~n6698 ^ n6697;
  assign n6006 = ~n4679 ^ REG3_REG_5__SCAN_IN;
  assign n5841 = ~n5816;
  assign n7266 = ~REG3_REG_20__SCAN_IN ^ n5072;
  assign n6557 = n6556 ^ n6555;
  assign n6959 = ~REG3_REG_22__SCAN_IN ^ n5096;
  assign n4529 = ~n4888 | ~n7650;
  assign n6831 = n4975 ^ n5005;
  assign n4975 = ~REG3_REG_18__SCAN_IN;
  assign n6830 = n6829 ^ n6828;
  assign n6021 = ~n4718 ^ REG3_REG_6__SCAN_IN;
  assign n7695 = ~n7694 ^ n7693;
  assign n7694 = ~n7690;
  assign n6634 = n6633 ^ n6632;
  assign n6990 = ~n5438 | ~n5437;
  assign n6133 = ~n6132 | ~n6131;
  assign n6834 = ~n7267;
  assign n6654 = ~n6915;
  assign n5879 = ~n6063;
  assign n6022 = ~n5965;
  assign n5991 = ~n5871;
  assign n4406 = ~n5395;
  assign n6353 = ~n7383 | ~n6509;
  assign n6689 = ~n7631 | ~ADDR_REG_15__SCAN_IN;
  assign n6867 = ~n6858 | ~n6857;
  assign n7673 = ~n7795 | ~n7668;
  assign n7497 = n7322 ^ n7321;
  assign n7251 = ~n7245;
  assign n6825 = n6888 ^ n7024;
  assign n6775 = n6741 ^ n6719;
  assign n6790 = ~n6789 ^ n6788;
  assign n6844 = ~n6648 ^ n7020;
  assign n6606 = ~n6605 ^ n7034;
  assign n6414 = ~REG3_REG_14__SCAN_IN ^ n4890;
  assign n6416 = ~REG2_REG_14__SCAN_IN | ~n7832;
  assign n6548 = ~n6355 ^ n4505;
  assign n6340 = ~REG3_REG_10__SCAN_IN ^ n4794;
  assign n6233 = ~n6237 | ~n6779;
  assign n6276 = n4771 ^ REG3_REG_9__SCAN_IN;
  assign n6257 = ~n6249 | ~n6248;
  assign n5745 = ~n5744 | ~n5743;
  assign n5946 = ~n5945 | ~n5944;
  assign n5944 = ~n5950 | ~n7496;
  assign n7761 = ~n7760 & ~n7759;
  assign n5831 = ~n5828 | ~n5827;
  assign n5808 = ~n5805 | ~n5804;
  assign n5383 = ~n4443 | ~n4442;
  assign n4439 = ~n4443 & ~n4912;
  assign n7236 = ~n7239 | ~STATE_REG_SCAN_IN;
  assign n7176 = ~n4417 ^ IR_REG_21__SCAN_IN;
  assign n4417 = ~n4416 | ~IR_REG_31__SCAN_IN;
  assign n7115 = n4415 ^ n4414;
  assign n7622 = ~n4989 ^ IR_REG_18__SCAN_IN;
  assign n7463 = n4961 ^ n4960;
  assign n6868 = n4913 ^ IR_REG_15__SCAN_IN;
  assign n4522 = ~IR_REG_14__SCAN_IN;
  assign n6508 = ~n4869 ^ IR_REG_13__SCAN_IN;
  assign n6314 = n4830 ^ n4853;
  assign n4781 = ~IR_REG_9__SCAN_IN;
  assign n5767 = n4731 ^ n4802;
  assign n5704 = n4704 ^ IR_REG_6__SCAN_IN;
  assign n5722 = n4686 ^ IR_REG_5__SCAN_IN;
  assign n5600 = n4684 ^ IR_REG_4__SCAN_IN;
  assign n5726 = n4636 ^ n4635;
  assign n5571 = n4662 ^ n4633;
  assign n5622 = ~n4557 ^ IR_REG_1__SCAN_IN;
  assign n6077 = ~n6076 | ~n6206;
  assign n7821 = ~n7820 & ~n7819;
  assign n6158 = ~n6157 | ~n6315;
  assign n6320 = ~n6319 | ~n6349;
  assign n5978 = ~n5977 | ~n5976;
  assign n6060 = ~n7767 | ~n6059;
  assign n5986 = ~n7767 | ~n5988;
  assign n5919 = ~n7767 | ~n5918;
  assign n6057 = ~n7763 | ~n6059;
  assign n5989 = ~n7763 | ~n5988;
  assign n5916 = ~n7763 | ~n5918;
  assign n7649 = ~n7503;
  assign n4579 = ~REG1_REG_0__SCAN_IN;
  assign n4567 = ~REG2_REG_0__SCAN_IN;
  assign n7184 = ~n7178;
  assign n4378 = n7555 | n7554;
  assign n4607 = ~IR_REG_0__SCAN_IN;
  assign n7009 = ~n7007;
  assign n7139 = ~n7138;
  assign n4765 = ~n4764;
  assign n4856 = ~DATAI_12_;
  assign n4783 = ~DATAI_9_;
  assign n5210 = ~DATAI_27_;
  assign n4637 = ~DATAI_3_;
  assign n4946 = ~n4945;
  assign n4770 = ~n4769;
  assign n5173 = ~n6648 | ~n5171;
  assign n4503 = ~REG3_REG_6__SCAN_IN;
  assign n5100 = ~REG0_REG_23__SCAN_IN;
  assign n4952 = ~REG2_REG_17__SCAN_IN;
  assign n5819 = ~n5927;
  assign n7311 = ~n7491;
  assign n4448 = ~n5505;
  assign n7232 = ~n7236;
  assign n4380 = ~IR_REG_12__SCAN_IN & ~IR_REG_11__SCAN_IN;
  assign n4379 = ~IR_REG_10__SCAN_IN & ~IR_REG_8__SCAN_IN;
  assign n4382 = ~IR_REG_9__SCAN_IN & ~IR_REG_7__SCAN_IN;
  assign n4383 = ~n4382 | ~n4381;
  assign n4386 = ~IR_REG_1__SCAN_IN & ~IR_REG_4__SCAN_IN;
  assign n4385 = ~IR_REG_5__SCAN_IN & ~IR_REG_0__SCAN_IN;
  assign n4387 = ~n4386 | ~n4385;
  assign n4635 = ~IR_REG_3__SCAN_IN;
  assign n4660 = ~n4633 | ~n4635;
  assign n4730 = ~n4387 & ~n4660;
  assign n4414 = ~IR_REG_20__SCAN_IN;
  assign n4395 = ~n4394 | ~n4414;
  assign n4407 = ~n4411 & ~n4395;
  assign n4404 = ~n4407 | ~n4396;
  assign n4401 = ~n4404 & ~IR_REG_23__SCAN_IN;
  assign n4399 = ~n4401 | ~n4397;
  assign n4427 = ~n4399 & ~IR_REG_25__SCAN_IN;
  assign n4398 = ~n4427 & ~n4912;
  assign n4400 = ~n4399 | ~IR_REG_31__SCAN_IN;
  assign n4402 = ~n4401 & ~n4912;
  assign n4405 = ~n4404 | ~IR_REG_31__SCAN_IN;
  assign n5395 = ~n7239 & ~U3149;
  assign n4408 = ~n4407 & ~n4912;
  assign n4410 = ~n7238 | ~STATE_REG_SCAN_IN;
  assign n4409 = ~DATAI_22_ | ~U3149;
  assign U3330 = ~n4410 | ~n4409;
  assign n4413 = ~n7115 | ~STATE_REG_SCAN_IN;
  assign n4412 = ~DATAI_20_ | ~U3149;
  assign U3332 = ~n4413 | ~n4412;
  assign n4419 = ~n7176 | ~STATE_REG_SCAN_IN;
  assign n4418 = ~DATAI_21_ | ~U3149;
  assign U3331 = ~n4419 | ~n4418;
  assign n4421 = ~n4492 | ~STATE_REG_SCAN_IN;
  assign n4420 = ~DATAI_24_ | ~U3149;
  assign U3328 = ~n4421 | ~n4420;
  assign n4423 = ~n4490 | ~STATE_REG_SCAN_IN;
  assign n4422 = ~DATAI_25_ | ~U3149;
  assign U3327 = ~n4423 | ~n4422;
  assign n4425 = ~n5392 | ~STATE_REG_SCAN_IN;
  assign n4424 = ~DATAI_26_ | ~U3149;
  assign U3326 = ~n4425 | ~n4424;
  assign n4438 = ~n4427 | ~n4426;
  assign n4429 = ~n7501 | ~STATE_REG_SCAN_IN;
  assign n4428 = ~DATAI_27_ | ~U3149;
  assign U3325 = ~n4429 | ~n4428;
  assign n4431 = ~n4430 | ~n4435;
  assign n4434 = ~n5581 | ~STATE_REG_SCAN_IN;
  assign n4433 = ~DATAI_28_ | ~U3149;
  assign U3324 = ~n4434 | ~n4433;
  assign n4437 = ~n4436 | ~n4435;
  assign n4443 = ~n4438 & ~n4437;
  assign n4441 = ~n4510 | ~STATE_REG_SCAN_IN;
  assign n4440 = ~DATAI_29_ | ~U3149;
  assign U3323 = ~n4441 | ~n4440;
  assign n4446 = ~n4506 | ~STATE_REG_SCAN_IN;
  assign n4445 = ~DATAI_30_ | ~U3149;
  assign U3322 = ~n4446 | ~n4445;
  assign n4447 = ~n5105 & ~n7239;
  assign n5506 = ~n6996 & ~n4447;
  assign n7631 = ~n5506 & ~n4448;
  assign U4043 = ~n6193;
  assign U3148 = ~n7631 & ~U4043;
  assign n4450 = ~n4449 & ~n4912;
  assign n7636 = n4450 ^ IR_REG_19__SCAN_IN;
  assign n5401 = ~n7108 | ~n4527;
  assign n7725 = ~n5474 | ~n7115;
  assign n4454 = ~n7234 & ~n7650;
  assign n4452 = ~n5401 & ~n7485;
  assign n4453 = ~n4452 & ~n5095;
  assign n4456 = ~D_REG_12__SCAN_IN & ~D_REG_13__SCAN_IN;
  assign n4455 = ~D_REG_10__SCAN_IN & ~D_REG_11__SCAN_IN;
  assign n4460 = ~n4456 | ~n4455;
  assign n4458 = ~D_REG_8__SCAN_IN & ~D_REG_9__SCAN_IN;
  assign n4457 = ~D_REG_6__SCAN_IN & ~D_REG_7__SCAN_IN;
  assign n4459 = ~n4458 | ~n4457;
  assign n4482 = n4460 | n4459;
  assign n4462 = ~D_REG_4__SCAN_IN & ~D_REG_5__SCAN_IN;
  assign n4461 = ~D_REG_2__SCAN_IN & ~D_REG_3__SCAN_IN;
  assign n4463 = ~n4462 | ~n4461;
  assign n4480 = ~n4463 & ~D_REG_29__SCAN_IN;
  assign n4465 = ~D_REG_28__SCAN_IN & ~D_REG_31__SCAN_IN;
  assign n4464 = ~D_REG_26__SCAN_IN & ~D_REG_27__SCAN_IN;
  assign n4469 = ~n4465 | ~n4464;
  assign n4467 = ~D_REG_15__SCAN_IN & ~D_REG_17__SCAN_IN;
  assign n4466 = ~D_REG_16__SCAN_IN & ~D_REG_14__SCAN_IN;
  assign n4468 = ~n4467 | ~n4466;
  assign n4477 = ~n4469 & ~n4468;
  assign n4471 = ~D_REG_24__SCAN_IN & ~D_REG_25__SCAN_IN;
  assign n4470 = ~D_REG_22__SCAN_IN & ~D_REG_23__SCAN_IN;
  assign n4475 = ~n4471 | ~n4470;
  assign n4473 = ~D_REG_20__SCAN_IN & ~D_REG_21__SCAN_IN;
  assign n4472 = ~D_REG_18__SCAN_IN & ~D_REG_19__SCAN_IN;
  assign n4474 = ~n4473 | ~n4472;
  assign n4476 = ~n4475 & ~n4474;
  assign n4478 = ~n4477 | ~n4476;
  assign n4479 = ~n4478 & ~D_REG_30__SCAN_IN;
  assign n5387 = ~n4488 | ~n5392;
  assign n5468 = n4489 | n5387;
  assign n5469 = ~n4491 & ~n5396;
  assign n5471 = ~n4494 & ~n4493;
  assign n4499 = ~n4584;
  assign n4497 = ~n7239;
  assign n4498 = ~n5112 | ~n4497;
  assign n4500 = ~n4499 & ~n4498;
  assign n7794 = ~n5532 & ~U3149;
  assign n4521 = ~n7521 & ~n6414;
  assign n4516 = n6548 | n6123;
  assign n4511 = ~n4506;
  assign n6125 = ~n4511 | ~n4510;
  assign n5324 = ~n6130;
  assign n4513 = ~n5324 & ~n4512;
  assign n4517 = ~n7234;
  assign n4518 = ~n4898;
  assign n5583 = ~n5581;
  assign n7790 = ~n4518 & ~n5583;
  assign n4519 = ~n6407 | ~n7790;
  assign n6498 = ~REG3_REG_14__SCAN_IN | ~U3149;
  assign n4520 = ~n4519 | ~n6498;
  assign n4531 = ~n4521 & ~n4520;
  assign n4525 = ~n6985 | ~DATAI_14_;
  assign n4523 = ~n4911 | ~IR_REG_31__SCAN_IN;
  assign n4524 = ~n6996 | ~n6680;
  assign n6395 = ~n4525 | ~n4524;
  assign n7700 = ~n4529 | ~n7746;
  assign n4530 = ~n6395 | ~n7700;
  assign n4902 = ~n4531 | ~n4530;
  assign n4538 = n6414 | n6123;
  assign n4535 = ~n5324 & ~n4534;
  assign n6627 = ~n4538 | ~n4537;
  assign n5657 = ~n7176 | ~n4539;
  assign n5211 = ~n4584 | ~n5657;
  assign n7772 = ~n5211;
  assign n7542 = ~n5401 & ~n7115;
  assign n4547 = ~REG2_REG_1__SCAN_IN;
  assign n4550 = ~n5324 & ~n4547;
  assign n4548 = ~REG0_REG_1__SCAN_IN;
  assign n4551 = ~REG3_REG_1__SCAN_IN;
  assign n4552 = ~REG1_REG_1__SCAN_IN;
  assign n5924 = ~n4556 | ~n4555;
  assign n4562 = ~n5924 | ~n7779;
  assign n4560 = n6996 & n5622;
  assign n4558 = ~DATAI_1_;
  assign n4559 = ~n6996 & ~n4558;
  assign n5190 = ~n4560 & ~n4559;
  assign n4561 = ~n5663 | ~n7772;
  assign n4563 = ~n4562 | ~n4561;
  assign n5641 = n4563 ^ n7775;
  assign n4565 = ~n5924 | ~n7777;
  assign n4564 = ~n5663 | ~n7779;
  assign n4592 = ~n5641 & ~n4566;
  assign n4569 = ~n5324 & ~n4567;
  assign n4568 = ~n6125 & ~n4579;
  assign n4570 = ~REG3_REG_0__SCAN_IN;
  assign n4573 = ~n6123 & ~n4570;
  assign n4571 = ~REG0_REG_0__SCAN_IN;
  assign n5662 = ~n4575 | ~n4574;
  assign n4583 = ~n5662 | ~n7779;
  assign n4578 = n6996 & IR_REG_0__SCAN_IN;
  assign n4576 = ~DATAI_0_;
  assign n4577 = ~n6996 & ~n4576;
  assign n5658 = ~n4578 & ~n4577;
  assign n4581 = ~n5658 & ~n5211;
  assign n4580 = ~n4584 & ~n4579;
  assign n4588 = ~n5662 | ~n7777;
  assign n4586 = ~n5658 & ~n5209;
  assign n4585 = ~n4584 & ~n4607;
  assign n4587 = ~n4586 & ~n4585;
  assign n4590 = ~n4589 & ~n5272;
  assign n5639 = ~n4591 & ~n4590;
  assign n5614 = ~n4595 & ~n4594;
  assign n4596 = ~REG2_REG_2__SCAN_IN;
  assign n4599 = ~n5324 & ~n4596;
  assign n4597 = ~REG3_REG_2__SCAN_IN;
  assign n4598 = ~n6123 & ~n4597;
  assign n4605 = ~n4599 & ~n4598;
  assign n4600 = ~REG1_REG_2__SCAN_IN;
  assign n4603 = ~n6125 & ~n4600;
  assign n4601 = ~REG0_REG_2__SCAN_IN;
  assign n4602 = ~n6127 & ~n4601;
  assign n4604 = ~n4603 & ~n4602;
  assign n5794 = ~n4605 | ~n4604;
  assign n4613 = ~n5794 | ~n7779;
  assign n4662 = ~n4608 | ~IR_REG_31__SCAN_IN;
  assign n4611 = n6996 & n5571;
  assign n4610 = ~n6996 & ~n4609;
  assign n5124 = ~n4611 & ~n4610;
  assign n4612 = ~n5937 | ~n7772;
  assign n4616 = ~n5794 | ~n7777;
  assign n4615 = ~n5937 | ~n7779;
  assign n5617 = ~n5614 | ~n5613;
  assign n5786 = ~n5617 | ~n4623;
  assign n4624 = ~REG2_REG_3__SCAN_IN;
  assign n4626 = ~n5324 & ~n4624;
  assign n4627 = ~REG1_REG_3__SCAN_IN;
  assign n4628 = ~REG0_REG_3__SCAN_IN;
  assign n5927 = ~n4632 | ~n4631;
  assign n4641 = ~n5927 | ~n7779;
  assign n4639 = n6996 & n5726;
  assign n4638 = ~n6996 & ~n4637;
  assign n5759 = ~n4639 & ~n4638;
  assign n4640 = ~n5789 | ~n7772;
  assign n4644 = ~n5927 | ~n7777;
  assign n4643 = ~n5789 | ~n7779;
  assign n4649 = ~n5786 & ~n5787;
  assign n5845 = ~n4649 & ~n4648;
  assign n4653 = ~REG3_REG_3__SCAN_IN;
  assign n4652 = ~REG3_REG_4__SCAN_IN;
  assign n4656 = ~n6130 | ~REG2_REG_4__SCAN_IN;
  assign n4664 = ~n6985 | ~DATAI_4_;
  assign n4661 = ~n4660 | ~IR_REG_31__SCAN_IN;
  assign n4663 = ~n6996 | ~n5600;
  assign n5847 = ~n5845 | ~n5844;
  assign n5998 = ~n5847 | ~n4676;
  assign n4680 = ~n6130 | ~REG2_REG_5__SCAN_IN;
  assign n4688 = ~n6985 | ~DATAI_5_;
  assign n4687 = ~n6996 | ~n5722;
  assign n6000 = ~n5998 | ~n5997;
  assign n4700 = ~n6130 | ~REG2_REG_6__SCAN_IN;
  assign n4706 = ~n6985 | ~DATAI_6_;
  assign n4704 = ~n4730 & ~n4912;
  assign n4705 = ~n6996 | ~n5704;
  assign n6074 = ~n4716 & ~n4715;
  assign n4722 = ~n5324 & ~n4717;
  assign n4805 = ~n4730 | ~n4729;
  assign n4734 = n6996 & n5767;
  assign n4733 = ~n6996 & ~n4732;
  assign n6206 = ~n6074 | ~n6073;
  assign n4750 = ~n6130 | ~REG2_REG_8__SCAN_IN;
  assign n4757 = ~n6985 | ~DATAI_8_;
  assign n4756 = ~n6996 | ~n5902;
  assign n6202 = ~n4768 | ~n6204;
  assign n6268 = ~n6202 | ~n4770;
  assign n4774 = ~n6130 | ~REG2_REG_9__SCAN_IN;
  assign n6224 = ~n4777 & ~n4776;
  assign n4785 = n6996 & n6091;
  assign n4784 = ~n6996 & ~n4783;
  assign n6264 = ~n4785 & ~n4784;
  assign n6270 = ~n6268 | ~n6267;
  assign n6332 = ~n6270 | ~n4793;
  assign n4801 = n6340 | n6123;
  assign n4798 = ~n5324 & ~n4797;
  assign n4808 = ~n6985 | ~DATAI_10_;
  assign n4807 = ~n6996 | ~n6151;
  assign n6335 = ~n4808 | ~n4807;
  assign n4827 = n6421 | n6123;
  assign n4824 = ~n5324 & ~n4823;
  assign n4833 = n6996 & n6314;
  assign n4832 = ~n6996 & ~n4831;
  assign n6280 = ~n4833 & ~n4832;
  assign n4843 = ~n6426 & ~n6424;
  assign n6476 = ~n4843 & ~n6423;
  assign n4848 = ~n5324 & ~n4847;
  assign n4858 = n6996 & n6357;
  assign n4857 = ~n6996 & ~n4856;
  assign n6470 = ~n4858 & ~n4857;
  assign n4872 = n6996 & n6508;
  assign n4871 = ~n6996 & ~n4870;
  assign n6539 = ~n4872 & ~n4871;
  assign n4904 = ~n4885 & ~n6551;
  assign n4897 = n6625 | n6123;
  assign n4894 = ~n5324 & ~n4893;
  assign n7788 = ~n4898 | ~n5583;
  assign n4899 = ~n6706 | ~n7532;
  assign U3212 = n4902 | n4901;
  assign n4910 = ~n4904 | ~n4903;
  assign n4987 = ~n4911 & ~IR_REG_14__SCAN_IN;
  assign n4916 = n6996 & n6868;
  assign n4915 = ~n6996 & ~n4914;
  assign n6562 = ~n4916 & ~n4915;
  assign n4926 = ~n6633 | ~n6632;
  assign n4925 = ~n4924 | ~n4923;
  assign n4934 = n6705 | n6123;
  assign n4931 = ~n5324 & ~n4930;
  assign n4938 = ~n6985 | ~DATAI_16_;
  assign n4937 = ~n6996 | ~n7387;
  assign n6700 = ~n4938 | ~n4937;
  assign n6917 = ~n4948 & ~n6696;
  assign n4953 = ~n5324 & ~n4952;
  assign n4963 = ~n6985 | ~DATAI_17_;
  assign n4962 = ~n6996 | ~n7463;
  assign n6924 = ~n4963 | ~n4962;
  assign n4976 = ~REG1_REG_18__SCAN_IN;
  assign n4977 = ~REG0_REG_18__SCAN_IN;
  assign n4980 = ~n6130 | ~REG2_REG_18__SCAN_IN;
  assign n6915 = ~n4983 & ~n4982;
  assign n4991 = ~n6985 | ~DATAI_18_;
  assign n4985 = ~n4984;
  assign n4990 = ~n6996 | ~n7622;
  assign n6792 = ~n4991 | ~n4990;
  assign n5002 = ~n6829 | ~n6828;
  assign n5006 = ~n6130 | ~REG2_REG_19__SCAN_IN;
  assign n7267 = ~n5009 & ~n5008;
  assign n5013 = ~n7267 & ~n5209;
  assign n5011 = ~n6985 | ~DATAI_19_;
  assign n5010 = ~n6996 | ~n7636;
  assign n6722 = ~n5011 | ~n5010;
  assign n5012 = ~n6731 & ~n5211;
  assign n5016 = ~n6731 & ~n5209;
  assign n5021 = ~n5018;
  assign n5020 = ~n5019;
  assign n5039 = ~n7794 | ~n6767;
  assign n7697 = ~n7790;
  assign n5037 = ~n6915 & ~n7697;
  assign n5025 = n6130 & REG2_REG_20__SCAN_IN;
  assign n5023 = ~REG1_REG_20__SCAN_IN;
  assign n5072 = ~n5026 & ~n5032;
  assign n5027 = ~REG0_REG_20__SCAN_IN;
  assign n5033 = ~n7788 & ~n6895;
  assign n5035 = ~n5033 & ~n7629;
  assign n5034 = ~n7700 | ~n6722;
  assign n5036 = ~n5035 | ~n5034;
  assign n5038 = ~n5037 & ~n5036;
  assign n5040 = ~n5039 | ~n5038;
  assign U3216 = n5041 | n5040;
  assign n5043 = ~n5794 & ~n5124;
  assign n7188 = ~n5749 & ~n5937;
  assign n5929 = ~n5043 & ~n7188;
  assign n7185 = ~n5924 & ~n5190;
  assign n7180 = ~n5121 & ~n5663;
  assign n5044 = ~n5929 | ~n5928;
  assign n5741 = ~n7013 & ~n7008;
  assign n6718 = ~n6789 | ~n7073;
  assign n7286 = ~n5067 | ~n7015;
  assign n5180 = ~n6985 | ~DATAI_20_;
  assign n6893 = ~n6745 | ~n5068;
  assign n5071 = n6130 & REG2_REG_21__SCAN_IN;
  assign n5069 = ~REG1_REG_21__SCAN_IN;
  assign n5073 = ~REG0_REG_21__SCAN_IN;
  assign n6904 = ~n6985 | ~DATAI_21_;
  assign n5082 = n6130 & REG2_REG_22__SCAN_IN;
  assign n5083 = ~REG1_REG_22__SCAN_IN;
  assign n5084 = ~REG0_REG_22__SCAN_IN;
  assign n6943 = ~n6985 | ~DATAI_22_;
  assign n7046 = ~n7084 | ~n7178;
  assign n5093 = ~n7176 | ~n7115;
  assign n5092 = ~n7238 | ~n7636;
  assign n7720 = n5093 & n5092;
  assign n7424 = ~n5581 | ~n5095;
  assign n5109 = ~n5186 & ~n7424;
  assign n5098 = n6130 & REG2_REG_23__SCAN_IN;
  assign n5099 = ~REG1_REG_23__SCAN_IN;
  assign n7503 = ~n5581 & ~n5105;
  assign n5107 = ~n7527 | ~n7503;
  assign n5106 = ~n6964 | ~n7650;
  assign n5108 = ~n5107 | ~n5106;
  assign n5117 = ~n5116 & ~n5115;
  assign n7037 = ~n5929;
  assign n5120 = ~n5924 & ~n5663;
  assign n5122 = ~n5121 & ~n5190;
  assign n5921 = ~n5123 & ~n5122;
  assign n5922 = ~n7037 | ~n5921;
  assign n5125 = ~n5749 | ~n5124;
  assign n5742 = ~n5922 | ~n5125;
  assign n5127 = ~n5742 | ~n5754;
  assign n5130 = ~n5128 | ~n5825;
  assign n5134 = ~n5886 | ~n5131;
  assign n5960 = ~n5134 | ~n5133;
  assign n5138 = ~n5960 | ~n5136;
  assign n6036 = ~n5138 | ~n5137;
  assign n5140 = ~n6036 | ~n7036;
  assign n6114 = ~n5140 | ~n5139;
  assign n5143 = ~n6114 | ~n5141;
  assign n6171 = ~n5143 | ~n5142;
  assign n5146 = ~n6171 | ~n5144;
  assign n6221 = ~n5146 | ~n5145;
  assign n6371 = ~n5154 | ~n5153;
  assign n6402 = ~n6400 | ~n6404;
  assign n7045 = ~n5165 | ~n7064;
  assign n5167 = ~n6568 | ~n7045;
  assign n6597 = ~n5167 | ~n5166;
  assign n6778 = ~n5173 | ~n5172;
  assign n5188 = ~n5185 | ~n5184;
  assign n7740 = ~n5402 | ~n7775;
  assign n5938 = ~n5190 | ~n5658;
  assign n6780 = ~n6663 | ~n6662;
  assign n6754 = ~n6782 | ~n6731;
  assign n5192 = ~n6905 | ~n6904;
  assign n5194 = ~n7746 & ~n6959;
  assign U3268 = n5199 | n5198;
  assign n5329 = ~REG3_REG_27__SCAN_IN;
  assign n5276 = n5261 & REG3_REG_24__SCAN_IN;
  assign n5300 = ~n5276 | ~REG3_REG_25__SCAN_IN;
  assign n5319 = ~n5300 & ~n5301;
  assign n5201 = ~REG1_REG_27__SCAN_IN;
  assign n5204 = ~n6125 & ~n5201;
  assign n5202 = ~REG0_REG_27__SCAN_IN;
  assign n5205 = ~n6130 | ~REG2_REG_27__SCAN_IN;
  assign n7696 = ~n5208 & ~n5207;
  assign n7657 = ~n6996 & ~n5210;
  assign n5212 = ~n7506 & ~n5211;
  assign n5215 = ~n7657 | ~n7779;
  assign n5243 = ~n7258 | ~n5230;
  assign n6955 = ~n5243 | ~n5242;
  assign n6957 = ~n6955 | ~n6954;
  assign n7350 = ~n6957 | ~n5252;
  assign n7305 = ~n6985 | ~DATAI_23_;
  assign n7352 = ~n7350 | ~n7349;
  assign n7518 = ~n7352 | ~n5260;
  assign n5263 = n6130 & REG2_REG_24__SCAN_IN;
  assign n5264 = ~REG1_REG_24__SCAN_IN;
  assign n5265 = ~REG0_REG_24__SCAN_IN;
  assign n7522 = ~n6985 | ~DATAI_24_;
  assign n5274 = ~n7308 | ~n7779;
  assign n5291 = ~n7518 | ~n7514;
  assign n7367 = ~REG2_REG_25__SCAN_IN;
  assign n5279 = ~n5324 & ~n7367;
  assign n7325 = ~n6996 & ~n5283;
  assign n7473 = ~REG2_REG_26__SCAN_IN;
  assign n5304 = ~n5324 & ~n7473;
  assign n7573 = ~n6985 | ~DATAI_26_;
  assign n5308 = ~n7699 | ~n7772;
  assign n5311 = ~n7699 | ~n7779;
  assign n5317 = ~n7690 | ~n7692;
  assign n7806 = ~n5317 | ~n7691;
  assign n7664 = ~REG2_REG_28__SCAN_IN;
  assign n5325 = ~n5324 & ~n7664;
  assign n5337 = ~n7778 | ~n7532;
  assign n5335 = ~n7596 & ~n7521;
  assign n5333 = ~n7579 | ~n7790;
  assign n5331 = ~n7793 & ~n7506;
  assign n5330 = ~n5329 & ~STATE_REG_SCAN_IN;
  assign n5332 = ~n5331 & ~n5330;
  assign n5334 = ~n5333 | ~n5332;
  assign n5336 = ~n5335 & ~n5334;
  assign n5338 = ~n5337 | ~n5336;
  assign U3211 = n5339 | n5338;
  assign n5341 = ~STATE_REG_SCAN_IN | ~IR_REG_0__SCAN_IN;
  assign n5340 = ~DATAI_0_ | ~U3149;
  assign U3352 = ~n5341 | ~n5340;
  assign n5343 = ~STATE_REG_SCAN_IN | ~n5622;
  assign n5342 = ~DATAI_1_ | ~U3149;
  assign U3351 = ~n5343 | ~n5342;
  assign n5345 = ~STATE_REG_SCAN_IN | ~n5571;
  assign n5344 = ~DATAI_2_ | ~U3149;
  assign U3350 = ~n5345 | ~n5344;
  assign n5347 = ~STATE_REG_SCAN_IN | ~n5600;
  assign n5346 = ~DATAI_4_ | ~U3149;
  assign U3348 = ~n5347 | ~n5346;
  assign n5349 = ~STATE_REG_SCAN_IN | ~n5726;
  assign n5348 = ~DATAI_3_ | ~U3149;
  assign U3349 = ~n5349 | ~n5348;
  assign n5351 = ~STATE_REG_SCAN_IN | ~n5704;
  assign n5350 = ~DATAI_6_ | ~U3149;
  assign U3346 = ~n5351 | ~n5350;
  assign n5353 = ~STATE_REG_SCAN_IN | ~n5722;
  assign n5352 = ~DATAI_5_ | ~U3149;
  assign U3347 = ~n5353 | ~n5352;
  assign n5355 = ~STATE_REG_SCAN_IN | ~n5767;
  assign n5354 = ~DATAI_7_ | ~U3149;
  assign U3345 = ~n5355 | ~n5354;
  assign n5357 = ~STATE_REG_SCAN_IN | ~n6680;
  assign n5356 = ~DATAI_14_ | ~U3149;
  assign U3338 = ~n5357 | ~n5356;
  assign n5359 = ~STATE_REG_SCAN_IN | ~n6151;
  assign n5358 = ~DATAI_10_ | ~U3149;
  assign U3342 = ~n5359 | ~n5358;
  assign n5361 = ~STATE_REG_SCAN_IN | ~n6868;
  assign n5360 = ~DATAI_15_ | ~U3149;
  assign U3337 = ~n5361 | ~n5360;
  assign n5363 = ~STATE_REG_SCAN_IN | ~n5902;
  assign n5362 = ~DATAI_8_ | ~U3149;
  assign U3344 = ~n5363 | ~n5362;
  assign n5365 = ~STATE_REG_SCAN_IN | ~n6314;
  assign n5364 = ~DATAI_11_ | ~U3149;
  assign U3341 = ~n5365 | ~n5364;
  assign n5367 = ~n7622 | ~STATE_REG_SCAN_IN;
  assign n5366 = ~DATAI_18_ | ~U3149;
  assign U3334 = ~n5367 | ~n5366;
  assign n5369 = ~STATE_REG_SCAN_IN | ~n6091;
  assign n5368 = ~DATAI_9_ | ~U3149;
  assign U3343 = ~n5369 | ~n5368;
  assign n5371 = ~STATE_REG_SCAN_IN | ~n7387;
  assign n5370 = ~DATAI_16_ | ~U3149;
  assign U3336 = ~n5371 | ~n5370;
  assign n5373 = ~STATE_REG_SCAN_IN | ~n6357;
  assign n5372 = ~DATAI_12_ | ~U3149;
  assign U3340 = ~n5373 | ~n5372;
  assign n5375 = ~STATE_REG_SCAN_IN | ~n7463;
  assign n5374 = ~DATAI_17_ | ~U3149;
  assign U3335 = ~n5375 | ~n5374;
  assign n5377 = ~STATE_REG_SCAN_IN | ~n6508;
  assign n5376 = ~DATAI_13_ | ~U3149;
  assign U3339 = ~n5377 | ~n5376;
  assign n5378 = ~DATAI_23_ | ~U3149;
  assign U3329 = ~n7236 | ~n5378;
  assign n5380 = ~n7636 | ~STATE_REG_SCAN_IN;
  assign n5379 = ~DATAI_19_ | ~U3149;
  assign U3333 = ~n5380 | ~n5379;
  assign n5382 = ~n5381 | ~STATE_REG_SCAN_IN;
  assign n5384 = ~n5383 & ~n5382;
  assign n5386 = ~n5384 | ~IR_REG_31__SCAN_IN;
  assign n5385 = ~DATAI_31_ | ~U3149;
  assign U3321 = ~n5386 | ~n5385;
  assign n5389 = ~n5387;
  assign n5399 = ~n5389 & ~n5388;
  assign n5394 = ~D_REG_0__SCAN_IN & ~n5399;
  assign n5391 = ~n5390 | ~n5395;
  assign n5393 = ~n5392 & ~n5391;
  assign U3458 = ~n5394 & ~n5393;
  assign n5398 = ~D_REG_1__SCAN_IN & ~n5399;
  assign n5397 = n5396 & n5395;
  assign U3459 = ~n5398 & ~n5397;
  assign U3299 = D_REG_23__SCAN_IN & n5400;
  assign U3297 = D_REG_25__SCAN_IN & n5400;
  assign U3298 = D_REG_24__SCAN_IN & n5400;
  assign U3320 = D_REG_2__SCAN_IN & n5400;
  assign U3300 = D_REG_22__SCAN_IN & n5400;
  assign U3318 = D_REG_4__SCAN_IN & n5400;
  assign U3317 = D_REG_5__SCAN_IN & n5400;
  assign U3316 = D_REG_6__SCAN_IN & n5400;
  assign U3315 = D_REG_7__SCAN_IN & n5400;
  assign U3314 = D_REG_8__SCAN_IN & n5400;
  assign U3319 = D_REG_3__SCAN_IN & n5400;
  assign U3307 = D_REG_15__SCAN_IN & n5400;
  assign U3306 = D_REG_16__SCAN_IN & n5400;
  assign U3305 = D_REG_17__SCAN_IN & n5400;
  assign U3304 = D_REG_18__SCAN_IN & n5400;
  assign U3303 = D_REG_19__SCAN_IN & n5400;
  assign U3302 = D_REG_20__SCAN_IN & n5400;
  assign U3301 = D_REG_21__SCAN_IN & n5400;
  assign U3308 = D_REG_14__SCAN_IN & n5400;
  assign U3313 = D_REG_9__SCAN_IN & n5400;
  assign U3312 = D_REG_10__SCAN_IN & n5400;
  assign U3311 = D_REG_11__SCAN_IN & n5400;
  assign U3310 = D_REG_12__SCAN_IN & n5400;
  assign U3309 = D_REG_13__SCAN_IN & n5400;
  assign U3292 = D_REG_30__SCAN_IN & n5400;
  assign U3296 = D_REG_26__SCAN_IN & n5400;
  assign U3293 = D_REG_29__SCAN_IN & n5400;
  assign U3291 = D_REG_31__SCAN_IN & n5400;
  assign U3295 = D_REG_27__SCAN_IN & n5400;
  assign U3294 = D_REG_28__SCAN_IN & n5400;
  assign n7181 = n5662 & n5658;
  assign n6987 = ~n7181 & ~n7177;
  assign n5403 = ~n5402 | ~n5401;
  assign n5408 = ~n6987 & ~n5403;
  assign n5476 = ~n5924 | ~n7503;
  assign n5404 = ~n5474 | ~n7485;
  assign n5405 = ~n7725 | ~n5404;
  assign n5406 = ~n5535 | ~n5405;
  assign n5407 = ~n5476 | ~n5406;
  assign n5410 = ~n5408 & ~n5407;
  assign n5409 = ~REG3_REG_0__SCAN_IN | ~n7668;
  assign n5411 = ~n5410 | ~n5409;
  assign n5413 = ~n7743 | ~n5411;
  assign n5412 = ~n7832 | ~REG2_REG_0__SCAN_IN;
  assign U3290 = ~n5413 | ~n5412;
  assign n5415 = ~n6193 | ~DATAO_REG_10__SCAN_IN;
  assign n5414 = ~n6422 | ~U4043;
  assign U3560 = ~n5415 | ~n5414;
  assign n5417 = ~n6193 | ~DATAO_REG_11__SCAN_IN;
  assign n5416 = ~n6467 | ~U4043;
  assign U3561 = ~n5417 | ~n5416;
  assign n5419 = ~n6193 | ~DATAO_REG_15__SCAN_IN;
  assign n5418 = ~n6706 | ~U4043;
  assign U3565 = ~n5419 | ~n5418;
  assign n5421 = ~n6193 | ~DATAO_REG_14__SCAN_IN;
  assign n5420 = ~n6627 | ~U4043;
  assign U3564 = ~n5421 | ~n5420;
  assign n5423 = ~n6193 | ~DATAO_REG_13__SCAN_IN;
  assign n5422 = ~n6407 | ~U4043;
  assign U3563 = ~n5423 | ~n5422;
  assign n5425 = ~n6193 | ~DATAO_REG_12__SCAN_IN;
  assign n5424 = ~n6543 | ~U4043;
  assign U3562 = ~n5425 | ~n5424;
  assign n5432 = ~n6193 | ~DATAO_REG_31__SCAN_IN;
  assign n5427 = ~n5436 | ~REG0_REG_31__SCAN_IN;
  assign n5426 = ~n6130 | ~REG2_REG_31__SCAN_IN;
  assign n5430 = ~n5427 | ~n5426;
  assign n5428 = ~REG1_REG_31__SCAN_IN;
  assign n5429 = ~n6125 & ~n5428;
  assign n6992 = ~n7504;
  assign n5431 = ~n6992 | ~U4043;
  assign U3581 = ~n5432 | ~n5431;
  assign n5440 = ~n6193 | ~DATAO_REG_30__SCAN_IN;
  assign n5435 = n6130 & REG2_REG_30__SCAN_IN;
  assign n5433 = ~REG1_REG_30__SCAN_IN;
  assign n5434 = ~n6125 & ~n5433;
  assign n5438 = ~n5435 & ~n5434;
  assign n5437 = ~n5436 | ~REG0_REG_30__SCAN_IN;
  assign n5439 = ~n6990 | ~U4043;
  assign U3580 = ~n5440 | ~n5439;
  assign n5442 = ~n6193 | ~DATAO_REG_18__SCAN_IN;
  assign n5441 = ~n6654 | ~U4043;
  assign U3568 = ~n5442 | ~n5441;
  assign n5444 = ~n6193 | ~DATAO_REG_17__SCAN_IN;
  assign n5443 = ~n6832 | ~U4043;
  assign U3567 = ~n5444 | ~n5443;
  assign n5446 = ~n6193 | ~DATAO_REG_16__SCAN_IN;
  assign n5445 = ~n6928 | ~U4043;
  assign U3566 = ~n5446 | ~n5445;
  assign n5448 = ~n5991 | ~U4043;
  assign n5447 = ~n6193 | ~DATAO_REG_4__SCAN_IN;
  assign U3554 = ~n5448 | ~n5447;
  assign n5450 = ~n6341 | ~U4043;
  assign n5449 = ~n6193 | ~DATAO_REG_9__SCAN_IN;
  assign U3559 = ~n5450 | ~n5449;
  assign n5452 = ~n6022 | ~U4043;
  assign n5451 = ~n6193 | ~DATAO_REG_5__SCAN_IN;
  assign U3555 = ~n5452 | ~n5451;
  assign n5454 = ~n5927 | ~U4043;
  assign n5453 = ~n6193 | ~DATAO_REG_3__SCAN_IN;
  assign U3553 = ~n5454 | ~n5453;
  assign n5456 = ~n5794 | ~U4043;
  assign n5455 = ~n6193 | ~DATAO_REG_2__SCAN_IN;
  assign U3552 = ~n5456 | ~n5455;
  assign n5458 = ~n5924 | ~U4043;
  assign n5457 = ~n6193 | ~DATAO_REG_1__SCAN_IN;
  assign U3551 = ~n5458 | ~n5457;
  assign n5460 = ~n5662 | ~U4043;
  assign n5459 = ~n6193 | ~DATAO_REG_0__SCAN_IN;
  assign U3550 = ~n5460 | ~n5459;
  assign n5462 = ~n6261 | ~U4043;
  assign n5461 = ~n6193 | ~DATAO_REG_8__SCAN_IN;
  assign U3558 = ~n5462 | ~n5461;
  assign n5464 = ~n5879 | ~U4043;
  assign n5463 = ~n6193 | ~DATAO_REG_6__SCAN_IN;
  assign U3556 = ~n5464 | ~n5463;
  assign n5482 = ~n5470 & ~n5469;
  assign n5480 = ~REG1_REG_0__SCAN_IN | ~n7769;
  assign n5472 = ~n7740 & ~n7636;
  assign n7755 = ~n5472 & ~n7312;
  assign n5473 = ~n6878 & ~n7647;
  assign n5478 = ~n6987 & ~n5473;
  assign n5475 = ~n5535 | ~n5474;
  assign n5477 = ~n5476 | ~n5475;
  assign n5483 = n5478 | n5477;
  assign n5479 = ~n7767 | ~n5483;
  assign U3518 = ~n5480 | ~n5479;
  assign n5485 = ~REG0_REG_0__SCAN_IN | ~n7764;
  assign n5484 = ~n7763 | ~n5483;
  assign U3467 = ~n5485 | ~n5484;
  assign n5487 = ~n6193 | ~DATAO_REG_19__SCAN_IN;
  assign n5486 = ~n6834 | ~U4043;
  assign U3569 = ~n5487 | ~n5486;
  assign n5489 = ~n6193 | ~DATAO_REG_20__SCAN_IN;
  assign n5488 = ~n7411 | ~U4043;
  assign U3570 = ~n5489 | ~n5488;
  assign n5491 = ~n6193 | ~DATAO_REG_21__SCAN_IN;
  assign n5490 = ~n7268 | ~U4043;
  assign U3571 = ~n5491 | ~n5490;
  assign n5493 = ~n6196 | ~U4043;
  assign n5492 = ~n6193 | ~DATAO_REG_7__SCAN_IN;
  assign U3557 = ~n5493 | ~n5492;
  assign n5564 = ~n5563 | ~n5562;
  assign n5509 = ~n5504 & ~n5503;
  assign n5768 = ~n5504 | ~n5503;
  assign n5507 = ~n5529;
  assign n5511 = ~n7501;
  assign n5508 = ~n5768 | ~n7392;
  assign n5528 = ~n5509 & ~n5508;
  assign n6064 = ~STATE_REG_SCAN_IN & ~n5510;
  assign n7235 = ~n5583 & ~n5511;
  assign n5512 = ~n7235;
  assign n5522 = ~n5779 & ~n5778;
  assign n5523 = ~n5522 ^ n5777;
  assign n5524 = ~n7620 & ~n5523;
  assign n5526 = ~n6064 & ~n5524;
  assign n5525 = ~n7631 | ~ADDR_REG_7__SCAN_IN;
  assign n5527 = ~n5526 | ~n5525;
  assign n5531 = ~n5528 & ~n5527;
  assign n7637 = ~n5529 & ~n5581;
  assign n5530 = ~n7637 | ~n5767;
  assign U3247 = ~n5531 | ~n5530;
  assign n5651 = ~STATE_REG_SCAN_IN | ~n5532;
  assign n5541 = ~REG3_REG_0__SCAN_IN | ~n5651;
  assign n5576 = n5534 ^ n5533;
  assign n5539 = ~n5576 & ~n7813;
  assign n5537 = ~n7700 | ~n5535;
  assign n5536 = ~n7532 | ~n5924;
  assign n5538 = ~n5537 | ~n5536;
  assign n5540 = ~n5539 & ~n5538;
  assign U3229 = ~n5541 | ~n5540;
  assign n5544 = ~n7383 | ~n4567;
  assign n5542 = n7392 & n4579;
  assign n5543 = ~n5542 & ~n7637;
  assign n5545 = n5544 & n5543;
  assign n5552 = ~n5545 & ~n4607;
  assign n5550 = ~ADDR_REG_0__SCAN_IN | ~n7631;
  assign n5547 = ~n7392 | ~REG1_REG_0__SCAN_IN;
  assign n5546 = ~n7383 | ~REG2_REG_0__SCAN_IN;
  assign n5548 = ~n5547 | ~n5546;
  assign n5549 = ~n5548 | ~n4607;
  assign n5551 = ~n5550 | ~n5549;
  assign n5554 = ~n5552 & ~n5551;
  assign n5553 = ~REG3_REG_0__SCAN_IN | ~U3149;
  assign U3240 = ~n5554 | ~n5553;
  assign n5556 = ~n6193 | ~DATAO_REG_22__SCAN_IN;
  assign n5555 = ~n6937 | ~U4043;
  assign U3572 = ~n5556 | ~n5555;
  assign n5561 = ~n5558 & ~n5557;
  assign n5560 = ~n7383 | ~n5559;
  assign n5575 = ~n5561 & ~n5560;
  assign n5566 = ~n5563 & ~n5562;
  assign n5565 = ~n5564 | ~n7392;
  assign n5570 = ~n5566 & ~n5565;
  assign n5568 = ~ADDR_REG_2__SCAN_IN | ~n7631;
  assign n5567 = ~REG3_REG_2__SCAN_IN | ~U3149;
  assign n5569 = ~n5568 | ~n5567;
  assign n5573 = ~n5570 & ~n5569;
  assign n5572 = ~n7637 | ~n5571;
  assign n5574 = ~n5573 | ~n5572;
  assign n5588 = ~n5575 & ~n5574;
  assign n5580 = n5576 | n7501;
  assign n5577 = ~IR_REG_0__SCAN_IN & ~REG2_REG_0__SCAN_IN;
  assign n5578 = ~n5577 & ~n5623;
  assign n5579 = ~n7501 | ~n5578;
  assign n5582 = ~n5580 | ~n5579;
  assign n5585 = ~n5582 | ~n5581;
  assign n5584 = ~n5583 | ~IR_REG_0__SCAN_IN;
  assign n5587 = ~n5585 | ~n5584;
  assign n5605 = ~n5587 | ~U4043;
  assign U3242 = ~n5588 | ~n5605;
  assign n5592 = ~n5589 & ~REG1_REG_4__SCAN_IN;
  assign n5591 = ~n5590 | ~n7392;
  assign n5604 = ~n5592 & ~n5591;
  assign n5596 = ~n5593 & ~REG2_REG_4__SCAN_IN;
  assign n5595 = ~n7383 | ~n5594;
  assign n5599 = ~n5596 & ~n5595;
  assign n5834 = ~REG3_REG_4__SCAN_IN | ~U3149;
  assign n5597 = ~n7631 | ~ADDR_REG_4__SCAN_IN;
  assign n5598 = ~n5834 | ~n5597;
  assign n5602 = ~n5599 & ~n5598;
  assign n5601 = ~n7637 | ~n5600;
  assign n5603 = ~n5602 | ~n5601;
  assign n5606 = ~n5604 & ~n5603;
  assign U3244 = ~n5606 | ~n5605;
  assign n5608 = ~n7790 | ~n5924;
  assign n5607 = ~n7532 | ~n5927;
  assign n5612 = ~n5608 | ~n5607;
  assign n5610 = ~REG3_REG_2__SCAN_IN | ~n5651;
  assign n5609 = ~n7700 | ~n5937;
  assign n5611 = ~n5610 | ~n5609;
  assign n5619 = ~n5612 & ~n5611;
  assign n5615 = ~n5614 & ~n5613;
  assign n5616 = ~n5615 & ~n7813;
  assign n5618 = ~n5617 | ~n5616;
  assign U3234 = ~n5619 | ~n5618;
  assign n5621 = ~ADDR_REG_1__SCAN_IN | ~n7631;
  assign n5620 = ~REG3_REG_1__SCAN_IN | ~U3149;
  assign n5631 = ~n5621 | ~n5620;
  assign n5629 = ~n7637 | ~n5622;
  assign n5625 = ~n5624 & ~n5623;
  assign n5627 = ~n5625 & ~n7620;
  assign n5628 = ~n5627 | ~n5626;
  assign n5630 = ~n5629 | ~n5628;
  assign n5638 = ~n5631 & ~n5630;
  assign n5634 = ~n5633 & ~n5632;
  assign n5636 = ~n7628 & ~n5634;
  assign n5637 = ~n5636 | ~n5635;
  assign U3241 = ~n5638 | ~n5637;
  assign n5642 = ~n5640 ^ n5639;
  assign n5643 = ~n5642 ^ n5641;
  assign n5650 = ~n5643 & ~n7813;
  assign n5644 = ~n5662;
  assign n5646 = ~n7697 & ~n5644;
  assign n5645 = ~n5749 & ~n7788;
  assign n5648 = ~n5646 & ~n5645;
  assign n5647 = ~n7700 | ~n5663;
  assign n5649 = ~n5648 | ~n5647;
  assign n5653 = ~n5650 & ~n5649;
  assign n5652 = ~REG3_REG_1__SCAN_IN | ~n5651;
  assign U3219 = ~n5653 | ~n5652;
  assign n5655 = ~n6193 | ~DATAO_REG_23__SCAN_IN;
  assign n5654 = ~n7527 | ~U4043;
  assign U3573 = ~n5655 | ~n5654;
  assign n5683 = n7038 ^ n5656;
  assign n5661 = ~n5683 | ~n6779;
  assign n5659 = n5663 ^ n5658;
  assign n5682 = ~n5659 & ~n7757;
  assign n5660 = ~n5682 | ~n7485;
  assign n5675 = ~n5661 | ~n5660;
  assign n5665 = ~n5662 | ~n7722;
  assign n5664 = ~n5663 | ~n7650;
  assign n5672 = ~n5665 | ~n5664;
  assign n5667 = n7038 | n7177;
  assign n5668 = ~n5667 | ~n5666;
  assign n5670 = ~n5668 | ~n7647;
  assign n5669 = ~n5794 | ~n7503;
  assign n5671 = ~n5670 | ~n5669;
  assign n5674 = ~n5672 & ~n5671;
  assign n5673 = ~n5683 | ~n5472;
  assign n5681 = ~n5674 | ~n5673;
  assign n5676 = ~n5675 & ~n5681;
  assign n5678 = ~n5676 | ~n7743;
  assign n5677 = REG2_REG_1__SCAN_IN | n7743;
  assign n5680 = ~n5678 | ~n5677;
  assign n5679 = ~REG3_REG_1__SCAN_IN | ~n7668;
  assign U3289 = ~n5680 | ~n5679;
  assign n5687 = ~REG0_REG_1__SCAN_IN | ~n7764;
  assign n5685 = ~n5682 & ~n5681;
  assign n5684 = ~n5683 | ~n7312;
  assign n5688 = ~n5685 | ~n5684;
  assign n5686 = ~n7763 | ~n5688;
  assign U3469 = ~n5687 | ~n5686;
  assign n5690 = ~REG1_REG_1__SCAN_IN | ~n7769;
  assign n5689 = ~n7767 | ~n5688;
  assign U3519 = ~n5690 | ~n5689;
  assign n6023 = ~REG3_REG_6__SCAN_IN | ~U3149;
  assign n5691 = ~n7631 | ~ADDR_REG_6__SCAN_IN;
  assign n5703 = ~n6023 | ~n5691;
  assign n5693 = ~REG1_REG_6__SCAN_IN & ~n5692;
  assign n5695 = ~n5693 & ~n7628;
  assign n5701 = ~n5695 | ~n5694;
  assign n5697 = ~REG2_REG_6__SCAN_IN & ~n5696;
  assign n5699 = ~n5697 & ~n7620;
  assign n5700 = ~n5699 | ~n5698;
  assign n5702 = ~n5701 | ~n5700;
  assign n5706 = ~n5703 & ~n5702;
  assign n5705 = ~n7637 | ~n5704;
  assign U3246 = ~n5706 | ~n5705;
  assign n5992 = ~REG3_REG_5__SCAN_IN | ~U3149;
  assign n5707 = ~n7631 | ~ADDR_REG_5__SCAN_IN;
  assign n5721 = ~n5992 | ~n5707;
  assign n5710 = ~n5709 & ~n5708;
  assign n5712 = ~n5710 & ~n7628;
  assign n5719 = ~n5712 | ~n5711;
  assign n5715 = ~n5714 & ~n5713;
  assign n5717 = ~n5715 & ~n7620;
  assign n5718 = ~n5717 | ~n5716;
  assign n5720 = ~n5719 | ~n5718;
  assign n5724 = ~n5721 & ~n5720;
  assign n5723 = ~n7637 | ~n5722;
  assign U3245 = ~n5724 | ~n5723;
  assign n5795 = ~REG3_REG_3__SCAN_IN | ~U3149;
  assign n5725 = ~n7631 | ~ADDR_REG_3__SCAN_IN;
  assign n5734 = ~n5795 | ~n5725;
  assign n5732 = ~n7637 | ~n5726;
  assign n5728 = ~REG1_REG_3__SCAN_IN & ~n5727;
  assign n5730 = ~n5728 & ~n7628;
  assign n5731 = ~n5730 | ~n5729;
  assign n5733 = ~n5732 | ~n5731;
  assign n5740 = ~n5734 & ~n5733;
  assign n5736 = ~REG2_REG_3__SCAN_IN & ~n5735;
  assign n5738 = ~n5736 & ~n7620;
  assign n5739 = ~n5738 | ~n5737;
  assign U3243 = ~n5740 | ~n5739;
  assign n5746 = ~n7746 & ~REG3_REG_3__SCAN_IN;
  assign n5744 = ~REG2_REG_3__SCAN_IN | ~n7832;
  assign n5801 = n5742 ^ n5741;
  assign n5743 = ~n5801 | ~n7496;
  assign n5765 = ~n5746 & ~n5745;
  assign n5753 = ~n5801 | ~n5472;
  assign n5748 = ~n5991 | ~n7503;
  assign n5747 = ~n5789 | ~n7650;
  assign n5751 = ~n5748 | ~n5747;
  assign n5750 = ~n5749 & ~n7424;
  assign n5752 = ~n5751 & ~n5750;
  assign n5758 = ~n5753 | ~n5752;
  assign n5756 = ~n5755 ^ n5754;
  assign n5757 = ~n5756 & ~n7720;
  assign n5805 = ~n5758 & ~n5757;
  assign n5760 = ~n5940 & ~n5759;
  assign n5761 = ~n5760 & ~n7757;
  assign n5802 = n5761 & n5811;
  assign n5762 = ~n5802 | ~n7485;
  assign n5763 = ~n5805 | ~n5762;
  assign n5764 = ~n5763 | ~n7743;
  assign U3287 = ~n5765 | ~n5764;
  assign n6197 = ~REG3_REG_8__SCAN_IN | ~U3149;
  assign n5766 = ~n7631 | ~ADDR_REG_8__SCAN_IN;
  assign n5776 = ~n6197 | ~n5766;
  assign n5774 = ~n7637 | ~n5902;
  assign n5890 = ~n5769 | ~n5768;
  assign n5770 = ~REG1_REG_8__SCAN_IN & ~n5771;
  assign n5772 = ~n5770 & ~n7628;
  assign n5773 = ~n5772 | ~n5891;
  assign n5775 = ~n5774 | ~n5773;
  assign n5785 = ~n5776 & ~n5775;
  assign n5781 = ~REG2_REG_8__SCAN_IN & ~n5782;
  assign n5783 = ~n5781 & ~n7620;
  assign n5784 = ~n5783 | ~n5903;
  assign U3248 = ~n5785 | ~n5784;
  assign n5788 = n5787 ^ n5786;
  assign n5793 = ~n5788 & ~n7813;
  assign n5791 = ~n7700 | ~n5789;
  assign n5790 = ~n7532 | ~n5991;
  assign n5792 = ~n5791 | ~n5790;
  assign n5800 = ~n5793 & ~n5792;
  assign n5798 = ~REG3_REG_3__SCAN_IN & ~n7521;
  assign n5796 = ~n7790 | ~n5794;
  assign n5797 = ~n5796 | ~n5795;
  assign n5799 = ~n5798 & ~n5797;
  assign U3215 = ~n5800 | ~n5799;
  assign n5807 = ~REG1_REG_3__SCAN_IN | ~n7769;
  assign n5803 = n5801 & n7312;
  assign n5804 = ~n5803 & ~n5802;
  assign n5806 = ~n7767 | ~n5808;
  assign U3521 = ~n5807 | ~n5806;
  assign n5810 = ~REG0_REG_3__SCAN_IN | ~n7764;
  assign n5809 = ~n7763 | ~n5808;
  assign U3473 = ~n5810 | ~n5809;
  assign n5830 = ~REG1_REG_4__SCAN_IN | ~n7769;
  assign n5813 = ~n5876;
  assign n5812 = ~n5811 | ~n5816;
  assign n5857 = ~n5813 | ~n5812;
  assign n5824 = ~n5857 & ~n7757;
  assign n5815 = n5814 ^ n5825;
  assign n5823 = ~n5815 | ~n7647;
  assign n5818 = ~n6022 | ~n7503;
  assign n5817 = ~n5816 | ~n7650;
  assign n5821 = ~n5818 | ~n5817;
  assign n5820 = ~n5819 & ~n7424;
  assign n5822 = ~n5821 & ~n5820;
  assign n5828 = ~n5824 & ~n5854;
  assign n5864 = ~n5826 ^ n5825;
  assign n5827 = ~n5864 | ~n6878;
  assign n5829 = ~n7767 | ~n5831;
  assign U3522 = ~n5830 | ~n5829;
  assign n5833 = ~REG0_REG_4__SCAN_IN | ~n7764;
  assign n5832 = ~n7763 | ~n5831;
  assign U3475 = ~n5833 | ~n5832;
  assign n5838 = ~n7788 & ~n5965;
  assign n5836 = ~n5834;
  assign n5835 = ~n7521 & ~n5856;
  assign n5837 = n5836 | n5835;
  assign n5840 = ~n5838 & ~n5837;
  assign n5839 = ~n7790 | ~n5927;
  assign n5843 = ~n5840 | ~n5839;
  assign n5842 = ~n7793 & ~n5841;
  assign n5850 = ~n5843 & ~n5842;
  assign n5846 = ~n5845 & ~n5844;
  assign n5848 = ~n5846 & ~n7813;
  assign n5849 = ~n5848 | ~n5847;
  assign U3227 = ~n5850 | ~n5849;
  assign n5852 = ~n6193 | ~DATAO_REG_24__SCAN_IN;
  assign n5851 = ~n7560 | ~U4043;
  assign U3574 = ~n5852 | ~n5851;
  assign n5853 = n5864 & n5472;
  assign n5855 = ~n5854 & ~n5853;
  assign n5863 = ~n7832 & ~n5855;
  assign n5859 = ~n5856 & ~n7746;
  assign n7750 = ~n6819 | ~n7542;
  assign n5858 = ~n5857 & ~n7750;
  assign n5861 = ~n5859 & ~n5858;
  assign n5860 = ~n7832 | ~REG2_REG_4__SCAN_IN;
  assign n5862 = ~n5861 | ~n5860;
  assign n5866 = ~n5863 & ~n5862;
  assign n5865 = ~n5864 | ~n7496;
  assign U3286 = ~n5866 | ~n5865;
  assign n5868 = ~n7668 | ~n6006;
  assign n5867 = ~n7832 | ~REG2_REG_5__SCAN_IN;
  assign n5885 = ~n5868 | ~n5867;
  assign n5870 = ~n5869 ^ n6983;
  assign n5873 = ~n5871 & ~n7424;
  assign n5872 = ~n5994 & ~n7725;
  assign n5874 = ~n5873 & ~n5872;
  assign n5877 = ~n5876 & ~n5994;
  assign n5878 = ~n5877 & ~n7757;
  assign n5881 = ~n5878 | ~n5971;
  assign n5880 = ~n5879 | ~n7503;
  assign n5911 = ~n5881 | ~n5880;
  assign n5882 = n5911 & n7485;
  assign n5883 = ~n5912 & ~n5882;
  assign n5884 = ~n5883 & ~n7832;
  assign n5888 = ~n5885 & ~n5884;
  assign n5913 = n5886 ^ n6983;
  assign n5887 = ~n5913 | ~n6974;
  assign U3285 = ~n5888 | ~n5887;
  assign n6262 = ~REG3_REG_9__SCAN_IN | ~U3149;
  assign n5889 = ~n7631 | ~ADDR_REG_9__SCAN_IN;
  assign n5900 = ~n6262 | ~n5889;
  assign n5898 = ~n7637 | ~n6091;
  assign n5893 = ~n5894 & ~n5895;
  assign n5896 = ~n5893 & ~n7628;
  assign n6082 = ~n5895 | ~n5894;
  assign n5897 = ~n5896 | ~n6082;
  assign n5899 = ~n5898 | ~n5897;
  assign n5910 = ~n5900 & ~n5899;
  assign n5905 = ~n5906 & ~n5907;
  assign n5908 = ~n5905 & ~n7620;
  assign n5909 = ~n5908 | ~n6092;
  assign U3249 = ~n5910 | ~n5909;
  assign n5917 = ~REG0_REG_5__SCAN_IN | ~n7764;
  assign n5915 = ~n5912 & ~n5911;
  assign n5914 = ~n5913 | ~n6878;
  assign U3477 = ~n5917 | ~n5916;
  assign n5920 = ~REG1_REG_5__SCAN_IN | ~n7769;
  assign U3523 = ~n5920 | ~n5919;
  assign n5923 = n5921 | n7037;
  assign n5936 = ~n5950 | ~n5472;
  assign n5926 = ~n7650 | ~n5937;
  assign n5925 = ~n7722 | ~n5924;
  assign n5934 = ~n5926 | ~n5925;
  assign n5932 = ~n7503 | ~n5927;
  assign n5930 = ~n5929 ^ n5928;
  assign n5931 = ~n5930 | ~n7647;
  assign n5933 = ~n5932 | ~n5931;
  assign n5935 = ~n5934 & ~n5933;
  assign n5939 = ~n5938 | ~n5937;
  assign n5941 = ~n5939 | ~n7542;
  assign n5952 = n5941 | n5940;
  assign n5942 = ~n5952 & ~n7636;
  assign n5943 = ~n5954 & ~n5942;
  assign n5947 = ~n7832 & ~n5943;
  assign n5945 = ~REG3_REG_2__SCAN_IN | ~n7668;
  assign n5949 = ~n5947 & ~n5946;
  assign n5948 = ~n7832 | ~REG2_REG_2__SCAN_IN;
  assign U3288 = ~n5949 | ~n5948;
  assign n5956 = ~REG0_REG_2__SCAN_IN | ~n7764;
  assign n5951 = ~n5950 | ~n7312;
  assign n5953 = ~n5952 | ~n5951;
  assign n5957 = n5954 | n5953;
  assign n5955 = ~n7763 | ~n5957;
  assign U3471 = ~n5956 | ~n5955;
  assign n5959 = ~REG1_REG_2__SCAN_IN | ~n7769;
  assign n5958 = ~n7767 | ~n5957;
  assign U3520 = ~n5959 | ~n5958;
  assign n5970 = ~n5981 & ~n7740;
  assign n5964 = ~n6196 | ~n7503;
  assign n5963 = ~n6016 | ~n7650;
  assign n5967 = ~n5964 | ~n5963;
  assign n5966 = ~n5965 & ~n7424;
  assign n5968 = ~n5967 & ~n5966;
  assign n5977 = ~n5970 & ~n5982;
  assign n5972 = ~n5971 | ~n6016;
  assign n5973 = ~n5972 | ~n7542;
  assign n5984 = n5973 | n6030;
  assign n5975 = ~n5984 & ~n7636;
  assign n5974 = ~n7746 & ~n6021;
  assign n5976 = ~n5975 & ~n5974;
  assign n5980 = ~n7743 | ~n5978;
  assign n5979 = ~n7832 | ~REG2_REG_6__SCAN_IN;
  assign U3284 = ~n5980 | ~n5979;
  assign n5987 = ~REG1_REG_6__SCAN_IN | ~n7769;
  assign n5983 = ~n5981 & ~n7755;
  assign U3524 = ~n5987 | ~n5986;
  assign n5990 = ~REG0_REG_6__SCAN_IN | ~n7764;
  assign U3479 = ~n5990 | ~n5989;
  assign n5993 = ~n7790 | ~n5991;
  assign n6005 = ~n5993 | ~n5992;
  assign n5996 = ~n7793 & ~n5994;
  assign n5995 = ~n7788 & ~n6063;
  assign n6003 = ~n5996 & ~n5995;
  assign n5999 = ~n5998 & ~n5997;
  assign n6001 = ~n5999 & ~n7813;
  assign n6002 = ~n6001 | ~n6000;
  assign n6004 = ~n6003 | ~n6002;
  assign n6008 = ~n6005 & ~n6004;
  assign n6007 = ~n6006 | ~n7794;
  assign U3224 = ~n6008 | ~n6007;
  assign n6010 = ~n6193 | ~DATAO_REG_25__SCAN_IN;
  assign n6009 = ~n7533 | ~U4043;
  assign U3575 = ~n6010 | ~n6009;
  assign n6013 = ~n6012 ^ n6011;
  assign n6015 = ~n6014 ^ n6013;
  assign n6020 = ~n6015 & ~n7813;
  assign n6018 = ~n7700 | ~n6016;
  assign n6017 = ~n7532 | ~n6196;
  assign n6019 = ~n6018 | ~n6017;
  assign n6028 = ~n6020 & ~n6019;
  assign n6026 = ~n7521 & ~n6021;
  assign n6024 = ~n7790 | ~n6022;
  assign n6025 = ~n6024 | ~n6023;
  assign n6027 = ~n6026 & ~n6025;
  assign U3236 = ~n6028 | ~n6027;
  assign n6031 = n6030 | n6029;
  assign n6051 = ~n6031 | ~n6110;
  assign n6035 = ~n6051 & ~n7750;
  assign n6033 = n7746 | n6062;
  assign n6032 = ~n7832 | ~REG2_REG_7__SCAN_IN;
  assign n6034 = ~n6033 | ~n6032;
  assign n6050 = ~n6035 & ~n6034;
  assign n6046 = ~n6052 & ~n7661;
  assign n6044 = ~n6038 | ~n7647;
  assign n6040 = ~n6261 | ~n7503;
  assign n6039 = ~n6068 | ~n7650;
  assign n6042 = ~n6040 | ~n6039;
  assign n6041 = ~n6063 & ~n7424;
  assign n6043 = ~n6042 & ~n6041;
  assign n6048 = ~n7832 & ~n6056;
  assign n6047 = ~n6052 & ~n7667;
  assign n6049 = ~n6048 & ~n6047;
  assign U3283 = ~n6050 | ~n6049;
  assign n6058 = ~REG0_REG_7__SCAN_IN | ~n7764;
  assign n6054 = ~n6051 & ~n7757;
  assign n6053 = ~n6052 & ~n7678;
  assign n6055 = ~n6054 & ~n6053;
  assign U3481 = ~n6058 | ~n6057;
  assign n6061 = ~REG1_REG_7__SCAN_IN | ~n7769;
  assign U3525 = ~n6061 | ~n6060;
  assign n6072 = ~n6062 & ~n7521;
  assign n6065 = ~n7697 & ~n6063;
  assign n6067 = n6065 | n6064;
  assign n6066 = ~n7788 & ~n6162;
  assign n6070 = ~n6067 & ~n6066;
  assign n6069 = ~n7700 | ~n6068;
  assign n6071 = ~n6070 | ~n6069;
  assign n6078 = ~n6072 & ~n6071;
  assign n6075 = ~n6074 & ~n6073;
  assign n6076 = ~n6075 & ~n7813;
  assign U3210 = ~n6078 | ~n6077;
  assign n6080 = ~n6193 | ~DATAO_REG_26__SCAN_IN;
  assign n6079 = ~n7579 | ~U4043;
  assign U3576 = ~n6080 | ~n6079;
  assign n6342 = ~REG3_REG_10__SCAN_IN | ~U3149;
  assign n6081 = ~n7631 | ~ADDR_REG_10__SCAN_IN;
  assign n6090 = ~n6342 | ~n6081;
  assign n6088 = ~n7637 | ~n6151;
  assign n6139 = ~n6083 | ~n6082;
  assign n6084 = ~REG1_REG_10__SCAN_IN & ~n6085;
  assign n6086 = ~n6084 & ~n7628;
  assign n6140 = ~REG1_REG_10__SCAN_IN | ~n6085;
  assign n6089 = ~n6088 | ~n6087;
  assign n6098 = ~n6090 & ~n6089;
  assign n6094 = ~REG2_REG_10__SCAN_IN & ~n6095;
  assign n6096 = ~n6094 & ~n7620;
  assign n6097 = ~n6096 | ~n6152;
  assign U3250 = ~n6098 | ~n6097;
  assign n6100 = ~n6193 | ~DATAO_REG_27__SCAN_IN;
  assign n6099 = ~n7791 | ~U4043;
  assign U3577 = ~n6100 | ~n6099;
  assign n6118 = ~REG1_REG_8__SCAN_IN | ~n7769;
  assign n6103 = ~n6341 | ~n7503;
  assign n6106 = ~n6196 | ~n7722;
  assign n6105 = ~n6109 | ~n7650;
  assign n6107 = ~n6106 | ~n6105;
  assign n6111 = ~n6110 | ~n6109;
  assign n6112 = ~n6111 | ~n7542;
  assign n6253 = ~n6112 & ~n6172;
  assign n6115 = n6249 & n6878;
  assign U3526 = ~n6118 | ~n6117;
  assign n6121 = ~REG0_REG_8__SCAN_IN | ~n7764;
  assign U3483 = ~n6121 | ~n6120;
  assign n6137 = ~n6193 | ~DATAO_REG_29__SCAN_IN;
  assign n6124 = ~REG1_REG_29__SCAN_IN;
  assign n6129 = ~n6125 & ~n6124;
  assign n6126 = ~REG0_REG_29__SCAN_IN;
  assign n6128 = ~n6127 & ~n6126;
  assign n6132 = ~n6129 & ~n6128;
  assign n6131 = ~n6130 | ~REG2_REG_29__SCAN_IN;
  assign n6135 = ~n7789;
  assign n6136 = ~n6135 | ~U4043;
  assign U3579 = ~n6137 | ~n6136;
  assign n6138 = ~n7631 | ~ADDR_REG_11__SCAN_IN;
  assign n6149 = ~n6432 | ~n6138;
  assign n6147 = ~n7637 | ~n6314;
  assign n6143 = ~n6141 | ~n6140;
  assign n6142 = ~n6143 & ~n6144;
  assign n6145 = ~n6142 & ~n7628;
  assign n6305 = ~n6144 | ~n6143;
  assign n6159 = ~n6149 & ~n6148;
  assign n6154 = ~n6155 & ~n6156;
  assign n6157 = ~n6154 & ~n7620;
  assign U3251 = ~n6159 | ~n6158;
  assign n6178 = ~REG1_REG_9__SCAN_IN | ~n7769;
  assign n6170 = ~n7011 & ~n7148;
  assign n6167 = ~n6162 & ~n7424;
  assign n6165 = ~n7650 | ~n6163;
  assign n6164 = ~n7503 | ~n6422;
  assign n6166 = ~n6165 | ~n6164;
  assign n6168 = n6167 | n6166;
  assign n6173 = ~n6172 & ~n6264;
  assign n6174 = ~n6173 & ~n7757;
  assign U3527 = ~n6178 | ~n6177;
  assign n6181 = ~REG0_REG_9__SCAN_IN | ~n7764;
  assign U3485 = ~n6181 | ~n6180;
  assign n6190 = REG2_REG_9__SCAN_IN & n7832;
  assign n6183 = ~n6182 | ~n7485;
  assign n6186 = ~n6185 & ~n7740;
  assign n6191 = ~n7668 | ~n6276;
  assign U3281 = ~n6192 | ~n6191;
  assign n6195 = ~n6193 | ~DATAO_REG_28__SCAN_IN;
  assign n6194 = ~n7778 | ~U4043;
  assign U3578 = ~n6195 | ~n6194;
  assign n6198 = ~n7790 | ~n6196;
  assign n6213 = ~n6198 | ~n6197;
  assign n6201 = ~n7793 & ~n6199;
  assign n6200 = ~n7788 & ~n6224;
  assign n6211 = ~n6201 & ~n6200;
  assign n6209 = ~n6202;
  assign n6205 = ~n6204 & ~n6203;
  assign n6210 = n6209 | n6208;
  assign n6214 = ~n6250 | ~n7794;
  assign U3218 = ~n6215 | ~n6214;
  assign n6220 = ~n6340 & ~n7746;
  assign n6218 = ~n6238 | ~n7830;
  assign n6217 = ~n7832 | ~REG2_REG_10__SCAN_IN;
  assign n6219 = ~n6218 | ~n6217;
  assign n6236 = ~n6220 & ~n6219;
  assign n6228 = ~n6224 & ~n7424;
  assign n6226 = ~n7503 | ~n6467;
  assign n6225 = ~n7650 | ~n6335;
  assign n6227 = ~n6226 | ~n6225;
  assign n6229 = ~n6228 & ~n6227;
  assign U3280 = ~n6236 | ~n6235;
  assign n6244 = ~REG1_REG_10__SCAN_IN | ~n7769;
  assign n6239 = n6238 & n7542;
  assign U3528 = ~n6244 | ~n6243;
  assign n6247 = ~REG0_REG_10__SCAN_IN | ~n7764;
  assign U3487 = ~n6247 | ~n6246;
  assign n6248 = ~n7740;
  assign n6251 = ~n6250 | ~n7668;
  assign n6254 = n6253 & n7485;
  assign n6256 = ~n6255 & ~n6254;
  assign n6259 = ~REG2_REG_8__SCAN_IN | ~n7832;
  assign U3282 = ~n6260 | ~n6259;
  assign n6263 = ~n7790 | ~n6261;
  assign n6275 = ~n6263 | ~n6262;
  assign n6266 = ~n6290 & ~n7788;
  assign n6265 = ~n6264 & ~n7793;
  assign n6273 = ~n6266 & ~n6265;
  assign n6269 = ~n6268 & ~n6267;
  assign n6271 = ~n6269 & ~n7813;
  assign n6277 = ~n6276 | ~n7794;
  assign U3228 = ~n6278 | ~n6277;
  assign n6287 = ~n6421 & ~n7746;
  assign n6282 = ~n6281 & ~n6280;
  assign n6283 = ~n7757 & ~n6282;
  assign n6284 = ~n6324 | ~n7485;
  assign n6294 = ~n6290 & ~n7424;
  assign n6292 = ~n6436 | ~n7650;
  assign n6291 = ~n6543 | ~n7503;
  assign n6293 = ~n6292 | ~n6291;
  assign n6297 = ~n6294 & ~n6293;
  assign n6302 = ~n7832 | ~REG2_REG_11__SCAN_IN;
  assign U3279 = ~n6303 | ~n6302;
  assign n6469 = ~REG3_REG_12__SCAN_IN | ~U3149;
  assign n6304 = ~n7631 | ~ADDR_REG_12__SCAN_IN;
  assign n6313 = ~n6469 | ~n6304;
  assign n6311 = ~n7637 | ~n6357;
  assign n6356 = ~n6306 | ~n6305;
  assign n6358 = ~REG1_REG_12__SCAN_IN | ~n6308;
  assign n6348 = ~n6316 | ~n6315;
  assign n6317 = ~REG2_REG_12__SCAN_IN & ~n6318;
  assign n6319 = ~n6317 & ~n7620;
  assign U3252 = ~n6321 | ~n6320;
  assign n6328 = ~REG1_REG_11__SCAN_IN | ~n7769;
  assign U3529 = ~n6328 | ~n6327;
  assign n6331 = ~REG0_REG_11__SCAN_IN | ~n7764;
  assign U3489 = ~n6331 | ~n6330;
  assign n6337 = ~n7700 | ~n6335;
  assign n6336 = ~n6467 | ~n7532;
  assign n6338 = ~n6337 | ~n6336;
  assign n6345 = ~n7521 & ~n6340;
  assign n6343 = ~n7790 | ~n6341;
  assign n6344 = ~n6343 | ~n6342;
  assign n6346 = ~n6345 & ~n6344;
  assign U3214 = ~n6347 | ~n6346;
  assign n6351 = ~n6350 | ~n6349;
  assign n6509 = ~n6352 | ~n6351;
  assign n6541 = ~STATE_REG_SCAN_IN & ~n6355;
  assign n6360 = ~n6359 | ~n6358;
  assign n6499 = ~n6361 | ~n6360;
  assign n6365 = ~n7631 | ~ADDR_REG_13__SCAN_IN;
  assign n6369 = ~n7637 | ~n6508;
  assign U3253 = ~n6370 | ~n6369;
  assign n6389 = ~REG1_REG_12__SCAN_IN | ~n7769;
  assign n6375 = ~n6382 | ~n7650;
  assign n6374 = ~n6407 | ~n7503;
  assign n6376 = ~n6375 | ~n6374;
  assign n6531 = n6458 | n6385;
  assign U3530 = ~n6389 | ~n6388;
  assign n6392 = ~REG0_REG_12__SCAN_IN | ~n7764;
  assign U3491 = ~n6392 | ~n6391;
  assign n6394 = ~n6706 | ~n7503;
  assign n6393 = ~n6395 | ~n7650;
  assign n6485 = n6563 | n6398;
  assign n6399 = ~n6485 & ~n7636;
  assign n6412 = ~n6488 & ~n6399;
  assign n6401 = ~n6400;
  assign n6489 = ~n6403 | ~n6402;
  assign n6408 = ~n6407 | ~n7722;
  assign n6418 = ~n7746 & ~n6414;
  assign U3276 = ~n6420 | ~n6419;
  assign n6435 = ~n6439 & ~n7788;
  assign n6431 = ~n7521 & ~n6421;
  assign n6425 = ~n6424 & ~n6423;
  assign n6437 = ~n6436 | ~n7700;
  assign U3233 = ~n6438 | ~n6437;
  assign n6463 = ~REG1_REG_13__SCAN_IN | ~n7769;
  assign n6446 = ~n6457 | ~n7650;
  assign n6445 = ~n6627 | ~n7503;
  assign n6451 = ~n6450 | ~n6449;
  assign n6524 = ~n6452 | ~n6451;
  assign U3531 = ~n6463 | ~n6462;
  assign n6466 = ~REG0_REG_13__SCAN_IN | ~n7764;
  assign U3493 = ~n6466 | ~n6465;
  assign n6468 = ~n6467 | ~n7790;
  assign n6482 = ~n6469 | ~n6468;
  assign n6473 = ~n6470 & ~n7793;
  assign n6472 = ~n6471 & ~n7788;
  assign n6480 = ~n6473 & ~n6472;
  assign n6553 = ~n6476 & ~n6475;
  assign n6477 = ~n6476 | ~n6475;
  assign n6483 = ~n6528 | ~n7794;
  assign U3221 = ~n6484 | ~n6483;
  assign n6493 = ~REG0_REG_14__SCAN_IN | ~n7764;
  assign U3495 = ~n6493 | ~n6492;
  assign n6496 = ~REG1_REG_14__SCAN_IN | ~n7769;
  assign U3532 = ~n6496 | ~n6495;
  assign n6497 = ~n7631 | ~ADDR_REG_14__SCAN_IN;
  assign n6507 = ~n6498 | ~n6497;
  assign n6679 = ~n6500 | ~n6499;
  assign n6681 = ~REG1_REG_14__SCAN_IN | ~n6502;
  assign n6672 = ~n6510 | ~n6509;
  assign U3254 = ~n6515 | ~n6514;
  assign n6523 = ~n7746 & ~n6548;
  assign n6518 = ~n6517 & ~n7750;
  assign U3277 = ~n6526 | ~n6525;
  assign n6529 = ~n6528 | ~n7668;
  assign n6532 = ~n6531 & ~n7636;
  assign n6537 = ~REG2_REG_12__SCAN_IN | ~n7832;
  assign U3278 = ~n6538 | ~n6537;
  assign n6547 = ~n7793 & ~n6539;
  assign n6542 = ~n6540 & ~n7788;
  assign n6545 = ~n6542 & ~n6541;
  assign n6544 = ~n6543 | ~n7790;
  assign n6546 = ~n6545 | ~n6544;
  assign n6561 = ~n6547 & ~n6546;
  assign n6550 = ~n6549;
  assign n6556 = ~n6551 & ~n6550;
  assign U3231 = ~n6561 | ~n6560;
  assign n6567 = ~n7750 & ~n6587;
  assign n6565 = n7746 | n6625;
  assign n6564 = ~n7832 | ~REG2_REG_15__SCAN_IN;
  assign n6566 = ~n6565 | ~n6564;
  assign n6585 = ~n6567 & ~n6566;
  assign n6575 = ~n6621 | ~n7650;
  assign n6574 = ~n6928 | ~n7503;
  assign n6578 = ~n6627 | ~n7722;
  assign U3275 = ~n6585 | ~n6584;
  assign n6593 = ~REG0_REG_15__SCAN_IN | ~n7764;
  assign U3497 = ~n6593 | ~n6592;
  assign n6596 = ~REG1_REG_15__SCAN_IN | ~n7769;
  assign U3533 = ~n6596 | ~n6595;
  assign n6604 = ~n6705 & ~n7746;
  assign n6611 = ~n6607 & ~n7424;
  assign n6609 = ~n6700 | ~n7650;
  assign n6608 = ~n6832 | ~n7503;
  assign n6610 = ~n6609 | ~n6608;
  assign n6614 = ~n6611 & ~n6610;
  assign n6619 = ~n7832 | ~REG2_REG_16__SCAN_IN;
  assign U3274 = ~n6620 | ~n6619;
  assign n6623 = ~n7700 | ~n6621;
  assign n6622 = ~n6928 | ~n7532;
  assign n6631 = ~n6623 | ~n6622;
  assign n6626 = ~n6625 & ~n7521;
  assign n6629 = ~n6688 & ~n6626;
  assign n6628 = ~n6627 | ~n7790;
  assign n6630 = ~n6629 | ~n6628;
  assign n6636 = ~n6631 & ~n6630;
  assign U3238 = ~n6636 | ~n6635;
  assign n6643 = ~REG0_REG_16__SCAN_IN | ~n7764;
  assign U3499 = ~n6643 | ~n6642;
  assign n6646 = ~REG1_REG_16__SCAN_IN | ~n7769;
  assign U3534 = ~n6646 | ~n6645;
  assign n6668 = ~REG1_REG_17__SCAN_IN | ~n7769;
  assign n6849 = n6665 | n6664;
  assign U3535 = ~n6668 | ~n6667;
  assign n6671 = ~REG0_REG_17__SCAN_IN | ~n7764;
  assign U3501 = ~n6671 | ~n6670;
  assign n6675 = ~n6674 | ~n6673;
  assign n6869 = ~n6676 | ~n6675;
  assign n6683 = ~n6682 | ~n6681;
  assign n6859 = ~n6684 | ~n6683;
  assign n6693 = ~n7637 | ~n6868;
  assign U3255 = ~n6694 | ~n6693;
  assign n6697 = ~n6696 & ~n6695;
  assign n6702 = ~n7700 | ~n6700;
  assign n6701 = ~n6832 | ~n7532;
  assign n6703 = ~n6702 | ~n6701;
  assign n6709 = ~n7521 & ~n6705;
  assign n6707 = ~n6706 | ~n7790;
  assign n6858 = ~REG3_REG_16__SCAN_IN | ~U3149;
  assign n6708 = ~n6707 | ~n6858;
  assign n6710 = ~n6709 & ~n6708;
  assign U3223 = ~n6711 | ~n6710;
  assign n6715 = ~n6778 & ~n6788;
  assign n6741 = ~n6715 & ~n6714;
  assign n6717 = ~n6716;
  assign n6726 = ~n6915 & ~n7424;
  assign n6724 = ~n7411 | ~n7503;
  assign n6723 = ~n6722 | ~n7650;
  assign n6725 = ~n6724 | ~n6723;
  assign n6727 = ~n6726 & ~n6725;
  assign n6735 = ~n7764 | ~REG0_REG_19__SCAN_IN;
  assign U3505 = ~n6736 | ~n6735;
  assign n6738 = ~n7769 | ~REG1_REG_19__SCAN_IN;
  assign U3537 = ~n6739 | ~n6738;
  assign n6888 = ~n6743 & ~n6742;
  assign n6746 = n7286 | n6744;
  assign n6749 = ~n7268 | ~n7503;
  assign n6748 = ~n7273 | ~n7650;
  assign n6751 = ~n6749 | ~n6748;
  assign n6750 = ~n7267 & ~n7424;
  assign n6752 = ~n6751 & ~n6750;
  assign n6759 = ~n7764 | ~REG0_REG_20__SCAN_IN;
  assign U3506 = ~n6760 | ~n6759;
  assign n6762 = ~n7769 | ~REG1_REG_20__SCAN_IN;
  assign U3538 = ~n6763 | ~n6762;
  assign n6766 = n6764 | n7636;
  assign n6768 = ~n7668 | ~n6767;
  assign n6769 = ~n7743 | ~n6768;
  assign n6773 = n7743 | REG2_REG_19__SCAN_IN;
  assign n6776 = n6775 | n7667;
  assign U3271 = ~n6777 | ~n6776;
  assign n6796 = ~n6791 & ~n7424;
  assign n6794 = ~n6792 | ~n7650;
  assign n6793 = ~n6834 | ~n7503;
  assign n6795 = ~n6794 | ~n6793;
  assign n6804 = ~n7832 | ~REG2_REG_18__SCAN_IN;
  assign U3272 = ~n6805 | ~n6804;
  assign n6812 = ~REG1_REG_18__SCAN_IN | ~n7769;
  assign U3536 = ~n6812 | ~n6811;
  assign n6815 = ~REG0_REG_18__SCAN_IN | ~n7764;
  assign U3503 = ~n6815 | ~n6814;
  assign n6821 = n7746 | n7266;
  assign U3270 = ~n6827 | ~n6826;
  assign n6841 = ~n7521 & ~n6831;
  assign n6839 = ~n6832 | ~n7790;
  assign n6837 = ~n7793 & ~n6833;
  assign n6835 = ~n7532 | ~n6834;
  assign n7452 = ~U3149 | ~REG3_REG_18__SCAN_IN;
  assign n6836 = ~n6835 | ~n7452;
  assign n6838 = ~n6837 & ~n6836;
  assign n6840 = ~n6839 | ~n6838;
  assign n6842 = ~n6841 & ~n6840;
  assign U3235 = ~n6843 | ~n6842;
  assign n6855 = ~n7832 | ~REG2_REG_17__SCAN_IN;
  assign U3273 = ~n6856 | ~n6855;
  assign n6857 = ~n7631 | ~ADDR_REG_16__SCAN_IN;
  assign n7386 = ~n6860 | ~n6859;
  assign n7378 = ~n6870 | ~n6869;
  assign U3256 = ~n6875 | ~n6874;
  assign n6884 = ~n6881 | ~n6880;
  assign n6882 = ~n7769 | ~REG1_REG_22__SCAN_IN;
  assign U3540 = ~n6883 | ~n6882;
  assign n6885 = ~n7764 | ~REG0_REG_22__SCAN_IN;
  assign U3508 = ~n6886 | ~n6885;
  assign n6899 = ~n6895 & ~n7424;
  assign n6897 = ~n6937 | ~n7503;
  assign n6896 = ~n7417 | ~n7650;
  assign n6898 = ~n6897 | ~n6896;
  assign n6900 = ~n6899 & ~n6898;
  assign n6909 = ~n7764 | ~REG0_REG_21__SCAN_IN;
  assign U3507 = ~n6910 | ~n6909;
  assign n6912 = ~n7769 | ~REG1_REG_21__SCAN_IN;
  assign U3539 = ~n6913 | ~n6912;
  assign n6929 = ~n6928 | ~n7790;
  assign U3225 = ~n6930 | ~n6929;
  assign n7280 = ~n6932 | ~n7117;
  assign n6936 = ~n7336 & ~n7649;
  assign n6935 = ~n7305 & ~n7725;
  assign n6939 = ~n6936 & ~n6935;
  assign n6938 = ~n6937 | ~n7722;
  assign n6971 = ~n6941 & ~n6940;
  assign n6945 = ~n6942 | ~n7046;
  assign n7281 = ~n6945 | ~n6944;
  assign n6951 = ~n6971 | ~n6948;
  assign n6949 = ~n7764 | ~REG0_REG_23__SCAN_IN;
  assign U3509 = ~n6950 | ~n6949;
  assign n6952 = ~n7769 | ~REG1_REG_23__SCAN_IN;
  assign U3541 = ~n6953 | ~n6952;
  assign n6956 = ~n6955 & ~n6954;
  assign n6970 = ~n6958 | ~n6957;
  assign n6968 = ~n7521 & ~n6959;
  assign n6961 = ~n7790 | ~n7268;
  assign n6960 = ~U3149 | ~REG3_REG_22__SCAN_IN;
  assign n6963 = ~n6961 | ~n6960;
  assign n6962 = ~n7788 & ~n7282;
  assign n6966 = ~n6963 & ~n6962;
  assign n6965 = ~n7700 | ~n6964;
  assign n6967 = ~n6966 | ~n6965;
  assign n6969 = ~n6968 & ~n6967;
  assign U3232 = ~n6970 | ~n6969;
  assign n6972 = n7743 | REG2_REG_23__SCAN_IN;
  assign n6977 = ~n7746 & ~n7354;
  assign n6979 = n6978 | n6977;
  assign U3267 = ~n6982 | ~n6981;
  assign n6989 = ~n6984 & ~n6983;
  assign n7500 = ~n6985 | ~DATAI_30_;
  assign n7216 = ~n6990 & ~n7500;
  assign n6986 = ~DATAI_31_;
  assign n6991 = ~n6996 & ~n6986;
  assign n7221 = ~n7504 & ~n6991;
  assign n7099 = ~n7216 & ~n7221;
  assign n6988 = n6987 & n7099;
  assign n6998 = ~n6989 | ~n6988;
  assign n7724 = ~n6990;
  assign n7106 = ~n7724 & ~n7538;
  assign n6993 = ~n6992 & ~n7540;
  assign n7219 = ~n7106 & ~n6993;
  assign n6994 = ~DATAI_29_;
  assign n7748 = ~n6996 & ~n6994;
  assign n6995 = ~DATAI_28_;
  assign n7780 = ~n6996 & ~n6995;
  assign n7000 = ~n6999;
  assign n7137 = ~n7000 & ~n7148;
  assign n7002 = ~n7137 | ~n7121;
  assign n7027 = ~n7002 & ~n7001;
  assign n7006 = ~n7004 | ~n7003;
  assign n7023 = ~n7006 & ~n7005;
  assign n7194 = ~n7009 & ~n7008;
  assign n7012 = ~n7010;
  assign n7147 = ~n7012 & ~n7011;
  assign n7018 = ~n7194 | ~n7147;
  assign n7014 = ~n7196;
  assign n7016 = ~n7014 & ~n7013;
  assign n7017 = ~n7016 | ~n7015;
  assign n7019 = ~n7018 & ~n7017;
  assign n7021 = ~n7073 | ~n7019;
  assign n7022 = ~n7021 & ~n7020;
  assign n7025 = ~n7023 | ~n7022;
  assign n7026 = ~n7025 & ~n7024;
  assign n7028 = ~n7027 | ~n7026;
  assign n7572 = ~n7053 | ~n7093;
  assign n7331 = ~n7560 & ~n7522;
  assign n7321 = ~n7333 & ~n7331;
  assign n7438 = ~n7431 | ~n7055;
  assign n7033 = ~n7438 & ~n7280;
  assign n7035 = ~n7321 | ~n7033;
  assign n7049 = ~n7035 & ~n7034;
  assign n7039 = ~n7037 & ~n7036;
  assign n7040 = ~n7039 | ~n7038;
  assign n7042 = ~n7041 & ~n7040;
  assign n7044 = ~n7043 | ~n7042;
  assign n7047 = n7045 | n7044;
  assign n7048 = ~n7047 & ~n7046;
  assign n7075 = ~n7073 & ~n7072;
  assign n7076 = ~n7075 & ~n7074;
  assign n7098 = ~n7504 | ~n7538;
  assign n7107 = ~n7106 & ~n7504;
  assign n7109 = ~n7107 & ~n7540;
  assign n7110 = ~n7109 & ~n7108;
  assign n7118 = ~n7331 & ~n7117;
  assign n7210 = n7118 | n7430;
  assign n7127 = ~n7119 & ~n7123;
  assign n7122 = ~n7121 | ~n7120;
  assign n7165 = ~n7123 & ~n7122;
  assign n7128 = ~n7165 | ~n7124;
  assign n7126 = ~n7125 & ~n7128;
  assign n7157 = n7127 | n7126;
  assign n7129 = ~n7128;
  assign n7163 = ~n7130 | ~n7129;
  assign n7131 = n7158 | n7163;
  assign n7135 = ~n7132 & ~n7131;
  assign n7134 = ~n7133;
  assign n7142 = ~n7137 | ~n7136;
  assign n7202 = ~n7142 & ~n7139;
  assign n7141 = ~n7202;
  assign n7154 = ~n7141 & ~n7140;
  assign n7146 = ~n7142;
  assign n7145 = ~n7144 | ~n7143;
  assign n7152 = ~n7146 | ~n7145;
  assign n7150 = ~n7148 & ~n7147;
  assign n7151 = ~n7150 & ~n7149;
  assign n7153 = ~n7152 | ~n7151;
  assign n7155 = ~n7154 & ~n7153;
  assign n7156 = ~n7204 & ~n7155;
  assign n7172 = ~n7157 & ~n7156;
  assign n7160 = ~n7158;
  assign n7161 = ~n7160 | ~n7159;
  assign n7164 = n7162 & n7161;
  assign n7170 = ~n7164 & ~n7163;
  assign n7167 = ~n7166 | ~n7165;
  assign n7169 = ~n7168 | ~n7167;
  assign n7171 = ~n7170 & ~n7169;
  assign n7179 = ~n7177 & ~n7176;
  assign n7183 = ~n7179 & ~n7184;
  assign n7182 = ~n7181 & ~n7180;
  assign n7187 = ~n7183 | ~n7182;
  assign n7186 = ~n7178 | ~n7185;
  assign n7191 = ~n7187 | ~n7186;
  assign n7189 = ~n7194;
  assign n7190 = ~n7189 & ~n7188;
  assign n7200 = ~n7191 | ~n7190;
  assign n7195 = ~n7193 | ~n7192;
  assign n7197 = ~n7195 | ~n7194;
  assign n7198 = ~n7197 | ~n7196;
  assign n7199 = ~n7198 | ~n7178;
  assign n7206 = n7200 & n7199;
  assign n7203 = ~n7202 | ~n7201;
  assign n7205 = n7204 | n7203;
  assign n7222 = ~n7221;
  assign n7237 = ~n7235 | ~n7234;
  assign n7241 = ~n7237 | ~n7236;
  assign n7240 = ~n7239 | ~n7238;
  assign n7242 = ~n7241 | ~n7240;
  assign n7243 = ~n7242 | ~B_REG_SCAN_IN;
  assign U3239 = ~n7244 | ~n7243;
  assign n7247 = ~n7746 & ~n7410;
  assign n7248 = ~n7832 & ~n7247;
  assign U3269 = n7256 | n7255;
  assign n7260 = n7258 | n7257;
  assign n7263 = n7261 | n7403;
  assign n7279 = n7265 | n7404;
  assign n7277 = ~n7521 & ~n7266;
  assign n7272 = ~n7697 & ~n7267;
  assign n7270 = ~n7532 | ~n7268;
  assign n7269 = ~U3149 | ~REG3_REG_20__SCAN_IN;
  assign n7271 = ~n7270 | ~n7269;
  assign n7275 = ~n7272 & ~n7271;
  assign n7274 = ~n7700 | ~n7273;
  assign n7276 = ~n7275 | ~n7274;
  assign n7278 = ~n7277 & ~n7276;
  assign U3230 = ~n7279 | ~n7278;
  assign n7292 = ~n7322 & ~n7661;
  assign n7332 = ~n7290 | ~n7289;
  assign n7295 = ~n7527 | ~n7722;
  assign n7294 = ~n7308 | ~n7650;
  assign n7302 = ~n7322 | ~n5472;
  assign n7309 = ~n7306 | ~n7305;
  assign n7318 = n7493 | n7315;
  assign n7316 = ~n7769 | ~REG1_REG_24__SCAN_IN;
  assign U3542 = ~n7317 | ~n7316;
  assign n7319 = ~n7764 | ~REG0_REG_24__SCAN_IN;
  assign U3510 = ~n7320 | ~n7319;
  assign n7324 = ~n7322 & ~n7321;
  assign n7437 = ~n7324 & ~n7323;
  assign n7441 = ~n7327 | ~n7559;
  assign n7429 = ~n7332 & ~n7331;
  assign n7340 = ~n7579 | ~n7503;
  assign n7338 = ~n7336 & ~n7424;
  assign n7337 = ~n7559 & ~n7725;
  assign n7339 = ~n7338 & ~n7337;
  assign n7366 = ~n7342 & ~n7341;
  assign n7346 = ~n7343 | ~n7366;
  assign n7344 = ~n7764 | ~REG0_REG_25__SCAN_IN;
  assign U3511 = ~n7345 | ~n7344;
  assign n7347 = ~n7769 | ~REG1_REG_25__SCAN_IN;
  assign U3543 = ~n7348 | ~n7347;
  assign n7351 = ~n7350 & ~n7349;
  assign n7365 = ~n7353 | ~n7352;
  assign n7363 = ~n7521 & ~n7354;
  assign n7358 = ~n7697 & ~n7414;
  assign n7356 = ~n7532 | ~n7560;
  assign n7355 = ~U3149 | ~REG3_REG_23__SCAN_IN;
  assign n7357 = ~n7356 | ~n7355;
  assign n7361 = ~n7358 & ~n7357;
  assign n7360 = ~n7700 | ~n7359;
  assign n7362 = ~n7361 | ~n7360;
  assign n7364 = ~n7363 & ~n7362;
  assign U3213 = ~n7365 | ~n7364;
  assign n7373 = ~n7558 | ~n7668;
  assign n7372 = n7371 | n7750;
  assign U3265 = ~n7377 | ~n7376;
  assign n7390 = ~n7389 | ~n7388;
  assign n7453 = ~n7391 | ~n7390;
  assign n7401 = ~n7637 | ~n7463;
  assign U3257 = ~n7402 | ~n7401;
  assign n7421 = ~n7521 & ~n7410;
  assign n7413 = ~n7790 | ~n7411;
  assign n7412 = ~REG3_REG_21__SCAN_IN | ~U3149;
  assign n7416 = ~n7413 | ~n7412;
  assign n7415 = ~n7788 & ~n7414;
  assign n7419 = ~n7416 & ~n7415;
  assign n7418 = ~n7700 | ~n7417;
  assign n7420 = ~n7419 | ~n7418;
  assign n7422 = ~n7421 & ~n7420;
  assign U3220 = ~n7423 | ~n7422;
  assign n7426 = ~n7698 & ~n7424;
  assign n7425 = ~n7573 & ~n7725;
  assign n7427 = ~n7426 & ~n7425;
  assign n7584 = ~n7430 & ~n7429;
  assign n7472 = ~n7436 & ~n7435;
  assign n7440 = ~n7438 | ~n7437;
  assign n7507 = ~n7441 & ~n7699;
  assign n7448 = ~n7472 | ~n7445;
  assign n7446 = ~n7764 | ~REG0_REG_26__SCAN_IN;
  assign U3512 = ~n7447 | ~n7446;
  assign n7449 = ~n7769 | ~REG1_REG_26__SCAN_IN;
  assign U3544 = ~n7450 | ~n7449;
  assign n7451 = ~n7631 | ~ADDR_REG_18__SCAN_IN;
  assign n7456 = ~n7454 | ~n7453;
  assign U3258 = ~n7471 | ~n7470;
  assign n7480 = ~n7705 | ~n7668;
  assign n7479 = n7478 | n7750;
  assign U3264 = ~n7484 | ~n7483;
  assign n7487 = ~n7746 & ~n7520;
  assign n7488 = ~n7832 & ~n7487;
  assign n7494 = ~n7743 & ~REG2_REG_24__SCAN_IN;
  assign n7499 = n7495 | n7494;
  assign U3266 = ~n7499 | ~n7498;
  assign n7510 = ~REG0_REG_30__SCAN_IN | ~n7764;
  assign n7505 = ~n7500 & ~n7725;
  assign n7502 = ~n7501 | ~B_REG_SCAN_IN;
  assign n7723 = ~n7503 | ~n7502;
  assign n7536 = ~n7504 & ~n7723;
  assign n7669 = ~n7507 | ~n7506;
  assign n7749 = ~n7669 & ~n7780;
  assign n7539 = ~n7749 | ~n7726;
  assign U3516 = ~n7510 | ~n7509;
  assign n7513 = ~REG1_REG_30__SCAN_IN | ~n7769;
  assign U3548 = ~n7513 | ~n7512;
  assign n7516 = ~n7518 & ~n7517;
  assign n7553 = ~n7518 | ~n7517;
  assign n7524 = ~n7521 & ~n7520;
  assign n7523 = ~n7793 & ~n7522;
  assign n7529 = ~n7790 | ~n7527;
  assign n7528 = ~REG3_REG_24__SCAN_IN | ~U3149;
  assign n7534 = ~n7533 | ~n7532;
  assign U3226 = ~n7535 | ~n7534;
  assign n7545 = ~REG0_REG_31__SCAN_IN | ~n7764;
  assign n7537 = ~n7540 & ~n7725;
  assign n7541 = ~n7539 & ~n7538;
  assign U3517 = ~n7545 | ~n7544;
  assign n7548 = ~REG1_REG_31__SCAN_IN | ~n7769;
  assign U3549 = ~n7548 | ~n7547;
  assign n7568 = ~n7574 & ~n7788;
  assign n7566 = ~n7558 | ~n7794;
  assign n7564 = ~n7793 & ~n7559;
  assign n7562 = ~n7790 | ~n7560;
  assign n7561 = ~REG3_REG_25__SCAN_IN | ~U3149;
  assign n7563 = ~n7562 | ~n7561;
  assign n7565 = ~n7564 & ~n7563;
  assign n7567 = ~n7566 | ~n7565;
  assign n7569 = ~n7568 & ~n7567;
  assign U3222 = ~n7570 | ~n7569;
  assign n7588 = ~n7643 | ~n7644;
  assign n7576 = ~n7572 | ~n7571;
  assign n7577 = n7576 & n7575;
  assign n7578 = n7588 | n7577;
  assign n7659 = ~n7588 | ~n7577;
  assign n7605 = ~n7578 | ~n7659;
  assign n7580 = ~n7657 | ~n7650;
  assign n7591 = ~n7583 & ~n7582;
  assign n7642 = ~n7587 & ~n7586;
  assign n7610 = ~n7593 & ~n7592;
  assign n7594 = n7743 | REG2_REG_27__SCAN_IN;
  assign n7600 = ~n7596 & ~n7746;
  assign n7601 = n7600 | n7599;
  assign U3263 = ~n7604 | ~n7603;
  assign n7613 = ~n7610 | ~n7609;
  assign n7611 = ~n7764 | ~REG0_REG_27__SCAN_IN;
  assign U3513 = ~n7612 | ~n7611;
  assign n7614 = ~n7769 | ~REG1_REG_27__SCAN_IN;
  assign U3545 = ~n7615 | ~n7614;
  assign n7618 = ~n7636 ^ REG2_REG_19__SCAN_IN;
  assign n7638 = ~n7637 | ~n7636;
  assign U3259 = ~n7639 | ~n7638;
  assign n7712 = n7643 & n7642;
  assign n7654 = ~n7789 & ~n7649;
  assign n7652 = ~n7791 | ~n7722;
  assign n7651 = ~n7780 | ~n7650;
  assign n7684 = ~n7663 & ~n7662;
  assign n7672 = n7680 | n7750;
  assign U3262 = ~n7677 | ~n7676;
  assign n7687 = ~n7684 | ~n7683;
  assign n7685 = ~n7769 | ~REG1_REG_28__SCAN_IN;
  assign U3546 = ~n7686 | ~n7685;
  assign n7688 = ~n7764 | ~REG0_REG_28__SCAN_IN;
  assign U3514 = ~n7689 | ~n7688;
  assign n7709 = ~n7696 & ~n7788;
  assign n7704 = ~n7698 & ~n7697;
  assign n7702 = ~n7700 | ~n7699;
  assign n7701 = ~REG3_REG_26__SCAN_IN | ~U3149;
  assign n7703 = ~n7702 | ~n7701;
  assign n7707 = ~n7704 & ~n7703;
  assign n7706 = ~n7705 | ~n7794;
  assign n7708 = ~n7707 | ~n7706;
  assign n7710 = ~n7709 & ~n7708;
  assign U3237 = ~n7711 | ~n7710;
  assign n7719 = ~n7715 & ~n7714;
  assign n7728 = ~n7724 & ~n7723;
  assign n7727 = ~n7726 & ~n7725;
  assign n7729 = ~n7728 & ~n7727;
  assign n7762 = ~n7732 & ~n7731;
  assign n7737 = ~n7735 & ~n7734;
  assign n7738 = ~n7737 & ~n7736;
  assign n7756 = n7739 ^ n7738;
  assign n7741 = ~n7756 & ~n7740;
  assign n7742 = ~n7741 & ~n7832;
  assign n7745 = ~n7762 | ~n7742;
  assign n7744 = n7743 | REG2_REG_29__SCAN_IN;
  assign U3354 = ~n7754 | ~n7753;
  assign n7760 = ~n7756 & ~n7755;
  assign n7768 = ~n7762 | ~n7761;
  assign n7766 = ~n7768 | ~n7763;
  assign n7765 = ~n7764 | ~REG0_REG_29__SCAN_IN;
  assign U3515 = ~n7766 | ~n7765;
  assign n7771 = ~n7768 | ~n7767;
  assign n7770 = ~n7769 | ~REG1_REG_29__SCAN_IN;
  assign U3547 = ~n7771 | ~n7770;
  assign n7773 = ~n7780 | ~n7772;
  assign n7781 = ~n7780 | ~n7779;
  assign n7787 = ~n7812 & ~n7813;
  assign n7803 = ~n7789 & ~n7788;
  assign n7801 = ~n7791 | ~n7790;
  assign n7799 = ~n7793 & ~n7792;
  assign n7797 = ~U3149 | ~REG3_REG_28__SCAN_IN;
  assign n7796 = ~n7795 | ~n7794;
  assign n7798 = ~n7797 | ~n7796;
  assign n7800 = ~n7799 & ~n7798;
  assign n7802 = ~n7801 | ~n7800;
  assign n7804 = ~n7803 & ~n7802;
  assign n7822 = n7805 & n7804;
  assign n7809 = ~n7811 | ~n7808;
  assign n7820 = ~n7810 & ~n7809;
  assign n7816 = ~n7811;
  assign n7817 = ~n7816 | ~n7815;
  assign n7819 = ~n7818 & ~n7817;
  assign U3217 = ~n7822 | ~n7821;
  assign n7828 = ~n7832 & ~n7823;
  assign U3260 = n7828 | n7827;
  assign n7836 = ~n7832 & ~n7829;
  assign U3261 = n7836 | n7835;
endmodule


