// Benchmark "b17_C" written by ABC on Thu Mar  5 01:04:08 2020

module b17_C ( 
    P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
    DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
    DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
    DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
    DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
    DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
    P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
    P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
    P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
    P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
    P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
    P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
    P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
    P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
    P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
    P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
    P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
    P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
    P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
    P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
    P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
    P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
    P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
    P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
    P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
    P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
    P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
    P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
    P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
    P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
    P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
    P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
    P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
    P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
    P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
    P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
    P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
    P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
    P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
    P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
    P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
    P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
    P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
    P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
    P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
    P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
    P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
    P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN,
    P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN,
    P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN,
    P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN,
    P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN,
    P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN,
    P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN,
    P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN,
    P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN,
    P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN,
    P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN,
    P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN,
    P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN,
    P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN,
    P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN,
    P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN,
    P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN,
    P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN,
    P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN,
    P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN,
    P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN,
    P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN,
    P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN,
    P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN,
    P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN,
    P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN,
    P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN,
    P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN,
    P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN,
    P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN,
    P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN,
    P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN,
    P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN,
    P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN,
    P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN,
    P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN,
    P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN,
    P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN,
    P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN,
    P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN,
    P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN,
    P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN,
    P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN,
    P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN,
    P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN,
    P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN,
    P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN,
    P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN,
    P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN,
    P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN,
    P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN,
    P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN,
    P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN,
    P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN,
    P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN,
    P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN,
    P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN,
    P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN,
    P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN,
    P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN,
    P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN,
    P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN,
    BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN,
    BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN,
    BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN,
    BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN,
    BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN,
    BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN,
    BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN,
    BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN,
    BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN,
    BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN,
    BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN,
    BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN,
    BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN,
    BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN,
    BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN,
    BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN,
    BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN,
    BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN,
    BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN,
    BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN,
    BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN,
    READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN,
    P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN,
    P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN,
    P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN,
    P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN,
    P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN,
    P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN,
    P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN,
    P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN,
    P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN,
    P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN,
    P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN,
    P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN,
    P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN,
    P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN,
    P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN,
    P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN,
    P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN,
    P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN,
    P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN,
    P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN,
    P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN,
    P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN,
    P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN,
    P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN,
    P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN,
    P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN,
    P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN,
    P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN,
    P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN,
    P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN,
    P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN,
    P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN,
    P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN,
    P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN,
    P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN,
    P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN,
    P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN,
    P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN,
    P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN,
    P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN,
    P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN,
    P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN,
    P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN,
    P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN,
    P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN,
    P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN,
    P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN,
    P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN,
    P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN,
    P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN,
    P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN,
    P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN,
    P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN,
    P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN,
    P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN,
    P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN,
    P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN,
    P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN,
    P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN,
    P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN,
    P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN,
    P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN,
    P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN,
    P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN,
    P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN,
    P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN,
    P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN,
    P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN,
    P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN,
    P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN,
    P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN,
    P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN,
    P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN,
    P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN,
    P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN,
    P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN,
    P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN,
    P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN,
    P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN,
    P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN,
    P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN,
    P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN,
    P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN,
    P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN,
    P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN,
    P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN,
    P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN,
    P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN,
    P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN,
    P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN,
    P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN,
    P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN,
    P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN,
    P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN,
    P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN,
    P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN,
    P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN,
    P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN,
    P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN,
    P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
    P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
    P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
    P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
    P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
    P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
    P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN,
    P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN,
    P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN,
    P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN,
    P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN,
    P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN,
    P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN,
    P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN,
    P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN,
    P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN,
    P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
    P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
    P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
    P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
    P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
    P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
    P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
    P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
    P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
    P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
    P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
    P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
    P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
    P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
    P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
    P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
    P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
    P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
    P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
    P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
    P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
    P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
    P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
    P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
    P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
    P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
    P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
    P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
    P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
    P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
    P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
    P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
    P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
    P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
    P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
    P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN,
    P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
    P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN,
    P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
    P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN,
    P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
    P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
    P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
    P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
    P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
    P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN,
    P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
    P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN,
    P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
    P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN,
    P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
    P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN,
    P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
    P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN,
    P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
    P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
    P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
    P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
    P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
    P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
    P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
    P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
    P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
    P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
    P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
    P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
    P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
    P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
    P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
    P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
    P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
    P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
    P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
    P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
    P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN,
    P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN,
    P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN,
    P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN,
    P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN,
    P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN,
    P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN,
    P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN,
    P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN,
    P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN,
    P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN,
    P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN,
    P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN,
    P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN,
    P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN,
    P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN,
    P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN,
    P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN,
    P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN,
    P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN,
    P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN,
    P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN,
    P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN,
    P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN,
    P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN,
    P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN,
    P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN,
    P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN,
    P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN,
    P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN,
    P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN,
    P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN,
    P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN,
    P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN,
    P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN,
    P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN,
    P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN,
    P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN,
    P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN,
    P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN,
    P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN,
    P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN,
    P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN,
    P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN,
    P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN,
    P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN,
    P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN,
    P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN,
    P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN,
    P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN,
    P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN,
    P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN,
    P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN,
    P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN,
    P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN,
    P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN,
    P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN,
    P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN,
    P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN,
    P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN,
    P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN,
    P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN,
    P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN,
    P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN,
    P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN,
    P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN,
    P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN,
    P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN,
    P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN,
    P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN,
    P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN,
    P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN,
    P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN,
    P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN,
    P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN,
    P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN,
    P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN,
    P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN,
    P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN,
    P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN,
    P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN,
    P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN,
    P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN,
    P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN,
    P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN,
    P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN,
    P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN,
    P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN,
    P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN,
    P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN,
    P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN,
    P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN,
    P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN,
    P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN,
    P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN,
    P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN,
    P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN,
    P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN,
    P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN,
    P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
    P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
    P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
    P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
    P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
    P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN,
    P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN,
    P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN,
    P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN,
    P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN,
    P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN,
    P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN,
    P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN,
    P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN,
    P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN,
    P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
    P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
    P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
    P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
    P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
    P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
    P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
    P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
    P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
    P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
    P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
    P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
    P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
    P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
    P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
    P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
    P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
    P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
    P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
    P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
    P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
    P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
    P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
    P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
    P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
    P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
    P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
    P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
    P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
    P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
    P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
    P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
    P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
    P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
    P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
    P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
    P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
    P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
    P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
    P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
    P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
    P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
    P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN,
    P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN,
    P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN,
    P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN,
    P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN,
    P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN,
    P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN,
    P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN,
    P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN,
    P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN,
    P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN,
    P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN,
    P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN,
    P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN,
    P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN,
    P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN,
    P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN,
    P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN,
    P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN,
    P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN,
    P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN,
    P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN,
    P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN,
    P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN,
    P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN,
    P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN,
    P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN,
    P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN,
    P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN,
    P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN,
    P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN,
    P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN,
    P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN,
    P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN,
    P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN,
    P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN,
    P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN,
    P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN,
    P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN,
    P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN,
    P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN,
    P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN,
    P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN,
    P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN,
    P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN,
    P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN,
    P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN,
    P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN,
    P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN,
    P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN,
    P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN,
    P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN,
    P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN,
    P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN,
    P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN,
    P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN,
    P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN,
    P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN,
    P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN,
    P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN,
    P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN,
    P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN,
    P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN,
    P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN,
    P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN,
    P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN,
    P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN,
    P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN,
    P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN,
    P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN,
    P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN,
    P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN,
    P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN,
    P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN,
    P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN,
    P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN,
    P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN,
    P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN,
    P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN,
    P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN,
    P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN,
    P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN,
    U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367,
    U368, U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350,
    U351, U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242,
    U241, U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230,
    U229, U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218,
    U217, U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260,
    U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272,
    U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215,
    U213, U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060,
    P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053,
    P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046,
    P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039,
    P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032,
    P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027,
    P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020,
    P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013,
    P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006,
    P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999,
    P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993,
    P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986,
    P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979,
    P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972,
    P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965,
    P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958,
    P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951,
    P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944,
    P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937,
    P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930,
    P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923,
    P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916,
    P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909,
    P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902,
    P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895,
    P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888,
    P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881,
    P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874,
    P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284,
    P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865,
    P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858,
    P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851,
    P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844,
    P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837,
    P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830,
    P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823,
    P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816,
    P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809,
    P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802,
    P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795,
    P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788,
    P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781,
    P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774,
    P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767,
    P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760,
    P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753,
    P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746,
    P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739,
    P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732,
    P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725,
    P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718,
    P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711,
    P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704,
    P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697,
    P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690,
    P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683,
    P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676,
    P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669,
    P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662,
    P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655,
    P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648,
    P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641,
    P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637,
    P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633,
    P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213,
    P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208,
    P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201,
    P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194,
    P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187,
    P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180,
    P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174,
    P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167,
    P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160,
    P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153,
    P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146,
    P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139,
    P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132,
    P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125,
    P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118,
    P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111,
    P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104,
    P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097,
    P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090,
    P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083,
    P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076,
    P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069,
    P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062,
    P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055,
    P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048,
    P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602,
    P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043,
    P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036,
    P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029,
    P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022,
    P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015,
    P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008,
    P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001,
    P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994,
    P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987,
    P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980,
    P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973,
    P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966,
    P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959,
    P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952,
    P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945,
    P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938,
    P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931,
    P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924,
    P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917,
    P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910,
    P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903,
    P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896,
    P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889,
    P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882,
    P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875,
    P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868,
    P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861,
    P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854,
    P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847,
    P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840,
    P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833,
    P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826,
    P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608,
    P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816,
    P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461,
    P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220,
    P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213,
    P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206,
    P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199,
    P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465,
    P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187,
    P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180,
    P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173,
    P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166,
    P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160,
    P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153,
    P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146,
    P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139,
    P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132,
    P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125,
    P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118,
    P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111,
    P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104,
    P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097,
    P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090,
    P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083,
    P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076,
    P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069,
    P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062,
    P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055,
    P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048,
    P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041,
    P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034,
    P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032,
    P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029,
    P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022,
    P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015,
    P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008,
    P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001,
    P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994,
    P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987,
    P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980,
    P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973,
    P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966,
    P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959,
    P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952,
    P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945,
    P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938,
    P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931,
    P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924,
    P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917,
    P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910,
    P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903,
    P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896,
    P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889,
    P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882,
    P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875,
    P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868,
    P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861,
    P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854,
    P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847,
    P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840,
    P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833,
    P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826,
    P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819,
    P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812,
    P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482,
    P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486,
    P1_U2803, P1_U2802, P1_U3487, P1_U2801  );
  input  P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
    DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
    DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
    DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
    DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
    DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
    P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
    P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
    P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
    P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
    P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
    P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
    P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
    P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
    P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
    P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
    P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
    P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
    P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
    P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
    P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
    P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
    P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
    P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
    P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
    P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
    P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
    P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
    P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
    P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
    P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
    P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
    P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
    P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
    P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
    P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
    P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
    P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
    P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
    P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
    P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
    P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
    P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
    P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
    P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
    P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
    P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
    P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN,
    P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN,
    P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN,
    P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN,
    P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN,
    P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN,
    P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN,
    P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN,
    P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN,
    P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN,
    P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN,
    P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN,
    P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN,
    P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN,
    P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN,
    P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN,
    P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN,
    P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN,
    P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN,
    P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN,
    P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN,
    P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN,
    P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN,
    P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN,
    P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN,
    P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN,
    P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN,
    P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN,
    P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN,
    P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN,
    P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN,
    P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN,
    P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN,
    P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN,
    P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN,
    P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN,
    P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN,
    P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN,
    P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN,
    P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN,
    P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN,
    P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN,
    P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN,
    P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN,
    P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN,
    P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN,
    P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN,
    P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN,
    P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN,
    P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN,
    P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN,
    P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN,
    P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN,
    P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN,
    P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN,
    P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN,
    P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN,
    P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN,
    P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN,
    P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN,
    P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN,
    P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN,
    BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN,
    BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN,
    BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN,
    BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN,
    BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN,
    BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN,
    BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN,
    BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN,
    BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN,
    BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN,
    BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN,
    BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN,
    BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN,
    BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN,
    BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN,
    BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN,
    BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN,
    BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN,
    BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN,
    BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN,
    BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN,
    READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN,
    P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN,
    P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN,
    P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN,
    P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN,
    P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN,
    P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN,
    P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN,
    P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN,
    P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN,
    P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN,
    P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN,
    P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN,
    P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN,
    P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN,
    P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN,
    P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN,
    P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN,
    P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN,
    P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN,
    P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN,
    P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN,
    P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN,
    P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN,
    P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN,
    P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN,
    P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN,
    P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN,
    P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN,
    P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN,
    P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN,
    P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN,
    P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN,
    P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN,
    P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN,
    P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN,
    P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN,
    P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN,
    P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN,
    P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN,
    P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN,
    P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN,
    P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN,
    P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN,
    P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN,
    P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN,
    P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN,
    P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN,
    P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN,
    P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN,
    P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN,
    P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN,
    P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN,
    P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN,
    P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN,
    P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN,
    P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN,
    P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN,
    P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN,
    P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN,
    P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN,
    P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN,
    P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN,
    P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN,
    P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN,
    P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN,
    P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN,
    P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN,
    P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN,
    P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN,
    P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN,
    P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN,
    P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN,
    P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN,
    P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN,
    P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN,
    P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN,
    P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN,
    P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN,
    P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN,
    P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN,
    P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN,
    P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN,
    P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN,
    P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN,
    P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN,
    P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN,
    P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN,
    P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN,
    P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN,
    P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN,
    P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN,
    P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN,
    P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN,
    P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN,
    P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN,
    P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN,
    P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN,
    P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN,
    P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN,
    P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
    P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
    P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
    P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
    P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
    P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
    P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN,
    P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN,
    P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN,
    P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN,
    P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN,
    P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN,
    P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN,
    P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN,
    P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN,
    P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN,
    P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
    P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
    P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
    P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
    P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
    P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
    P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
    P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
    P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
    P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
    P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
    P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
    P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
    P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
    P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
    P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
    P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
    P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
    P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
    P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
    P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
    P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
    P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
    P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
    P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
    P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
    P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
    P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
    P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
    P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
    P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
    P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
    P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
    P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
    P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
    P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN,
    P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
    P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN,
    P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
    P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN,
    P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
    P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
    P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
    P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
    P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
    P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN,
    P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
    P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN,
    P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
    P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN,
    P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
    P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN,
    P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
    P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN,
    P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
    P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
    P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
    P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
    P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
    P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
    P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
    P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
    P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
    P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
    P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
    P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
    P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
    P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
    P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
    P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
    P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
    P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
    P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
    P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
    P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN,
    P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN,
    P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN,
    P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN,
    P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN,
    P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN,
    P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN,
    P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN,
    P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN,
    P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN,
    P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN,
    P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN,
    P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN,
    P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN,
    P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN,
    P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN,
    P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN,
    P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN,
    P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN,
    P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN,
    P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN,
    P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN,
    P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN,
    P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN,
    P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN,
    P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN,
    P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN,
    P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN,
    P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN,
    P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN,
    P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN,
    P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN,
    P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN,
    P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN,
    P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN,
    P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN,
    P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN,
    P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN,
    P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN,
    P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN,
    P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN,
    P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN,
    P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN,
    P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN,
    P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN,
    P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN,
    P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN,
    P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN,
    P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN,
    P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN,
    P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN,
    P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN,
    P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN,
    P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN,
    P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN,
    P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN,
    P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN,
    P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN,
    P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN,
    P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN,
    P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN,
    P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN,
    P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN,
    P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN,
    P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN,
    P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN,
    P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN,
    P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN,
    P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN,
    P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN,
    P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN,
    P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN,
    P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN,
    P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN,
    P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN,
    P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN,
    P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN,
    P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN,
    P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN,
    P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN,
    P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN,
    P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN,
    P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN,
    P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN,
    P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN,
    P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN,
    P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN,
    P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN,
    P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN,
    P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN,
    P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN,
    P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN,
    P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN,
    P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN,
    P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN,
    P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN,
    P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN,
    P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN,
    P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN,
    P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
    P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
    P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
    P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
    P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
    P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN,
    P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN,
    P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN,
    P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN,
    P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN,
    P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN,
    P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN,
    P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN,
    P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN,
    P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN,
    P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
    P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
    P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
    P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
    P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
    P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
    P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
    P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
    P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
    P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
    P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
    P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
    P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
    P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
    P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
    P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
    P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
    P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
    P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
    P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
    P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
    P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
    P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
    P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
    P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
    P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
    P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
    P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
    P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
    P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
    P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
    P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
    P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
    P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
    P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
    P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
    P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
    P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
    P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
    P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
    P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
    P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
    P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN,
    P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN,
    P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN,
    P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN,
    P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN,
    P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN,
    P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN,
    P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN,
    P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN,
    P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN,
    P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN,
    P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN,
    P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN,
    P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN,
    P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN,
    P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN,
    P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN,
    P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN,
    P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN,
    P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN,
    P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN,
    P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN,
    P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN,
    P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN,
    P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN,
    P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN,
    P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN,
    P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN,
    P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN,
    P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN,
    P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN,
    P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN,
    P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN,
    P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN,
    P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN,
    P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN,
    P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN,
    P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN,
    P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN,
    P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN,
    P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN,
    P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN,
    P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN,
    P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN,
    P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN,
    P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN,
    P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN,
    P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN,
    P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN,
    P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN,
    P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN,
    P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN,
    P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN,
    P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN,
    P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN,
    P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN,
    P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN,
    P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN,
    P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN,
    P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN,
    P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN,
    P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN,
    P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN,
    P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN,
    P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN,
    P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN,
    P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN,
    P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN,
    P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN,
    P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN,
    P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN,
    P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN,
    P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN,
    P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN,
    P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN,
    P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN,
    P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN,
    P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN,
    P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN,
    P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN,
    P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN,
    P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
    U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348, U349,
    U350, U351, U352, U353, U354, U365, U376, U247, U246, U245, U244, U243,
    U242, U241, U240, U239, U238, U237, U236, U235, U234, U233, U232, U231,
    U230, U229, U228, U227, U226, U225, U224, U223, U222, U221, U220, U219,
    U218, U217, U216, U251, U252, U253, U254, U255, U256, U257, U258, U259,
    U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271,
    U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U212,
    U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061,
    P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054,
    P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047,
    P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040,
    P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033,
    P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028,
    P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021,
    P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014,
    P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007,
    P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000,
    P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994,
    P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987,
    P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980,
    P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973,
    P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966,
    P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959,
    P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952,
    P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945,
    P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938,
    P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931,
    P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924,
    P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917,
    P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910,
    P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903,
    P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896,
    P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889,
    P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882,
    P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875,
    P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868,
    P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866,
    P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859,
    P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852,
    P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845,
    P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838,
    P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831,
    P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824,
    P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817,
    P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810,
    P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803,
    P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796,
    P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789,
    P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782,
    P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775,
    P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768,
    P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761,
    P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754,
    P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747,
    P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740,
    P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733,
    P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726,
    P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719,
    P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712,
    P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705,
    P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698,
    P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691,
    P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684,
    P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677,
    P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670,
    P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663,
    P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656,
    P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649,
    P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642,
    P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294,
    P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634,
    P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588,
    P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
    P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
    P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
    P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214,
    P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592,
    P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202,
    P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195,
    P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188,
    P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181,
    P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175,
    P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168,
    P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161,
    P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154,
    P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147,
    P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140,
    P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133,
    P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126,
    P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119,
    P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112,
    P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105,
    P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098,
    P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091,
    P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084,
    P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077,
    P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070,
    P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063,
    P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056,
    P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049,
    P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047,
    P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044,
    P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037,
    P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030,
    P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023,
    P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016,
    P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009,
    P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002,
    P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995,
    P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988,
    P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981,
    P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974,
    P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967,
    P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960,
    P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953,
    P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946,
    P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939,
    P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932,
    P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925,
    P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918,
    P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911,
    P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904,
    P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897,
    P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890,
    P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883,
    P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876,
    P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869,
    P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862,
    P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855,
    P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848,
    P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841,
    P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834,
    P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827,
    P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820,
    P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611,
    P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460,
    P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221,
    P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214,
    P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207,
    P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200,
    P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464,
    P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188,
    P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181,
    P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174,
    P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167,
    P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161,
    P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154,
    P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147,
    P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140,
    P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133,
    P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126,
    P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119,
    P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112,
    P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105,
    P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098,
    P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091,
    P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084,
    P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077,
    P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070,
    P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063,
    P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056,
    P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049,
    P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042,
    P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035,
    P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474,
    P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030,
    P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023,
    P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016,
    P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009,
    P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002,
    P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995,
    P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988,
    P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981,
    P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974,
    P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967,
    P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960,
    P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953,
    P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946,
    P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939,
    P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932,
    P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925,
    P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918,
    P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911,
    P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904,
    P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897,
    P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890,
    P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883,
    P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876,
    P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869,
    P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862,
    P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855,
    P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848,
    P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841,
    P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834,
    P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827,
    P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820,
    P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813,
    P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807,
    P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804,
    P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801;
  wire n43927, n43914, n33474, n43525, n32110, n43813, n42971, n41949,
    n42242, n36904, n27875, n39578, n26498, n43462, n27853, n34270, n26432,
    n24787, n23673, n40080, n40081, n39615, n25897, n24715, n37965, n37279,
    n32334, n24337, n24434, n34552, n23607, n35392, n36320, n22903, n32337,
    n22914, n22919, n36317, n37289, n31721, n43061, n23523, n39892, n23575,
    n36795, n22947, n25634, n23481, n22911, n23463, n28587, n32127, n43408,
    n35715, n26853, n33727, n32119, n22928, n35755, n32506, n26153, n24706,
    n43098, n43100, n26838, n43514, n24610, n24500, n23649, n22923, n22913,
    n28507, n26044, n43054, n33556, n31779, n34569, n41718, n23053, n43750,
    n39522, n41894, n42175, n31718, n26579, n40693, n40350, n23415, n32149,
    n32798, n42708, n39531, n29436, n44019, n43694, n41264, n33548, n31662,
    n42336, n43358, n33545, n43181, n43823, n42939, n43554, n43370, n42838,
    n43595, n43772, n42987, n42685, n43821, n42684, n43771, n42986, n42837,
    n43594, n43366, n43548, n43656, n42593, n43786, n42938, n42496, n28563,
    n43652, n43053, n43545, n43629, n43590, n43784, n43687, n42555, n43145,
    n43030, n28734, n43686, n43628, n42376, n42504, n28556, n42495, n42590,
    n42554, n43221, n43822, n43025, n43219, n43237, n42824, n43538, n43773,
    n42976, n42503, n28856, n28555, n41974, n42009, n42375, n43534, n43630,
    n43008, n43535, n43236, n43328, n41973, n42499, n43023, n43894, n43907,
    n43436, n42008, n43204, n43653, n28851, n28855, n43747, n42535, n28482,
    n42481, n43324, n43531, n43609, n43533, n42963, n42973, n43202, n43785,
    n43007, n42917, n43119, n41750, n43134, n42915, n43602, n42962, n43744,
    n42480, n28479, n28509, n42814, n43593, n42889, n43210, n42673, n41748,
    n43129, n42734, n28481, n43144, n43325, n43203, n41281, n42999, n42643,
    n42853, n42622, n43143, n42472, n42732, n41747, n43208, n43304, n42883,
    n42995, n41280, n28829, n42866, n42867, n43369, n43314, n42229, n42610,
    n43220, n42362, n42577, n41275, n43368, n42631, n42744, n42881, n42316,
    n42298, n42823, n42471, n42951, n43238, n43591, n42609, n42468, n42463,
    n42898, n43170, n43052, n42879, n43009, n42575, n42434, n41716, n42449,
    n42360, n42661, n42448, n42623, n42950, n42470, n42296, n42710, n42630,
    n42435, n42227, n42169, n42450, n42599, n42380, n42422, n42079, n42659,
    n42436, n42706, n42469, n42234, n42037, n41841, n42574, n42482, n42629,
    n28865, n28842, n43051, n43040, n41714, n42869, n42152, n41510, n42127,
    n42627, n42418, n42196, n40807, n42573, n28503, n42604, n28840, n42277,
    n42304, n41712, n42151, n42344, n42647, n42077, n28864, n28475, n42852,
    n42213, n42150, n27935, n42343, n28085, n42562, n41509, n42671, n28502,
    n41891, n28742, n42687, n26576, n28537, n41656, n42416, n42660, n41860,
    n41947, n41765, n42656, n41615, n39567, n43922, n43528, n41687, n28535,
    n41511, n42190, n28741, n42041, n41089, n43889, n42642, n26574, n42398,
    n41945, n41858, n43904, n42207, n43770, n42208, n41713, n43921, n41856,
    n39649, n42462, n41263, n43887, n40103, n25990, n42189, n42621, n42042,
    n43639, n41499, n26560, n43903, n43769, n42397, n39565, n28084, n28835,
    n28518, n27821, n28074, n42069, n43861, n42409, n42205, n42103, n26912,
    n40954, n27934, n40782, n41889, n42512, n41944, n42314, n42270, n41087,
    n41183, n28373, n27818, n39564, n25988, n43133, n41910, n41699, n28517,
    n43638, n41227, n43916, n41493, n40101, n43703, n43819, n43899, n43782,
    n42269, n38813, n43627, n43888, n41258, n28463, n27848, n42064, n26559,
    n28372, n41771, n40953, n39648, n42098, n42097, n42182, n43434, n41423,
    n41256, n41736, n43626, n42203, n41943, n43818, n43685, n41908, n38665,
    n42813, n28491, n39713, n42063, n27846, n28772, n43702, n27755, n26908,
    n42388, n42281, n28525, n41960, n41567, n42505, n41492, n39930, n41735,
    n28490, n42386, n43684, n39669, n41169, n42342, n41422, n40939, n42812,
    n39560, n43200, n27753, n41906, n43118, n40766, n28106, n41443, n26707,
    n43650, n28769, n38664, n42888, n41248, n41459, n40879, n42340, n41166,
    n43199, n28767, n39925, n43322, n41416, n26705, n27887, n41953, n41037,
    n28103, n40765, n40153, n41079, n41201, n40097, n42093, n39590, n41840,
    n43117, n41246, n40955, n41845, n38803, n28101, n39769, n26719, n42335,
    n37567, n40123, n43589, n25490, n38135, n41035, n43544, n38381, n27029,
    n41457, n41839, n41165, n41244, n37448, n37128, n38801, n41678, n28765,
    n43235, n40846, n41614, n27833, n41123, n39588, n41668, n28763, n40844,
    n43215, n38802, n40869, n43233, n41194, n41112, n41268, n40118, n41155,
    n41764, n41255, n40721, n41143, n26681, n41224, n42334, n41033, n39712,
    n39767, n37738, n39707, n26596, n41031, n41141, n37505, n43587, n42913,
    n37563, n27744, n40719, n43006, n36911, n40842, n41254, n41667, n42958,
    n40863, n41562, n37352, n37827, n41611, n41763, n41561, n40840, n39185,
    n39161, n39198, n40858, n38267, n39143, n39169, n41237, n39177, n39151,
    n39136, n41152, n41139, n40717, n37473, n37733, n43004, n42730, n38997,
    n42864, n39026, n39013, n38990, n26139, n36909, n40700, n38640, n39005,
    n43021, n38967, n26712, n38395, n39011, n39133, n39614, n39238, n39024,
    n40839, n39291, n38252, n41559, n39183, n39196, n39258, n38928, n39249,
    n39159, n36131, n38962, n37732, n39003, n37278, n39141, n39167, n38985,
    n40862, n39175, n40755, n39149, n40791, n42533, n37557, n26082, n24761,
    n39209, n41137, n39762, n36099, n39266, n37009, n38244, n38995, n39935,
    n39276, n42477, n37472, n38752, n41557, n37845, n40819, n37932, n38760,
    n41238, n37747, n26086, n37877, n37254, n37234, n39610, n26939, n38303,
    n40065, n38206, n37893, n37787, n37804, n38315, n37007, n37885, n37633,
    n38003, n37901, n38243, n39289, n26501, n38812, n39236, n37972, n38780,
    n37987, n38233, n38901, n37120, n38249, n39256, n27743, n38198, n38922,
    n39247, n39264, n39274, n38219, n40753, n37979, n38011, n42911, n37351,
    n38276, n40496, n28761, n24759, n26092, n38768, n37814, n26080, n39204,
    n38251, n40853, n42532, n40860, n39684, n37822, n37795, n38744, n37995,
    n38302, n38571, n38796, n38765, n36125, n38215, n38388, n39192, n38981,
    n38572, n37842, n38001, n38273, n37864, n43019, n37985, n38311, n38203,
    n39598, n38292, n38776, n37801, n37004, n37252, n36547, n27863, n37744,
    n26938, n37277, n38757, n38248, n37888, n39609, n37959, n37631, n25993,
    n37927, n38741, n37880, n38367, n37811, n38579, n38966, n38580, n38195,
    n37977, n38587, n42877, n42358, n39683, n38588, n37792, n38351, n38009,
    n40816, n38989, n38749, n38359, n38232, n38343, n37784, n37819, n37896,
    n26085, n38272, n37383, n37971, n37391, n36852, n38740, n40054, n38310,
    n37530, n27862, n37200, n38692, n37931, n37407, n37892, n37211, n37152,
    n37390, n39208, n42293, n36279, n40485, n37251, n37900, n37595, n37606,
    n38291, n37425, n38202, n38242, n38775, n39130, n38711, n38756, n37800,
    n37382, n37841, n37399, n40752, n38940, n38194, n38583, n37818, n37876,
    n38720, n38214, n37743, n37398, n37192, n37791, n38674, n37884, n38748,
    n37168, n37176, n38764, n37184, n38683, n37783, n38701, n37160, n37810,
    n38170, n37850, n43872, n41018, n37386, n37555, n37745, n40757, n43844,
    n38313, n42619, n25066, n38301, n39804, n35363, n27737, n37590, n43474,
    n40086, n40751, n39439, n43804, n37521, n38241, n37370, n36399, n36854,
    n39129, n37394, n28162, n40483, n42517, n37467, n38027, n38807, n43838,
    n43843, n43871, n42432, n37589, n38209, n43868, n38770, n37861, n26483,
    n38165, n41015, n42985, n37956, n38306, n39802, n37835, n37836, n38300,
    n25797, n42225, n39283, n40541, n38228, n39120, n39435, n40469, n43802,
    n38328, n43303, n26339, n38190, n39612, n40538, n40002, n37272, n37001,
    n43302, n37873, n37379, n39991, n40467, n38236, n37860, n40013, n39980,
    n40435, n40051, n38287, n39969, n36090, n37423, n41014, n42287, n37955,
    n39799, n37215, n42850, n43573, n37968, n40024, n40035, n38337, n41886,
    n39124, n43870, n26338, n39434, n39845, n37588, n38875, n37615, n39877,
    n39861, n38859, n38164, n39890, n38896, n38843, n38883, n39837, n38186,
    n39829, n38851, n37628, n39853, n39869, n38867, n43840, n38049, n35331,
    n37044, n38435, n38089, n38073, n38105, n38427, n38097, n38121, n40537,
    n38419, n38113, n40433, n38223, n26458, n38459, n37963, n39423, n39460,
    n43834, n39112, n28726, n43830, n37779, n38185, n43671, n38620, n40085,
    n38930, n41012, n37145, n37205, n37941, n40644, n38045, n42494, n42669,
    n38336, n38451, n37366, n38443, n38134, n39797, n38480, n37868, n38467,
    n38081, n38295, n37574, n43751, n36376, n38282, n40536, n37043, n37608,
    n37037, n35329, n38222, n38618, n39111, n35816, n38631, n36118, n43663,
    n37138, n37144, n40257, n37645, n41938, n39419, n42553, n40691, n39457,
    n43604, n39530, n36274, n38322, n37769, n37949, n40430, n43836, n28828,
    n37856, n36568, n38177, n43826, n27859, n36738, n38044, n36575, n40429,
    n41730, n36749, n39417, n37855, n43190, n38221, n43603, n39456, n38320,
    n36737, n37573, n38281, n38151, n42633, n40041, n37657, n43669, n38933,
    n43749, n28674, n36656, n40601, n39882, n37643, n39514, n42007, n42491,
    n39602, n37948, n37028, n42333, n35321, n37365, n38888, n38043, n36574,
    n36370, n36088, n43662, n40078, n39110, n27732, n37026, n41307, n39377,
    n41221, n39415, n42665, n38616, n39527, n35780, n40622, n36206, n39817,
    n42332, n25115, n41563, n39955, n43670, n37493, n36654, n42980, n38305,
    n36565, n37033, n37571, n38126, n28768, n38149, n38174, n42057, n35327,
    n43189, n43180, n39455, n38472, n42137, n39101, n43376, n38959, n35326,
    n39543, n37492, n38497, n42937, n40666, n39042, n42329, n26383, n43179,
    n39187, n42056, n37045, n42132, n41867, n42054, n38409, n39413, n43178,
    n28753, n36736, n39313, n38061, n35806, n35832, n43194, n38030, n41933,
    n42027, n37147, n39015, n37854, n38150, n43186, n42646, n39952, n24721,
    n24723, n24869, n38173, n43657, n37642, n39815, n28474, n38407, n26360,
    n43606, n35323, n43185, n42117, n41685, n28671, n43188, n38056, n41553,
    n42004, n41866, n36744, n39309, n42131, n37131, n39951, n35778, n42133,
    n42327, n42055, n39040, n38495, n41534, n37491, n28752, n35602, n25978,
    n43348, n40880, n35517, n25973, n36109, n28102, n38172, n39814, n38148,
    n36652, n42022, n43177, n25965, n38066, n24741, n40349, n34521, n41122,
    n42309, n36793, n40852, n40096, n42129, n34063, n38412, n41249, n28097,
    n34813, n37490, n39589, n25976, n39810, n41529, n37572, n42020, n37859,
    n34585, n39947, n43536, n23700, n24672, n42040, n40407, n28059, n38064,
    n40151, n38494, n24720, n43209, n24742, n42568, n25963, n39039, n35432,
    n28751, n42374, n42325, n42975, n42836, n28732, n41552, n34131, n42019,
    n40482, n25110, n41995, n39809, n40404, n36152, n34094, n28228, n26402,
    n24739, n35627, n42021, n42331, n27756, n39945, n40976, n40345, n38054,
    n40582, n35324, n39304, n42324, n24754, n28853, n41865, n38493, n35155,
    n41067, n28096, n26369, n28749, n26379, n39038, n41013, n41424, n38410,
    n26422, n41234, n43173, n40539, n26423, n40094, n26580, n28090, n26416,
    n37489, n26417, n26408, n42905, n43207, n43530, n41530, n41121, n41528,
    n26401, n42907, n26395, n39303, n26409, n41549, n38053, n26418, n38835,
    n40754, n26419, n26406, n26403, n40520, n26400, n42017, n26413, n26414,
    n43182, n40402, n26415, n34511, n42408, n33733, n38491, n42589, n41009,
    n34652, n41683, n42330, n36556, n41064, n35774, n39126, n26349, n42715,
    n26351, n26356, n28554, n26363, n26367, n26373, n39037, n39943, n41770,
    n26421, n40327, n38402, n41415, n40428, n41187, n40147, n39808, n40578,
    n26566, n28095, n40974, n40480, n28748, n37487, n27823, n41120, n40255,
    n40468, n41558, n28754, n40236, n41526, n40530, n40535, n42015, n34343,
    n41154, n41387, n41512, n34269, n42714, n23664, n26394, n40534, n42997,
    n43807, n43472, n27350, n26399, n40427, n41393, n26348, n26347, n39798,
    n27040, n42683, n41555, n41153, n28744, n34507, n40572, n41413, n38401,
    n26250, n24618, n41548, n43444, n41168, n42900, n24840, n39035, n28891,
    n38296, n24716, n37623, n42719, n27720, n40464, n26362, n38927, n39795,
    n26412, n39794, n40232, n23661, n40526, n26292, n42990, n42718, n43447,
    n42586, n39454, n41006, n40400, n26239, n41972, n41236, n40465, n41411,
    n41114, n40478, n41232, n42464, n40516, n37638, n39424, n41229, n40249,
    n41378, n40818, n42965, n44020, n42712, n27751, n43437, n43791, n38925,
    n40409, n33731, n43012, n35769, n41458, n42717, n24615, n40524, n40475,
    n39792, n39420, n43567, n39452, n24623, n39442, n38176, n40964, n39414,
    n41969, n42280, n40460, n42537, n40999, n34502, n42466, n28766, n40545,
    n42250, n37591, n28557, n41746, n22916, n41242, n40248, n24816, n24614,
    n28756, n37021, n38790, n42527, n42383, n28869, n28838, n42538, n42346,
    n42278, n42254, n43371, n43853, n41935, n38175, n42892, n42558, n33725,
    n42592, n39743, n27750, n38188, n41902, n40770, n42930, n40414, n38047,
    n41451, n42178, n42652, n41450, n38924, n40088, n42258, n42727, n24575,
    n24419, n37085, n28877, n40092, n37637, n41942, n33724, n42966, n41214,
    n42249, n41239, n41373, n39557, n41019, n42171, n43617, n23697, n42584,
    n41073, n42676, n41124, n42121, n41888, n35361, n42122, n42248, n43559,
    n28216, n38279, n41934, n41931, n39640, n41369, n39785, n41859, n36542,
    n34489, n41977, n42252, n42385, n41453, n41946, n28886, n36173, n43797,
    n37713, n43386, n41965, n36890, n39389, n43788, n40841, n40982, n41368,
    n42240, n43165, n39635, n34485, n40669, n36895, n40388, n28882, n41926,
    n36866, n31796, n35172, n23693, n43767, n35178, n36543, n37325, n43148,
    n42246, n42400, n43158, n41271, n43748, n43876, n32145, n27749, n28559,
    n27713, n24801, n41357, n38781, n40883, n41283, n26254, n42198, n40436,
    n23542, n41290, n42662, n42539, n42236, n42092, n36403, n41302, n39934,
    n38553, n38885, n41295, n39098, n40894, n40907, n40906, n39549, n43372,
    n39732, n41921, n41869, n41879, n39535, n38650, n43716, n36459, n39240,
    n38703, n40500, n39883, n35962, n36167, n34124, n39388, n40042, n40881,
    n41318, n43331, n40277, n40186, n41358, n43341, n41976, n40205, n26550,
    n41204, n34287, n32341, n39251, n42927, n38687, n35959, n41370, n39200,
    n39241, n42185, n39280, n39230, n43732, n37808, n42802, n41356, n43333,
    n23540, n25944, n39378, n33786, n32144, n42235, n40242, n42244, n42201,
    n36177, n27706, n42091, n26057, n41339, n44021, n39959, n42305, n36955,
    n41296, n39390, n35553, n41756, n43693, n38411, n42085, n26051, n24501,
    n22946, n39790, n27709, n39036, n37302, n34876, n24612, n35719, n43362,
    n40275, n41920, n41352, n41336, n39541, n36237, n40899, n42804, n36794,
    n43523, n26206, n43911, n40607, n43698, n24766, n43697, n25102, n42083,
    n39030, n35421, n39394, n43709, n27702, n31795, n31960, n27705, n37476,
    n35594, n27754, n26064, n40375, n35465, n26048, n41338, n36078, n41335,
    n44023, n43719, n36867, n40652, n35940, n31821, n43915, n39387, n42090,
    n24129, n36077, n41327, n41496, n26062, n43707, n31684, n34808, n34404,
    n31722, n37486, n26204, n24562, n43809, n24479, n43718, n34495, n38482,
    n41912, n35967, n39302, n41326, n35658, n26047, n41333, n28323, n31681,
    n24401, n38334, n28338, n34335, n28819, n39481, n31913, n40270, n28088,
    n40373, n44091, n40372, n33262, n34651, n28199, n40762, n44003, n33917,
    n35601, n35431, n33208, n28226, n39453, n28093, n28764, n31820, n41245,
    n25073, n36205, n35970, n27344, n37264, n41329, n24803, n40935, n27893,
    n35656, n24336, n39920, n36257, n41223, n39756, n27923, n35261, n41732,
    n35249, n41078, n28315, n28657, n27921, n28308, n27900, n28715, n28235,
    n26529, n39448, n27907, n24811, n28242, n26543, n28275, n28281, n39727,
    n31818, n28268, n27889, n28288, n28295, n26536, n28147, n38595, n28261,
    n34966, n43293, n28301, n28758, n28746, n35989, n28255, n28248, n27914,
    n36046, n28322, n36045, n41342, n31361, n32938, n32794, n35935, n23647,
    n23615, n41005, n33951, n35532, n28299, n28286, n32792, n23642, n35527,
    n32752, n31927, n40508, n35744, n28279, n28293, n28266, n41345, n41231,
    n27346, n28150, n36043, n28834, n35951, n26202, n32838, n27882, n23613,
    n28816, n31682, n35667, n28107, n26201, n32871, n28043, n23622, n23629,
    n35944, n28613, n36509, n36333, n28714, n35462, n42322, n32716, n36038,
    n24444, n34659, n36967, n32330, n27879, n31322, n31344, n27872, n32494,
    n32680, n34655, n28143, n26205, n28041, n36338, n36239, n25573, n34536,
    n26189, n26492, n23515, n31817, n32865, n36022, n36243, n36871, n26514,
    n34673, n28654, n28612, n40125, n28152, n28039, n32861, n33906, n40872,
    n36242, n28414, n35930, n27340, n33630, n36154, n23621, n28108, n34340,
    n24441, n36153, n26181, n23514, n23722, n34671, n36490, n24340, n26493,
    n31196, n31202, n41520, n32671, n33801, n23588, n34638, n24252, n27337,
    n26489, n28459, n36019, n42320, n32870, n32372, n34637, n26180, n32849,
    n35947, n23717, n31273, n27338, n27973, n36660, n33496, n27028, n33310,
    n28413, n41403, n33802, n26198, n27679, n23265, n33500, n26477, n34979,
    n28109, n32251, n24431, n26478, n32550, n31777, n23263, n40734, n27678,
    n28036, n31920, n31911, n41531, n32202, n33823, n25554, n23596, n28265,
    n28239, n26331, n23719, n28258, n23926, n26679, n31894, n28232, n24174,
    n26445, n24175, n27918, n27972, n33824, n26525, n28245, n27617, n31276,
    n27330, n27910, n23219, n32200, n27904, n26533, n23628, n27676, n27813,
    n28252, n26980, n27897, n28110, n26456, n24204, n23284, n41397, n26540,
    n23595, n40744, n24214, n35377, n27615, n23179, n26330, n26711, n33953,
    n43394, n36374, n39700, n39909, n26982, n32196, n40415, n32263, n28163,
    n23581, n36830, n26457, n24247, n23180, n35443, n37270, n26196, n25540,
    n23922, n25541, n37535, n33783, n36828, n32344, n23531, n23716, n36970,
    n32889, n31824, n28079, n26551, n23177, n39759, n24245, n41208, n34902,
    n27609, n25563, n34986, n23178, n27801, n25722, n25764, n37464, n23134,
    n26913, n25736, n23135, n26979, n41472, n35316, n25026, n23914, n27325,
    n27727, n26137, n31534, n25063, n40442, n41927, n25113, n37499, n26459,
    n37444, n33555, n32799, n23492, n31670, n26228, n24244, n25839, n23218,
    n23696, n27717, n27733, n25750, n34835, n26227, n25060, n24949, n26032,
    n26981, n36667, n28706, n25730, n25546, n25744, n34985, n41362, n41147,
    n25022, n27811, n25539, n26637, n25560, n28415, n27974, n27799, n26135,
    n27037, n27034, n26688, n23912, n26685, n28050, n26145, n28053, n23176,
    n23273, n26036, n41784, n23925, n28468, n23173, n23688, n25942, n23283,
    n25939, n25844, n28471, n25088, n23656, n24243, n25085, n24139, n25082,
    n25757, n25771, n25079, n23549, n27734, n24196, n23915, n26507, n24168,
    n24187, n24216, n24193, n24181, n24178, n42978, n27731, n24184, n36249,
    n24190, n23913, n24839, n26226, n26684, n23911, n23279, n23921, n26144,
    n23924, n25074, n26598, n23272, n27681, n23221, n24826, n26035, n27324,
    n25785, n35435, n24713, n24116, n25776, n25675, n24177, n25716, n26487,
    n25630, n25742, n24167, n27816, n24095, n31790, n27878, n25769, n25592,
    n28615, n28112, n24334, n34531, n25578, n25934, n26031, n25530, n42318,
    n25552, n25755, n32175, n25728, n25571, n23687, n23928, n23175, n26466,
    n23670, n37468, n31907, n24849, n23920, n27669, n24837, n25720, n23559,
    n23946, n23901, n24824, n24142, n24779, n25072, n40586, n27674, n23594,
    n32082, n24800, n23660, n31896, n24814, n23558, n25543, n41546, n27888,
    n40606, n25535, n25529, n41212, n26093, n28604, n25557, n23216, n27342,
    n25581, n33848, n26462, n33564, n25930, n23278, n24331, n28135, n39927,
    n34498, n32177, n23491, n24239, n32367, n35437, n24611, n23565, n27597,
    n27814, n23543, n27329, n37735, n25713, n27606, n27326, n24911, n24731,
    n24114, n24711, n24986, n24172, n39210, n27664, n39480, n31787, n24947,
    n26429, n31910, n25893, n40738, n24847, n24708, n24482, n22944, n27802,
    n31788, n24559, n27787, n26916, n23902, n24835, n27629, n23919, n24162,
    n24657, n35819, n24608, n31525, n24857, n24165, n33666, n26058, n26385,
    n27322, n25025, n23577, n31808, n24389, n28113, n24166, n27331, n27612,
    n31793, n24778, n27619, n23449, n24807, n25094, n23652, n31895, n23524,
    n24909, n25834, n24984, n25928, n24794, n23889, n23703, n26224, n23262,
    n24332, n31809, n26285, n22904, n31498, n24654, n31806, n33915, n27655,
    n24211, n23503, n25024, n24817, n27785, n24867, n24207, n24161, n23576,
    n24237, n24234, n26178, n27332, n24822, n23934, n25838, n33688, n24119,
    n23447, n24221, n24481, n24111, n27661, n24709, n32206, n26030, n33585,
    n27791, n35436, n27866, n24775, n25892, n24560, n27596, n23728, n23545,
    n27628, n23497, n24793, n28133, n26225, n24395, n36202, n27618, n24297,
    n31511, n24330, n23513, n28114, n31666, n40052, n24396, n35974, n27250,
    n37119, n24871, n27666, n27592, n24112, n35267, n32868, n27789, n32199,
    n27599, n34097, n26327, n27775, n27630, n26449, n37754, n43721, n26173,
    n24102, n25932, n24831, n24236, n25889, n31804, n38968, n38013, n22900,
    n41789, n35858, n25235, n34134, n27658, n25236, n38140, n23120, n23445,
    n23214, n43475, n23511, n25266, n25146, n23166, n27616, n25623, n27604,
    n32489, n27796, n27626, n24802, n24150, n34226, n25885, n32848, n34187,
    n25206, n27803, n28131, n24393, n32860, n33738, n25668, n23260, n24135,
    n23167, n25190, n23848, n25651, n23121, n23241, n25205, n23119, n24097,
    n27180, n23384, n24658, n24980, n31193, n25265, n23215, n25691, n25296,
    n28115, n25667, n25527, n23259, n25297, n25128, n27781, n24943, n34149,
    n23165, n23213, n25175, n25709, n37575, n25604, n24392, n41790, n25622,
    n27659, n25145, n23787, n27773, n25250, n24905, n27213, n27143, n27764,
    n23240, n23236, n24568, n27499, n27769, n27281, n27142, n28130, n27470,
    n27590, n37016, n23257, n24653, n24704, n24475, n23258, n24476, n23300,
    n24605, n25189, n23102, n25640, n25620, n23101, n25621, n23113, n25264,
    n25684, n23432, n25249, n24328, n27197, n25708, n25666, n25707, n24606,
    n24327, n25204, n27078, n23152, n25143, n25144, n23151, n23474, n25129,
    n27112, n25161, n24652, n25600, n25203, n25528, n23200, n27163, n27247,
    n24705, n33067, n25526, n23201, n24016, n24689, n23192, n24688, n24703,
    n23269, n23255, n23256, n23249, n24651, n23461, n23318, n23164, n24636,
    n23093, n23100, n23099, n23423, n23393, n24603, n27077, n27423, n24325,
    n27439, n27164, n23785, n27162, n25699, n27454, n25706, n27246, n24295,
    n24589, n23784, n24386, n27111, n24385, n27092, n27772, n24312, n27763,
    n27189, n27196, n27762, n24294, n27212, n24326, n27589, n24474, n27558,
    n24590, n27500, n27264, n25661, n27560, n25665, n27127, n27929, n27394,
    n24459, n27530, n27378, n27265, n27497, n27528, n24460, n27280, n27141,
    n25512, n36873, n25522, n27469, n27574, n25650, n24557, n31063, n25525,
    n24075, n25513, n27179, n24558, n23462, n23209, n24293, n23879, n27093,
    n27064, n27076, n23473, n23118, n25649, n36558, n24465, n24582, n25648,
    n23844, n24066, n28128, n24458, n24074, n23846, n25521, n24452, n39901,
    n24555, n24650, n24536, n24088, n27056, n24604, n27057, n24635, n24272,
    n25603, n24000, n23161, n25618, n24634, n24855, n25690, n25700, n25698,
    n25702, n23775, n25701, n25705, n27245, n24273, n24588, n23783, n25503,
    n24643, n25502, n27219, n25511, n25510, n25639, n24473, n27150, n27437,
    n23337, n27438, n27421, n24324, n36222, n23254, n24317, n23251, n23252,
    n23248, n27210, n27424, n23394, n27211, n24311, n23250, n27195, n27767,
    n27186, n24304, n27133, n27407, n27408, n27565, n27140, n27573, n27126,
    n27393, n27385, n24512, n27588, n27119, n27587, n27514, n27496, n27513,
    n27519, n27527, n42522, n27498, n27364, n27483, n27363, n27257, n27369,
    n27377, n27544, n27484, n27543, n27263, n27550, n27177, n27557, n27467,
    n27468, n23931, n27279, n24680, n27178, n27453, n24702, n27278, n27161,
    n27155, n27091, n24362, n23306, n23212, n27109, n23268, n23362, n23431,
    n24637, n24981, n27110, n23424, n27361, n27585, n27225, n27586, n27218,
    n27579, n25509, n27506, n27505, n27525, n27370, n27520, n23782, n27362,
    n27215, n27224, n23916, n24472, n27511, n27116, n27356, n27526, n27512,
    n27355, n27580, n24471, n27376, n24086, n27436, n24535, n24087, n27435,
    n24523, n27276, n24524, n27277, n27445, n24079, n27270, n24025, n23929,
    n27271, n27460, n24553, n24081, n27262, n27259, n27476, n27475, n27482,
    n24448, n27481, n24556, n27490, n24447, n27489, n24451, n24073, n27495,
    n28116, n24064, n27386, n24454, n27138, n24457, n27139, n27392, n27391,
    n27400, n27132, n27399, n27129, n24466, n27406, n23843, n27405, n27124,
    n27566, n27125, n24463, n25519, n27571, n27074, n24318, n27208, n27209,
    n27202, n23878, n27203, n24309, n24310, n27194, n24303, n24281, n27191,
    n24299, n24300, n27184, n24384, n27107, n27085, n27108, n24292, n27102,
    n27084, n27090, n27087, n27375, n24262, n25704, n27536, n27237, n27535,
    n25695, n27542, n27175, n27541, n27243, n27176, n23776, n25688, n25689,
    n27549, n27242, n27556, n25683, n25680, n27555, n27169, n27170, n27159,
    n27160, n29835, n27156, n27147, n27148, n25596, n24271, n27047, n23815,
    n27046, n27055, n23756, n24056, n27054, n24323, n24319, n27065, n27063,
    n24316, n27075, n23058, n23205, n23072, n24628, n23116, n23457, n23109,
    n22926, n23094, n23472, n23156, n23471, n23476, n24944, n24642, n23479,
    n24649, n24648, n25659, n25662, n23989, n23034, n23390, n23024, n23400,
    n23399, n23341, n23333, n23327, n23405, n23328, n24681, n23408, n23420,
    n23430, n23429, n23988, n23434, n23358, n24511, n23368, n23367, n23999,
    n23253, n26827, n26837, n26831, n23305, n26852, n23246, n23239, n23237,
    n27429, n23961, n37853, n30874, n36182, n24026, n27416, n27415, n27422,
    n27430, n24006, n24581, n24005, n23038, n25637, n23233, n23335, n24554,
    n29304, n23331, n23023, n23032, n23029, n24261, n24533, n24534, n23030,
    n23026, n24629, n24545, n24450, n24449, n39311, n28126, n24456, n24462,
    n24461, n23016, n24464, n24468, n24467, n24470, n26841, n43880, n23324,
    n39188, n23323, n23326, n25696, n23332, n25682, n25677, n27471, n24322,
    n28934, n24320, n24315, n23893, n24313, n24314, n24307, n27432, n27427,
    n24308, n27419, n24306, n24301, n24302, n27758, n28775, n39279, n27474,
    n42524, n27354, n27522, n27517, n27371, n27532, n27534, n27575, n27576,
    n27567, n27404, n27401, n27395, n24291, n24280, n24439, n24270, n23654,
    n35805, n41877, n24290, n24020, n27275, n27272, n27268, n24019, n27266,
    n24023, n27267, n27261, n24035, n27253, n27136, n27134, n27130, n27131,
    n27128, n27122, n27123, n27120, n23983, n24906, n23982, n23986, n23998,
    n27089, n27086, n23854, n27082, n27083, n27080, n23869, n32845, n27072,
    n27067, n27062, n27059, n27060, n27052, n27053, n27050, n23751, n27044,
    n27045, n23750, n27042, n23755, n23814, n27043, n23766, n23765, n27241,
    n27238, n27239, n27233, n27234, n27222, n27223, n27220, n23792, n27216,
    n27217, n27214, n24065, n24069, n24068, n24072, n23821, n24077, n24076,
    n23819, n23820, n24078, n24085, n24546, n24047, n27173, n27174, n27171,
    n27172, n27167, n27168, n27165, n27149, n24046, n24057, n24055, n27207,
    n27204, n27205, n27200, n27201, n27198, n27192, n27193, n27190, n23855,
    n29461, n27105, n27106, n27103, n27098, n27099, n27088, n27728, n23419,
    n23422, n23426, n23425, n23428, n23470, n23433, n23465, n26818, n23466,
    n23304, n23357, n23456, n43711, n43367, n23360, n43361, n23965, n23364,
    n23960, n23293, n23956, n23460, n43137, n23389, n23392, n23064, n23060,
    n23396, n23395, n22906, n23475, n28943, n23398, n23953, n23066, n23063,
    n23407, n23057, n23754, n23858, n24249, n28156, n24507, n24469, n34718,
    n23880, n23753, n24305, n23868, n23805, n23810, n23864, n23865, n23809,
    n23825, n24455, n23826, n23822, n43246, n37485, n39016, n24070, n24071,
    n43275, n23600, n23781, n23791, n23796, n24321, n23763, n22988, n23764,
    n27236, n23760, n36415, n27766, n23418, n23427, n23436, n23356, n23290,
    n41374, n23997, n23992, n23993, n23987, n23303, n23056, n39775, n23065,
    n24861, n23455, n38207, n23959, n26848, n23958, n28117, n26858, n23478,
    n23469, n25678, n23859, n24054, n24050, n23325, n24051, n24044, n24045,
    n23343, n24040, n23022, n24041, n23031, n37834, n23388, n24034, n23397,
    n24029, n24030, n23410, n24024, n22979, n22909, n39097, n22910, n23017,
    n23015, n24100, n23014, n22901, n27097, n37933, n37542, n24227, n26791,
    n41145, n22917, n24250, n22980, n41516, n23329, n22915, n23686, n23827,
    n23346, n37851, n23777, n22986, n23828, n24209, n23020, n27240, n39529,
    n23671, n39113, n26214, n42023, n23759, n38220, n22977, n27927, n38481,
    n27066, n23811, n24437, n23620, n23123, n22902, n23353, n22952, n42626,
    n23453, n24852, n38884, n23377, n36289, n23995, n27274, n23002, n23012,
    n23996, n23001, n26807, n23899, n22966, n27095, n23054, n23013, n43094,
    n24033, n35624, n27206, n23046, n23386, n23403, n43033, n22978, n23900,
    n22967, n23482, n28608, n27144, n23416, n36286, n24032, n23439, n27776,
    n23539, n22964, n27777, n23122, n44100, n34909, n22972, n22965, n23849,
    n36048, n26587, n22993, n27759, n22973, n23008, n23000, n27071, n22994,
    n40168, n23850, n42214, n29574, n23271, n23892, n27771, n29308, n40221,
    n22999, n41375, n23937, n32190, n22959, n23011, n39524, n23103, n23679,
    n31938, n29580, n38316, n23105, n23619, n22951, n22976, n22953, n22987,
    n22958, n23226, n39946, n23007, n22985, n24505, n43146, n24843, n43612,
    n37805, n42547, n37629, n22996, n22998, n42321, n22997, n22995, n22948,
    n43097, n33537, n43082, n23006, n23005, n41230, n26779, n22990, n43093,
    n23003, n22989, n35254, n23010, n22992, n23009, n22991, n23004, n42337,
    n22968, n42786, n22971, n23104, n39511, n28129, n36357, n42070, n34677,
    n38321, n24707, n22970, n32075, n28132, n37475, n22975, n23637, n40527,
    n22974, n39937, n37634, n35452, n22982, n32083, n23579, n22984, n22983,
    n37635, n31055, n23684, n33579, n39114, n22950, n41597, n22949, n39944,
    n41578, n22955, n22954, n24830, n32336, n22957, n22956, n22961, n22960,
    n35163, n23626, n22963, n41513, n22962, n22969, n42104, n29752, n39440,
    n26060, n23994, n23991, n23990, n23985, n23984, n23981, n27880, n27235,
    n41023, n33714, n26059, n33710, n41128, n40959, n42707, n40403, n27048,
    n41072, n35608, n23980, n38277, n35663, n35728, n29055, n33933, n43867,
    n43895, n43731, n43717, n43342, n28743, n28866, n43820, n42933, n42832,
    n42977, n43651, n43050, n43455, n43142, n43705, n28857, n43783, n28492,
    n43866, n43453, n43529, n43641, n42585, n28519, n28504, n43640, n43925,
    n42487, n42821, n43216, n42974, n43643, n42549, n28510, n28848, n43022,
    n42486, n43522, n43476, n43806, n43387, n43323, n43201, n42534, n41952,
    n28895, n28508, n42959, n43598, n41951, n42914, n42916, n43552, n42885,
    n43592, n42733, n42672, n43383, n27834, n42800, n42865, n43057, n42731,
    n42854, n42840, n43572, n43597, n28873, n43551, n42880, n43024, n42315,
    n42228, n42297, n43380, n28675, n42822, n42536, n28727, n42359, n42295,
    n42433, n42128, n41186, n42608, n42878, n42226, n41669, n28870, n42447,
    n41679, n43550, n41846, n42897, n42168, n42696, n42720, n42233, n42989,
    n42705, n43039, n42379, n42563, n40806, n42572, n42625, n41711, n41269,
    n41696, n28839, n42276, n42126, n26940, n42378, n42750, n27824, n42051,
    n42670, n28060, n41619, n28075, n39585, n42415, n42851, n42624, n28464,
    n43527, n28534, n42058, n42641, n26573, n41434, n41182, n42511, n42461,
    n41855, n39685, n41781, n42620, n42284, n39717, n40781, n43766, n42664,
    n28371, n27041, n41939, n25987, n41088, n28045, n43781, n40066, n43132,
    n41772, n40497, n40071, n26557, n40100, n41048, n42181, n28225, n39562,
    n41488, n39645, n42095, n38806, n39599, n41490, n41470, n41222, n41734,
    n27845, n42307, n26695, n27869, n41959, n38902, n41566, n39673, n42062,
    n25798, n41461, n27752, n41077, n41905, n41225, n40783, n41731, n43611,
    n38661, n27030, n39672, n40558, n39293, n38897, n43625, n43681, n43649,
    n39665, n42887, n41844, n41200, n43198, n26704, n40934, n40937, n26152,
    n43321, n41677, n39922, n37564, n41613, n39587, n26558, n41243, n41455,
    n27746, n43543, n42319, n39926, n26040, n39586, n28100, n39768, n27857,
    n27856, n41030, n27745, n28762, n37561, n39921, n37503, n40070, n39907,
    n43586, n39757, n36908, n40855, n40716, n38638, n26090, n40856, n41151,
    n38394, n38266, n25092, n39689, n38960, n38983, n36126, n39023, n41148,
    n39010, n41150, n39002, n42725, n41253, n26389, n41136, n38994, n40115,
    n40854, n36097, n37349, n37993, n39688, n40494, n39273, n38810, n42294,
    n39235, n39263, n37218, n44012, n39288, n26079, n39020, n39246, n39202,
    n39703, n39255, n40064, n39176, n37878, n39142, n37894, n41076, n36122,
    n37886, n37460, n39150, n27861, n38577, n38898, n38585, n39168, n39596,
    n27741, n42876, n36861, n38907, n39197, n37925, n38794, n38372, n38205,
    n39184, n38808, n38218, n38569, n38197, n37862, n39284, n39134, n37245,
    n27868, n38906, n26340, n36859, n38217, n27865, n37630, n37265, n36857,
    n36487, n36092, n41309, n42640, n37848, n36860, n43443, n42875, n37726,
    n36396, n37206, n40891, n38938, n39364, n40258, n39096, n37597, n39332,
    n39109, n38856, n37604, n39965, n38864, n38872, n39340, n37621, n38848,
    n43837, n37214, n38840, n39348, n38880, n38152, n38892, n39874, n39072,
    n39080, n37416, n39532, n39866, n26332, n40046, n39998, n39088, n39834,
    n39324, n39048, n40009, n39385, n40020, n39987, n39826, n39886, n39858,
    n37547, n39976, n39850, n39356, n39064, n39372, n39056, n40031, n39842,
    n38102, n38524, n38432, n38532, n42983, n37539, n38540, n38130, n38416,
    n38508, n38118, n28223, n38456, n38548, n41316, n38078, n38516, n38086,
    n38560, n38094, n42492, n38500, n39345, n39069, n39361, n38448, n39077,
    n39321, n39085, n39329, n39045, n39337, n38440, n39381, n28872, n38476,
    n36373, n39353, n39061, n39105, n38424, n37934, n28725, n39369, n38070,
    n39093, n36801, n39053, n38110, n37356, n37372, n38464, n28894, n41876,
    n38625, n27858, n39286, n42981, n42552, n28827, n37038, n37767, n37143,
    n40256, n43828, n43832, n36553, n43195, n28673, n38280, n41872, n37364,
    n36745, n38556, n42006, n44013, n38319, n38612, n43382, n37651, n38615,
    n39509, n37025, n41554, n39446, n26427, n36253, n44098, n28722, n38127,
    n36653, n39607, n26426, n39411, n26582, n37570, n37627, n24722, n41875,
    n26411, n28841, n37946, n43193, n42645, n42936, n37650, n37367, n42908,
    n43183, n38473, n39507, n43176, n43184, n26410, n28473, n34599, n26425,
    n43192, n26424, n43174, n40977, n39410, n26352, n26404, n43347, n43027,
    n35096, n34513, n41395, n40347, n34363, n41394, n38298, n35330, n26323,
    n39119, n25933, n25968, n43171, n37644, n28536, n24670, n24620, n25971,
    n39127, n35244, n34584, n26564, n42835, n26350, n34752, n28728, n26358,
    n26368, n40148, n27825, n25977, n42417, n38385, n41684, n42373, n24858,
    n38619, n42003, n42901, n33793, n43448, n28729, n40851, n34425, n24851,
    n28476, n27722, n26251, n26355, n24737, n41381, n25979, n41386, n42500,
    n38383, n24860, n40813, n38239, n25972, n26407, n25970, n35014, n41769,
    n22933, n38238, n42183, n26233, n26245, n27718, n41907, n37376, n40234,
    n40528, n25931, n41441, n37639, n28553, n40479, n37363, n28056, n28092,
    n41008, n41010, n42904, n42588, n33918, n27721, n40401, n41063, n40812,
    n37130, n41670, n41515, n40547, n41115, n36648, n40517, n40850, n35354,
    n41003, n39745, n39447, n41514, n40746, n26310, n42682, n26312, n42899,
    n41543, n24710, n24828, n26240, n27719, n41857, n24841, n35623, n35262,
    n39505, n27847, n40462, n27894, n41439, n40847, n40476, n42882, n42711,
    n32895, n32800, n24496, n40747, n36258, n42351, n27349, n42024, n24609,
    n41438, n38153, n32347, n40245, n32264, n39771, n41745, n27844, n40405,
    n26691, n39437, n39789, n39393, n26706, n26703, n32891, n41456, n35250,
    n23698, n42414, n37772, n40745, n37509, n26521, n26520, n40985, n42700,
    n36143, n37919, n32545, n41276, n41113, n40341, n41547, n40411, n41545,
    n27707, n42199, n26516, n41034, n32629, n42247, n39636, n42243, n43583,
    n23694, n34575, n40706, n42237, n35173, n40278, n36169, n43794, n28370,
    n40630, n28213, n28210, n38923, n24781, n34279, n41979, n43893, n25670,
    n40960, n41308, n40895, n37774, n40185, n35546, n40204, n42110, n41206,
    n39948, n38696, n43735, n39811, n38715, n43738, n43737, n43306, n40376,
    n38706, n36193, n43441, n36692, n40911, n24132, n43689, n23689, n36694,
    n36693, n36591, n36587, n36560, n36592, n36691, n32107, n36633, n34687,
    n36632, n39516, n36559, n36642, n25625, n36682, n36624, n35381, n36683,
    n36643, n36586, n40668, n36799, n36800, n40838, n36805, n36621, n36784,
    n37488, n36785, n36804, n36620, n43547, n41340, n41355, n36677, n36676,
    n40676, n36783, n43734, n39821, n36782, n43297, n36578, n39818, n42089,
    n26069, n26056, n36002, n40017, n40028, n40043, n39984, n39995, n40006,
    n39973, n39962, n36162, n35766, n32237, n43713, n24205, n40503, n23617,
    n39953, n34165, n35473, n34242, n42081, n25587, n34188, n25584, n41495,
    n41301, n34914, n43811, n43924, n26497, n40908, n40896, n27348, n40167,
    n24486, n24813, n34241, n43295, n31439, n41289, n39540, n40882, n32236,
    n39515, n26203, n41317, n24128, n32235, n26185, n28773, n34119, n34355,
    n37830, n28817, n34903, n37355, n41491, n36158, n24765, n37725, n40114,
    n36552, n26061, n36063, n23667, n39702, n31905, n37459, n36395, n24127,
    n35695, n35534, n39404, n36901, n26183, n23644, n24445, n36061, n36429,
    n36039, n23516, n24096, n24126, n28274, n28234, n28233, n28273, n28246,
    n27632, n35541, n28247, n26182, n28254, n28253, n28294, n27898, n27899,
    n26528, n28145, n28240, n26535, n28241, n26534, n31912, n41540, n27919,
    n27920, n26495, n36042, n26541, n28260, n26542, n28259, n28280, n28655,
    n28287, n27905, n27911, n28267, n26526, n39958, n25574, n26515, n24442,
    n42339, n24808, n27341, n27687, n41016, n40843, n36282, n35823, n40529,
    n34641, n26494, n33772, n24433, n40968, n31524, n31909, n23635, n32147,
    n25566, n34843, n31765, n32608, n28460, n42338, n36021, n28153, n32566,
    n31286, n41371, n32606, n32807, n34611, n35609, n25572, n41331, n25565,
    n26484, n36359, n27682, n23674, n32678, n26207, n26488, n28346, n28511,
    n28037, n23632, n28142, n25562, n27620, n23935, n23264, n32201, n32370,
    n25555, n31771, n27817, n31954, n26197, n23927, n41408, n23222, n24430,
    n24226, n27815, n32368, n27027, n32369, n28140, n27335, n23611, n23560,
    n32366, n31768, n23551, n23552, n32197, n24215, n27873, n32846, n32167,
    n23639, n28149, n24246, n25064, n26431, n32213, n25564, n26545, n31659,
    n27675, n41402, n26678, n28138, n37123, n32373, n23546, n26436, n25715,
    n26636, n26091, n41324, n25629, n27812, n28111, n36272, n25591, n31810,
    n25674, n41250, n37213, n25570, n23657, n25537, n32214, n24751, n37568,
    n25551, n35654, n43055, n24427, n23228, n25538, n23692, n23681, n27700,
    n26434, n25721, n23499, n27729, n27704, n25735, n25789, n25756, n26439,
    n23567, n27670, n26136, n25763, n32371, n23733, n23132, n25743, n27715,
    n23133, n28137, n38143, n25780, n26677, n24223, n25749, n26924, n23680,
    n27695, n35529, n23662, n28665, n25770, n23556, n23691, n25582, n27742,
    n23695, n23227, n42748, n27608, n25729, n31371, n25561, n24192, n31447,
    n24195, n24189, n25078, n25081, n27800, n25084, n24186, n25087, n25843,
    n31807, n25938, n25941, n23548, n41235, n24183, n24180, n25545, n31823,
    n24105, n27343, n27607, n23452, n26437, n27602, n23170, n41149, n24780,
    n23678, n23587, n23217, n25726, n25739, n25725, n24220, n25727, n25723,
    n25741, n23894, n23578, n23586, n25748, n25751, n25714, n25711, n25577,
    n26191, n27665, n41093, n25894, n23908, n24222, n25737, n24483, n27323,
    n23938, n26193, n23905, n24219, n25548, n25672, n25673, n25549, n25669,
    n23185, n24656, n24425, n27876, n40980, n26447, n27336, n23261, n23125,
    n25586, n26490, n25589, n25568, n25569, n27680, n28206, n25734, n25590,
    n25754, n41932, n25627, n25628, n25624, n25493, n43727, n27601, n26450,
    n36973, n25762, n23223, n25765, n25086, n25083, n25842, n23504, n23126,
    n23918, n25077, n23904, n25080, n24194, n24746, n27318, n24191, n24730,
    n26029, n32857, n24188, n35445, n23168, n24185, n25579, n25580, n24130,
    n27333, n28051, n28048, n26909, n27035, n27032, n26686, n31451, n25533,
    n25534, n27673, n26683, n25719, n25718, n27605, n27328, n26143, n42745,
    n26034, n25940, n25937, n24199, n24329, n33357, n24179, n24176, n24411,
    n24182, n27795, n24170, n24732, n26505, n25109, n31716, n25833, n24908,
    n25585, n31056, n25059, n24983, n27249, n24946, n24729, n24118, n24405,
    n23851, n31921, n24607, n25093, n24232, n23917, n23910, n23085, n38909,
    n23909, n27747, n31448, n24745, n23896, n26223, n27792, n24856, n24846,
    n24836, n24834, n25995, n27614, n25494, n25575, n26328, n23501, n26177,
    n36561, n25062, n27613, n27611, n35976, n27610, n35425, n26282, n27627,
    n24208, n24728, n24866, n27671, n24659, n24169, n26428, n24109, n27248,
    n31803, n25710, n23052, n24099, n34645, n27320, n27660, n26440, n25021,
    n28810, n33486, n27788, n27805, n27595, n31805, n36546, n27591, n23083,
    n35963, n27656, n25837, n24985, n24733, n23486, n23414, n23446, n24391,
    n34164, n40038, n39981, n39989, n40011, n39967, n23277, n39939, n39970,
    n40000, n40014, n40022, n40025, n39992, n40033, n40003, n40049, n39978,
    n23485, n23442, n27380, n27379, n27440, n23370, n27079, n24948, n23080,
    n27559, n23402, n23049, n24489, n23338, n24488, n27410, n27314, n23936,
    n23944, n27529, n25061, n23406, n23027, n23336, n23351, n23078, n23361,
    n23238, n23061, n23301, n23310, n23413, n23487, n31189, n27226, n27227,
    n24910, n25020, n25619, n25612, n27409, n23963, n23977, n24089, n27770,
    n27446, n27452, n23768, n27244, n23655, n24602, n24687, n24686, n23962,
    n23376, n24058, n24037, n23438, n23059, n23369, n23025, n23359, n23028,
    n23832, n23968, n23401, n23391, n23480, n23976, n23873, n23872, n23076,
    n24067, n24080, n23345, n23043, n23316, n23062, n24383, n23334, n23459,
    n23421, n23955, n23954, n23317, n23412, n23823, n27185, n23831, n27538,
    n27166, n23969, n23884, n23951, n24063, n23033, n27368, n23885, n23411,
    n23344, n23042, n24059, n23974, n27104, n27546, n27051, n23767, n23870,
    n27269, n23975, n23861, n23824, n27115, n24036, n27221, n27492, n24596,
    n24595, n24601, n27478, n27465, n39896, n23375, n27387, n24587, n27420,
    n23067, n27418, n23075, n23068, n27760, n24361, n27451, n23312, n23437,
    n24440, n27508, n23837, n27518, n23210, n23838, n27358, n27562, n27572,
    n27564, n23435, n27434, n27477, n24251, n27433, n23366, n27073, n25687,
    n27480, n27426, n23903, n23363, n27472, n27488, n27487, n23371, n27491,
    n26820, n23298, n24229, n23117, n27251, n27258, n27260, n23477, n27137,
    n23184, n38059, n22925, n27411, n23073, n23071, n24453, n27081, n31825,
    n27273, n32880, n23340, n27523, n36363, n27353, n27359, n23860, n23871,
    n27548, n27547, n27552, n27553, n24084, n27503, n23970, n23971, n27583,
    n27561, n27584, n27582, n23409, n27577, n23964, n23957, n23037, n27389,
    n27145, n23040, n24083, n27570, n23972, n27569, n27397, n23830, n24082,
    n27510, n27199, n43729, n27232, n27231, n32867, n23296, n23374, n23365,
    n35804, n23041, n34515, n41310, n41560, n24838, n22905, n23182, n23074,
    n27188, n27183, n27256, n23891, n27118, n23829, n22907, n23877, n27101,
    n29305, n27096, n28494, n27748, n31495, n22908, n24506, n43499, n23275,
    n29439, n22927, n23077, n24833, n22912, n27061, n27539, n36316, n24510,
    n29553, n24825, n24438, n39310, n24228, n23631, n44099, n27431, n29721,
    n27479, n23608, n26862, n23570, n23943, n23942, n35630, n23932, n25114,
    n27757, n24864, n26877, n43496, n23183, n23720, n27058, n36311, n40127,
    n35811, n36366, n31488, n26174, n24436, n42011, n24504, n24248, n35802,
    n37023, n27182, n27181, n36364, n24842, n23039, n24829, n34550, n31507,
    n41671, n33842, n40196, n31667, n40998, n27117, n26099, n29726, n28755,
    n34476, n29997, n41341, n29171, n27153, n31953, n33734, n36307, n23665,
    n23634, n42746, n42747, n34726, n43864, n43905, n43898, n43795, n43728,
    n32238, n27070, n36295, n23724, n36306, n34576, n22920, n22921, n22922,
    n40306, n36299, n26235, n22924, n23019, n23571, n24743, n24406, n24508,
    n24115, n24426, n23583, n23566, n23603, n42197, n27860, n23709, n23708,
    n27689, n42002, n25936, n42285, n42066, n40395, n27668, n41332, n43379,
    n25076, n37000, n35821, n43016, n39671, n42872, n38016, n37839, n34906,
    n36625, n36579, n24631, n24630, n24633, n24624, n24625, n24626, n24640,
    n24641, n24639, n24679, n24678, n24677, n24599, n24600, n24598, n24591,
    n24592, n24594, n24585, n24586, n24583, n23172, n25615, n25614, n25616,
    n25611, n25595, n23191, n23190, n23204, n23092, n23091, n23096, n23097,
    n23108, n23110, n23897, n27003, n27010, n24717, n24576, n23853, n23857,
    n25285, n25635, n25636, n23245, n23232, n23235, n27228, n27537, n27533,
    n27462, n27464, n27457, n27458, n27456, n27443, n24726, n24027, n24735,
    n35325, n24133, n24333, n24296, n24485, n31891, n24015, n33720, n33719,
    n33717, n23591, n43099, n25559, n28284, n42204, n42094, n42084, n38945,
    n26499, n26496, n23534, n23321, n23490, n23383, n26167, n23124, n35771,
    n35772, n27388, n27384, n27383, n27381, n27765, n27521, n27516, n27501,
    n27502, n27413, n27414, n27594, n27374, n27373, n40823, n39773, n41349,
    n41348, n24171, n26634, n26600, n24874, n25023, n37500, n24848, n34344,
    n40079, n42483, n41435, n26146, n26715, n26142, n25984, n25841, n37219,
    n36905, n23888, n24388, n24443, n24503, n24117, n31903, n23979, n33716,
    n34505, n23510, n23220, n26195, n28277, n42256, n40282, n39461, n37329,
    n28271, n25222, n25234, n25159, n25160, n25162, n25174, n25169, n42749,
    n43829, n43613, n28309, n37466, n28282, n42202, n23729, n23500, n23714,
    n26209, n37796, n42782, n39525, n39528, n27255, n40861, n27347, n27677,
    n27317, n39788, n40412, n40210, n39401, n27685, n40269, n38594, n43374,
    n28820, n28044, n28512, n26680, n28485, n26138, n25850, n36900, n37220,
    n34814, n41898, n25992, n37536, n31908, n43571, n28854, n28505, n26581,
    n25975, n38798, n37551, n43359, n43135, n42551, n28723, n42815, n42833,
    n42680, n41127, n37498, n35237, n38406, n28196, n40932, n37729, n37727,
    n37728, n23663, n23605, n41657, n41565, n36377, n42219, n35380, n42564,
    n43667, n43224, n42857, n42516, n42515, n42437, n42288, n42526, n42612,
    n42611, n42259, n42632, n42111, n42139, n36613, n36846, n27100, n39445,
    n28091, n40241, n40239, n40253, n40331, n40229, n40963, n40972, n41537,
    n40374, n39631, n43575, n28879, n28533, n42180, n37520, n36115, n35887,
    n36149, n35512, n42941, n28660, n28465, n26693, n26713, n26717, n26150,
    n26033, n26038, n41454, n41024, n40707, n39593, n43029, n42679, n41968,
    n40784, n26585, n38659, n40795, n40793, n26572, n40099, n24757, n24756,
    n35836, n39765, n39754, n39704, n42439, n36393, n38956, n39715, n39295,
    n42637, n42424, n38980, n38970, n25796, n38015, n40152, n42514, n42138,
    n39667, n37626, n37602, n37527, n37914, n37906, n37545, n37430, n37412,
    n37421, n37404, n38936, n38623, n40914, n40902, n40889, n41299, n41298,
    n41319, n41287, n41286, n35941, n40810, n36401, n41398, n41414, n37776,
    n38167, n38168, n38029, n37593, n40958, n40983, n40994, n40993, n40992,
    n38589, n38609, n41372, n26398, n26393, n26397, n26392, n25605, n26346,
    n28586, n26100, n24646, n24647, n24644, n24645, n24632, n24627, n24638,
    n24685, n24684, n24682, n24683, n24701, n24700, n24694, n24695, n24676,
    n24355, n24364, n24368, n24378, n24367, n24356, n26094, n24267, n24255,
    n23131, n23174, n43085, n26260, n26405, n26345, n23289, n23313, n23355,
    n23890, n23933, n23930, n26096, n28616, n23761, n23757, n23762, n43251,
    n43245, n43265, n24578, n24577, n24580, n24579, n24597, n24593, n24584,
    n24613, n24345, n24363, n23862, n23867, n23866, n23863, n28592, n24210,
    n24373, n24341, n24377, n24352, n24342, n24346, n24374, n24264, n24275,
    n43260, n43261, n43274, n43264, n43241, n43242, n40587, n28202, n26301,
    n25676, n43086, n41805, n26790, n26768, n41588, n26396, n25657, n25658,
    n25660, n25617, n25613, n25599, n42787, n26232, n25517, n25518, n25506,
    n25507, n25508, n43172, n28201, n25697, n23198, n23199, n23193, n23208,
    n23089, n23098, n23112, n41631, n26298, n23128, n23181, n27761, n27600,
    n27603, n27339, n27551, n27554, n27563, n27568, n27473, n27493, n27494,
    n23898, n24098, n43239, n24053, n24049, n24048, n24052, n24043, n24038,
    n24042, n24021, n24022, n24017, n27971, n26978, n26944, n23752, n23749,
    n25926, n25927, n25896, n24978, n24982, n24941, n24945, n24903, n24904,
    n24907, n24859, n24845, n24823, n43456, n24718, n24418, n24137, n23852,
    n23856, n24387, n24734, n24238, n24242, n24233, n24480, n34682, n33709,
    n23266, n23493, n23224, n28203, n42209, n28200, n26444, n23136, n26460,
    n28211, n43426, n25241, n25257, n25258, n26257, n25167, n41602, n41598,
    n43092, n41592, n26819, n25768, n25761, n25202, n25181, n25182, n25187,
    n25188, n25196, n25120, n25121, n25140, n25139, n25664, n25663, n25632,
    n23247, n23234, n25492, n25524, n25523, n26271, n23155, n43659, n28291,
    n42099, n27885, n23723, n25685, n25686, n25703, n25681, n26391, n26390,
    n26476, n23547, n26286, n23169, n23458, n25692, n23468, n26157, n23130,
    n26159, n27768, n27417, n27049, n34767, n33298, n27158, n27151, n27154,
    n27157, n27146, n34766, n27710, n27345, n27366, n27365, n27367, n27357,
    n27360, n28747, n42323, n27229, n27684, n27327, n27667, n27672, n27798,
    n32198, n27545, n27540, n27531, n27447, n27449, n27466, n27463, n27459,
    n27444, n27578, n27485, n27486, n41330, n26676, n26134, n25943, n24853,
    n24854, n24791, n24031, n24028, n26977, n28478, n25836, n25019, n24798,
    n24797, n40072, n28720, n28719, n28669, n28668, n28832, n28663, n28522,
    n28466, n28054, n28052, n28523, n28550, n28049, n28047, n27036, n41436,
    n27033, n26689, n26687, n41437, n26714, n26141, n25983, n25935, n25840,
    n37532, n37531, n24753, n24725, n24740, n34817, n24173, n32549, n34058,
    n24494, n24157, n26568, n31916, n24103, n24108, n32131, n32116, n24125,
    n24121, n34691, n34685, n38403, n38492, n38484, n38490, n39316, n38063,
    n34684, n34508, n23507, n43668, n43607, n39764, n37274, n36385, n25746,
    n25747, n40355, n26446, n38821, n39569, n43512, n43503, n28264, n28257,
    n25327, n25328, n25281, n25295, n23592, n23630, n28186, n40921, n41564,
    n26923, n25788, n25784, n25487, n25732, n25733, n26384, n25558, n25491,
    n28139, n28136, n28134, n35971, n28127, n28124, n28125, n23163, n23149,
    n23150, n23144, n23143, n43753, n28353, n41940, n28336, n28329, n28330,
    n43584, n28321, n28314, n28307, n28305, n28300, n28298, n28292, n26919,
    n42713, n28285, n42716, n42347, n42348, n42283, n25779, n42279, n42253,
    n42257, n25775, n42387, n42245, n26503, n26500, n42382, n36840, n25544,
    n36489, n36486, n23645, n32944, n32945, n25547, n41474, n34879, n23537,
    n23538, n43091, n37620, n38237, n38329, n37139, n36746, n37870, n24777,
    n38626, n37951, n36635, n37362, n26172, n26171, n23568, n35777, n27396,
    n27398, n27390, n27382, n27402, n27790, n27804, n27774, n31665, n35641,
    n33741, n36164, n35408, n35420, n33620, n27507, n27509, n27524, n27515,
    n27504, n27428, n27425, n27412, n36310, n36298, n27187, n27797, n38905,
    n32883, n39450, n40726, n27321, n27663, n36664, n27319, n35446, n27352,
    n27351, n27372, n41407, n28745, n40997, n37765, n39449, n39774, n40215,
    n40213, n40211, n35861, n27690, n36075, n35988, n36020, n40194, n27809,
    n27784, n29841, n33502, n36294, n41337, n41351, n42160, n28661, n28469,
    n42412, n42404, n42184, n41848, n27843, n27841, n26702, n27836, n40703,
    n37241, n34823, n36990, n26065, n39942, n28656, n28461, n27026, n25849,
    n33791, n31794, n31697, n25071, n28858, n28735, n42173, n26633, n26028,
    n37242, n31360, n31359, n43712, n43558, n43138, n43046, n43378, n28860,
    n43035, n28737, n28731, n42410, n42174, n42507, n42498, n41899, n41955,
    n41444, n41196, n41025, n40708, n26578, n41131, n40490, n38389, n39592,
    n38804, n36269, n24812, n43442, n43569, n43042, n42817, n42935, n42934,
    n43329, n42834, n42172, n41743, n43330, n26148, n41022, n40798, n40797,
    n26571, n40098, n38662, n38643, n35822, n36264, n35682, n34339, n34818,
    n35334, n33309, n33792, n36893, n32532, n24339, n39301, n34725, n33718,
    n34258, n35180, n34748, n34421, n35351, n34090, n34088, n35089, n35033,
    n33726, n44106, n29579, n23509, n26199, n27871, n43524, n41936, n41728,
    n43175, n42721, n42467, n28278, n40570, n41783, n41265, n37831, n28269,
    n28272, n35964, n36203, n35598, n28227, n25233, n35426, n34918, n25176,
    n25173, n35253, n36248, n43056, n43389, n43672, n41211, n42799, n42909,
    n40053, n38014, n37121, n41703, n32217, n43777, n28141, n42354, n42215,
    n42658, n42140, n42561, n41702, n26519, n33563, n43842, n43891, n43743,
    n43814, n43682, n43661, n43645, n43315, n43316, n43317, n43155, n43154,
    n43582, n43581, n43537, n39761, n43549, n43223, n43211, n42953, n42952,
    n42906, n42992, n43015, n43018, n43014, n42998, n42855, n42722, n42871,
    n42874, n42870, n42598, n42628, n42224, n42423, n42212, n42668, n42841,
    n42451, n28076, n41171, n27854, n42600, n39656, n25576, n26546, n36612,
    n35790, n43164, n26211, n26210, n36500, n37945, n32893, n32894, n32509,
    n37625, n37624, n37641, n37640, n38331, n38330, n39125, n37858, n37857,
    n38212, n37947, n38294, n38297, n38614, n37953, n37952, n36634, n37360,
    n37359, n37373, n39526, n41284, n32966, n36161, n41518, n34656, n32858,
    n32859, n33124, n33622, n33514, n41389, n32253, n32472, n34011, n35307,
    n32826, n32284, n27315, n41399, n41091, n40859, n41156, n40732, n41100,
    n41233, n40817, n40410, n40335, n36869, n32881, n36195, n36439, n36433,
    n36444, n36446, n40371, n36927, n36913, n36659, n27282, n27653, n27654,
    n41535, n41556, n40836, n41011, n39796, n40532, n40466, n40425, n40408,
    n39444, n39412, n39409, n41240, n40398, n40981, n40200, n27593, n40182,
    n40179, n38605, n27810, n27786, n43990, n41354, n36055, n36052, n42016,
    n42013, n31442, n43800, n43384, n42166, n43343, n41854, n41904, n26708,
    n40718, n40715, n41140, n26078, n26081, n38792, n37519, n37507, n43570,
    n35515, n43796, n28046, n40493, n38636, n44007, n37550, n34815, n42028,
    n41425, n41039, n40549, n41130, n32233, n44092, n31748, n31757, n42371,
    n28497, n28549, n28483, n41742, n40802, n40692, n40486, n39643, n39594,
    n37516, n37501, n37502, n37243, n37003, n37002, n36993, n35681, n36110,
    n35518, n42829, n41749, n41279, n41278, n40805, n40804, n25986, n25985,
    n39563, n24203, n32340, n39964, n39975, n40008, n39997, n39986, n40045,
    n40030, n40019, n39076, n39068, n39084, n39044, n39052, n39060, n39104,
    n39092, n38446, n38447, n38438, n38439, n38474, n38475, n38462, n38463,
    n38422, n38423, n38430, n38431, n38414, n38415, n38454, n38455, n38531,
    n38523, n38539, n38507, n38547, n38515, n38559, n38499, n34730, n39328,
    n39360, n39344, n39336, n39352, n39368, n39380, n39320, n38108, n38109,
    n38068, n38069, n38100, n38101, n38116, n38117, n38084, n38085, n38092,
    n38093, n38076, n38077, n38128, n38129, n39873, n39865, n39833, n39885,
    n39825, n39849, n39857, n39841, n38855, n38863, n38847, n38839, n38891,
    n38879, n38871, n29568, n44000, n28151, n29550, n41916, n28148, n28222,
    n41737, n40933, n37470, n37461, n37275, n37267, n42352, n37731, n37730,
    n40687, n42452, n40663, n39491, n39470, n37338, n40367, n38833, n40579,
    n40324, n28368, n43633, n41755, n26911, n40069, n42616, n42842, n42565,
    n35599, n34917, n40580, n40325, n43130, n41842, n41675, n40067, n40298,
    n25097, n36958, n36957, n36011, n31353, n43912, n43808, n43013, n42709,
    n42431, n42059, n42076, n41170, n38379, n38377, n37556, n36493, n36492,
    n43812, n43754, n43776, n43775, n43644, n43578, n43156, n43222, n42894,
    n42520, n42519, n42868, n42282, n42289, n42560, n41697, n40941, n40758,
    n28061, n40769, n39651, n36862, n36616, n36615, n34913, n36532, n37782,
    n37739, n37799, n37840, n37817, n37790, n37809, n36940, n36680, n37596,
    n37648, n37939, n38567, n38565, n38357, n38356, n38341, n38340, n38349,
    n38348, n38581, n38575, n38573, n38365, n38364, n37150, n37209, n37198,
    n37174, n37158, n37182, n37166, n37190, n39147, n39173, n39165, n39139,
    n39157, n39181, n39194, n37048, n37081, n37064, n37072, n37056, n39203,
    n38709, n38718, n38672, n38681, n38690, n38929, n38699, n37976, n37957,
    n38008, n37992, n38000, n38304, n37984, n36729, n36808, n36788, n36705,
    n36697, n36796, n36713, n37368, n37392, n37384, n38769, n41314, n38814,
    n29204, n29221, n41365, n36168, n35644, n34545, n33756, n35525, n41864,
    n41681, n41863, n34400, n43933, n42135, n41059, n36281, n33062, n32501,
    n33095, n32193, n43984, n41532, n41118, n41111, n40848, n40815, n37024,
    n36868, n36479, n36963, n36978, n41259, n41002, n40254, n40531, n40484,
    n40431, n40421, n40344, n40231, n40146, n40142, n40973, n40515, n40459,
    n39633, n39620, n40191, n38731, n36352, n40418, n29449, n43992, n43577,
    n28896, n28880, n28845, n28844, n28538, n42191, n27851, n36116, n35891,
    n36150, n28826, n28724, n28672, n41442, n26694, n26718, n26151, n26039,
    n25948, n37537, n43741, n39936, n37825, n43365, n43141, n42820, n43038,
    n42510, n41958, n38396, n35687, n42988, n42556, n26575, n35838, n37494,
    n34524, n34522, n39929, n39770, n40119, n39708, n36398, n39228, n40641,
    n40598, n40618, n39583, n39716, n39296, n39297, n38138, n38139, n38982,
    n38028, n33424, n33428, n33432, n33436, n33440, n33444, n33448, n33452,
    n33456, n33460, n33477, n33464, n33468, n33472, n43909, n42479, n42446,
    n42268, n42396, n42149, n40164, n42125, n39668, n37605, n37529, n37917,
    n37909, n39613, n37549, n37433, n37414, n37424, n37406, n38939, n38635,
    n38314, n38275, n38751, n38743, n38779, n38759, n38767, n40916, n40904,
    n40892, n40893, n41306, n41294, n35781, n35958, n35660, n40546, n39744,
    n39504, n37922, n37327, n36405, n36179, n35555, n41421, n41167, n39438,
    n37778, n37777, n38169, n38189, n37594, n38048, n36887, n36673, n27820,
    n28105, n28771, n40986, n38610, n42026, n27152, n28191, n22929, n22930,
    n22931, n22932, n43540, n23127, n22934, n34812, n22935, n22936, n22937,
    n27697, n34858, n26859, n28062, n26522, n28316, n22938, n22939, n22940,
    n22941, n23758, n27696, n22942, n25556, n25758, n26849, n28236, n24862,
    n28249, n29669, n28229, n28331, n25724, n22943, n35543, n33191, n24804,
    n28345, n26537, n27915, n29493, n29749, n24818, n24788, n29506, n28324,
    n23636, n28262, n27901, n26530, n25671, n25738, n29462, n22945, n28289,
    n43850, n25583, n24283, n24537, n23225, n26302, n24287, n24351, n24665,
    n38489, n25644, n27625, n24039, n24018, n24432, n42783, n26806, n23618,
    n27094, n28648, n24435, n24565, n24335, n40672, n23467, n43833, n26479,
    n39772, n24422, n28354, n28302, n42754, n25626, n42465, n26283, n27301,
    n26179, n40312, n42206, n26486, n43660, n42096, n35439, n26063, n42546,
    n35366, n42801, n37271, n42657, n41173, n43605, n42255, n27867, n36562,
    n38325, n37374, n35711, n37577, n40441, n25065, n41191, n26570, n34679,
    n26910, n43539, n28123, n36918, n40748, n37694, n36661, n30837, n28928,
    n26046, n32136, n28822, n37846, n31989, n34243, n43351, n40089, n39710,
    n41785, n38969, n43390, n32271, n31252, n28144, n27852, n37286, n43599,
    n42303, n39600, n29471, n39502, n41391, n34402, n33527, n31633, n32499,
    n34844, n36220, n40820, n38732, n36966, n29381, n44105, n39741, n35551,
    n43931, n36283, n43967, n22981, n36557, n27891, n32176, n31487, n35800,
    n23018, n23541, n23021, n23045, n35718, n23036, n23464, n23035, n25645,
    n26832, n25652, n23051, n23044, n25656, n26726, n23047, n26878, n23048,
    n23050, n23055, n23070, n23069, n23084, n23082, n26828, n23079, n23081,
    n23088, n26789, n23086, n23087, n23090, n25495, n23095, n25440, n23107,
    n26808, n23106, n23111, n25641, n23114, n23115, n23129, n26154, n39534,
    n23138, n23137, n23140, n23139, n23142, n23141, n23146, n23145, n23148,
    n23147, n23153, n23157, n23154, n23159, n23158, n23160, n23162, n34885,
    n23171, n23267, n26317, n23187, n23186, n23189, n23188, n23195, n23194,
    n23197, n23196, n23203, n23202, n23207, n23206, n23211, n23564, n23281,
    n23231, n23229, n23230, n26780, n26737, n23244, n23242, n23243, n26341,
    n23270, n23282, n23274, n23276, n26168, n23280, n23285, n23512, n23288,
    n23286, n26192, n23287, n31493, n25653, n23291, n23295, n23292, n23294,
    n23297, n23299, n23302, n23308, n23307, n23309, n23319, n23311, n23315,
    n23314, n23320, n23322, n23339, n23330, n23352, n23342, n23347, n23349,
    n23348, n23350, n36779, n23385, n23354, n23372, n23373, n23382, n23378,
    n23380, n23379, n23381, n23448, n23387, n23404, n23417, n23444, n23440,
    n23441, n23443, n36688, n26184, n23585, n23450, n23451, n23544, n23454,
    n23489, n23483, n23484, n23488, n23520, n23495, n23494, n23496, n26200,
    n23498, n23502, n23505, n23711, n23730, n23706, n31058, n23506, n23508,
    n31770, n25099, n32148, n31057, n29085, n23518, n23517, n31819, n23532,
    n23519, n23521, n23522, n23527, n23562, n23554, n23525, n23526, n23530,
    n23553, n23528, n23529, n23533, n31766, n28197, n23535, n23536, n23701,
    n23550, n23555, n23715, n23557, n25096, n23702, n23593, n23561, n23574,
    n25532, n23563, n23731, n23569, n35707, n23572, n23573, n23582, n23598,
    n23580, n23590, n41873, n23584, n23659, n23610, n27912, n23589, n23614,
    n23597, n39573, n23601, n23599, n23602, n23604, n26527, n23606, n23675,
    n23612, n23609, n23676, n23616, n23623, n23633, n23666, n26512, n23625,
    n23624, n23627, n26518, n23646, n23643, n28361, n23640, n23638, n23641,
    n26513, n23650, n23648, n23651, n36607, n38820, n31816, n23658, n23685,
    n23653, n39508, n42796, n25105, n25107, n23699, n23668, n23669, n23672,
    n23677, n23683, n23682, n23690, n32143, n37852, n32892, n32896, n25106,
    n36533, n23744, n23710, n23704, n23705, n23707, n23713, n23712, n31522,
    n26506, n35750, n23742, n23718, n35725, n35721, n23721, n23740, n26509,
    n23725, n35722, n43484, n23726, n23727, n23738, n26508, n23732, n23734,
    n35752, n23736, n35729, n23735, n23737, n23739, n23741, n35714, n23743,
    n23745, n23747, n23746, n35113, n23748, n35112, n34283, n35099, n25950,
    n33721, n23772, n24795, n24515, n31922, n24517, n32084, n32118, n32121,
    n23769, n24539, n26095, n24526, n24527, n23788, n27006, n23771, n31937,
    n28585, n23770, n27004, n23774, n28591, n23773, n27011, n23779, n26659,
    n23778, n28593, n27009, n23780, n23786, n39891, n23790, n23789, n23794,
    n23793, n23802, n23795, n23800, n23798, n23797, n23799, n23801, n23818,
    n23804, n23803, n23808, n23806, n23807, n23816, n23812, n23813, n23817,
    n31382, n23847, n23834, n43270, n23833, n23836, n23835, n23840, n23839,
    n23842, n23841, n23845, n23875, n23874, n43271, n23876, n23887, n23881,
    n23883, n23882, n23886, n24122, n23895, n24394, n24872, n23945, n24655,
    n23923, n23906, n24200, n23907, n35466, n23941, n23940, n23939, n23947,
    n24101, n23949, n23948, n23950, n23952, n23967, n23966, n23973, n23978,
    n24002, n24001, n24004, n24003, n24014, n24008, n24007, n24012, n24010,
    n24009, n24011, n24013, n24061, n24060, n24092, n25069, n24062, n24091,
    n24090, n24093, n31478, n39895, n24094, n24107, n31374, n24104, n24106,
    n32239, n24149, n24110, n24113, n24120, n24134, n24123, n24124, n31715,
    n24509, n44102, n35474, n31892, n24131, n32080, n42922, n24148, n31477,
    n24136, n24240, n40073, n28825, n24235, n24138, n24206, n24146, n24144,
    n24140, n24141, n24143, n24145, n24147, n24151, n25068, n32123, n24152,
    n42924, n24154, n36891, n24420, n32540, n34290, n35100, n25952, n24153,
    n24155, n24752, n24738, n25951, n24156, n24762, n24158, n39315, n32552,
    n24160, n24159, n35833, n24760, n32232, n24163, n31358, n24164, n43344,
    n31705, n37246, n24758, n24198, n24197, n24202, n24201, n31449, n36906,
    n24213, n31898, n24424, n24212, n24217, n24727, n24218, n24241, n24231,
    n24224, n24225, n24230, n24338, n31936, n24429, n24253, n24298, n24477,
    n24254, n24257, n24256, n24258, n24260, n24259, n24263, n24266, n24265,
    n24269, n24268, n24274, n24277, n24276, n24279, n24278, n24282, n24285,
    n24284, n24286, n24289, n24288, n24749, n24399, n24390, n24344, n24343,
    n24350, n24348, n24347, n24349, n24354, n24353, n24360, n24358, n24357,
    n24359, n24366, n24365, n24372, n24370, n24369, n24371, n24376, n24375,
    n24382, n24380, n24379, n24381, n24412, n24397, n24398, n25895, n24400,
    n24403, n24402, n24484, n34560, n24410, n24404, n24408, n24407, n24409,
    n24416, n34551, n24415, n24413, n24491, n24414, n31687, n24417, n32062,
    n32556, n32061, n24421, n24495, n24423, n32546, n24428, n35165, n24446,
    n36136, n24563, n24478, n24499, n24487, n24497, n24564, n24490, n24492,
    n24493, n32547, n34057, n24498, n24502, n24513, n24514, n24519, n24516,
    n24518, n24520, n24522, n24521, n24525, n24529, n24528, n26662, n24532,
    n24530, n24531, n24541, n24538, n24540, n24542, n24544, n28590, n24543,
    n24547, n24549, n28584, n24548, n26658, n24552, n24550, n24551, n24561,
    n24573, n24569, n24566, n24567, n24571, n24570, n24572, n35322, n34055,
    n24574, n24622, n24616, n24617, n35332, n24619, n24621, n24674, n24664,
    n24712, n24668, n24661, n24663, n24660, n24662, n24666, n24667, n24669,
    n36128, n24671, n24675, n36086, n24673, n36091, n35109, n24691, n24690,
    n24693, n24692, n24697, n24696, n24699, n24698, n24714, n24719, n35104,
    n24724, n35108, n35110, n35831, n24747, n24736, n24744, n25962, n24748,
    n24750, n24755, n43469, n37006, n24764, n24763, n37285, n24767, n28146,
    n28122, n28118, n24769, n24768, n24774, n36365, n24770, n35756, n35751,
    n24772, n24771, n35749, n24773, n24783, n24776, n24782, n24784, n24786,
    n24785, n24873, n43722, n24815, n24792, n24790, n43294, n36144, n24789,
    n32630, n24799, n24796, n24806, n24805, n24809, n24810, n32631, n33313,
    n24827, n35889, n43725, n24821, n24819, n24820, n33314, n33794, n24832,
    n24850, n24844, n35820, n36992, n24868, n24863, n24865, n24870, n36273,
    n24876, n24875, n24880, n24878, n24877, n24879, n24888, n24882, n24881,
    n24886, n24884, n24883, n24885, n24887, n24890, n24889, n24894, n24892,
    n24891, n24893, n24902, n24896, n24895, n24900, n24898, n24897, n24899,
    n24901, n24912, n24914, n24913, n24918, n24916, n24915, n24917, n24926,
    n24920, n24919, n24924, n24922, n24921, n24923, n24925, n24942, n24928,
    n24927, n24932, n24930, n24929, n24931, n24940, n24934, n24933, n24938,
    n24936, n24935, n24937, n24939, n24951, n24950, n24955, n24953, n24952,
    n24954, n24963, n24957, n24956, n24961, n24959, n24958, n24960, n24962,
    n24979, n24965, n24964, n24969, n24967, n24966, n24968, n24977, n24971,
    n24970, n24975, n24973, n24972, n24974, n24976, n24987, n24989, n24988,
    n24993, n24991, n24990, n24992, n25001, n24995, n24994, n24999, n24997,
    n24996, n24998, n25000, n25017, n25003, n25002, n25007, n25005, n25004,
    n25006, n25015, n25009, n25008, n25013, n25011, n25010, n25012, n25014,
    n25016, n25018, n25028, n25027, n25032, n25030, n25029, n25031, n25040,
    n25034, n25033, n25038, n25036, n25035, n25037, n25039, n25056, n25042,
    n25041, n25046, n25044, n25043, n25045, n25054, n25048, n25047, n25052,
    n25050, n25049, n25051, n25053, n25055, n25057, n25058, n25067, n25070,
    n31904, n25075, n35626, n43300, n43298, n25090, n25089, n25091, n25095,
    n25098, n25100, n41759, n25101, n25104, n43690, n25103, n25800, n25112,
    n25108, n25111, n25117, n25116, n25119, n25118, n25123, n25122, n25127,
    n25125, n25124, n25126, n25377, n25132, n25130, n25131, n25136, n25134,
    n25133, n25135, n25138, n25137, n26891, n25142, n25360, n25141, n25717,
    n34646, n25150, n25148, n25147, n25149, n25154, n25152, n25151, n25153,
    n25156, n25155, n25158, n25157, n25164, n25499, n25163, n25170, n25168,
    n25166, n25165, n25172, n25171, n25178, n25177, n25180, n25179, n25184,
    n25183, n25186, n25185, n25424, n25192, n25191, n25194, n25193, n41648,
    n25195, n25198, n25197, n25200, n25199, n25201, n25731, n41804, n25208,
    n25469, n25207, n25214, n41822, n25212, n25210, n25209, n25211, n25213,
    n25216, n25215, n25220, n25218, n25217, n25219, n25221, n25224, n25223,
    n25226, n25225, n25230, n25228, n25227, n25229, n25232, n25231, n25238,
    n25237, n25242, n25240, n25239, n25244, n25243, n25248, n25246, n25245,
    n25247, n25252, n25251, n25254, n25253, n25256, n25255, n25260, n25259,
    n25262, n25261, n25263, n25745, n25268, n25267, n25272, n25270, n25269,
    n25271, n25282, n25274, n25273, n25280, n25276, n25275, n25278, n25277,
    n25279, n25284, n25283, n25291, n25289, n25287, n25286, n25288, n25290,
    n25293, n25292, n25294, n25299, n25298, n25303, n25301, n25300, n25302,
    n25311, n25305, n25304, n25309, n25307, n25306, n25308, n25310, n43425,
    n25314, n25312, n25313, n25316, n25315, n25320, n25318, n25317, n25319,
    n25326, n25324, n25322, n25321, n25323, n25325, n25759, n25330, n25329,
    n25334, n25332, n25331, n25333, n25344, n25336, n25335, n25338, n25337,
    n25342, n25340, n25339, n25341, n25343, n25359, n25345, n25349, n25347,
    n25346, n25348, n25353, n25351, n25350, n25352, n25357, n25355, n25354,
    n25356, n25358, n25362, n25361, n25364, n25363, n25368, n25366, n25365,
    n25367, n25376, n25370, n25369, n25374, n25372, n25371, n25373, n25375,
    n25391, n25379, n25378, n25381, n25380, n25385, n25383, n25382, n25384,
    n25389, n25387, n25386, n25388, n25390, n37442, n25393, n25392, n25397,
    n25395, n25394, n25396, n25405, n25399, n25398, n25403, n25401, n25400,
    n25402, n25404, n25421, n41601, n25407, n25406, n25411, n41591, n25409,
    n25408, n25410, n25415, n25413, n25412, n25414, n25419, n25417, n25416,
    n25418, n25420, n37441, n25423, n25422, n25430, n25426, n25425, n25428,
    n25427, n25429, n25438, n25432, n25431, n25436, n25434, n25433, n25435,
    n25437, n25454, n25439, n25442, n25441, n25444, n25443, n25448, n25446,
    n25445, n25447, n25452, n25450, n25449, n25451, n25453, n25456, n25455,
    n25460, n25458, n25457, n25459, n25468, n25462, n25461, n25466, n25464,
    n25463, n25465, n25467, n25486, n25471, n25470, n25475, n25473, n41821,
    n25472, n25474, n25479, n25477, n25476, n25478, n25484, n26288, n25482,
    n25480, n25481, n25483, n25485, n25488, n25489, n41754, n25497, n25496,
    n25498, n25501, n25500, n25505, n25504, n25514, n25516, n25515, n25520,
    n25531, n25550, n25536, n25553, n32168, n25542, n26914, n41473, n32890,
    n25567, n36831, n25588, n25594, n25593, n25598, n25597, n25602, n25601,
    n25607, n43072, n25606, n25609, n25608, n25610, n36829, n25633, n25631,
    n25638, n25643, n43409, n25642, n25647, n26817, n25646, n25655, n25654,
    n43407, n26552, n25712, n25679, n25694, n25693, n42353, n43835, n32345,
    n31210, n25740, n33784, n34836, n42100, n25753, n31223, n25752, n35378,
    n25760, n35376, n25767, n31268, n25766, n37124, n25774, n25772, n25773,
    n37445, n25778, n25777, n36375, n25783, n25781, n25782, n25787, n25786,
    n43695, n25790, n25792, n25791, n36792, n36001, n25794, n31214, n25793,
    n25795, n25799, n25802, n25801, n25806, n25804, n25803, n25805, n25814,
    n25808, n25807, n25812, n25810, n25809, n25811, n25813, n25830, n25816,
    n25815, n25820, n25818, n25817, n25819, n25828, n25822, n25821, n25826,
    n25824, n25823, n25825, n25827, n25829, n25831, n25835, n25832, n25848,
    n25846, n25845, n25847, n25852, n25851, n25856, n25854, n25853, n25855,
    n25864, n25858, n25857, n25862, n25860, n25859, n25861, n25863, n25880,
    n25866, n25865, n25870, n25868, n25867, n25869, n25878, n25872, n25871,
    n25876, n25874, n25873, n25875, n25877, n25879, n25881, n25888, n44034,
    n25884, n25882, n25883, n25887, n25886, n26084, n40709, n25890, n25891,
    n25899, n25898, n25903, n25901, n25900, n25902, n25911, n25905, n25904,
    n25909, n25907, n25906, n25908, n25910, n25913, n25912, n25917, n25915,
    n25914, n25916, n25925, n25919, n25918, n25923, n25921, n25920, n25922,
    n25924, n25929, n26569, n25949, n25945, n25947, n25946, n38642, n25957,
    n38641, n39555, n36889, n36894, n38652, n38645, n38648, n25958, n25953,
    n28539, n25981, n40091, n25954, n25955, n25991, n25956, n28545, n25961,
    n28541, n25959, n25960, n25989, n25964, n25966, n25969, n25967, n38799,
    n25974, n38384, n40093, n25980, n26565, n25982, n40786, n25994, n25997,
    n25996, n26001, n25999, n25998, n26000, n26009, n26003, n26002, n26007,
    n26005, n26004, n26006, n26008, n26025, n26011, n26010, n26015, n26013,
    n26012, n26014, n26023, n26017, n26016, n26021, n26019, n26018, n26020,
    n26022, n26024, n26026, n43286, n26027, n26037, n37237, n35875, n35877,
    n35501, n35502, n26041, n34829, n37235, n26042, n37227, n38256, n26043,
    n26696, n31717, n26045, n42405, n26049, n26055, n26050, n26586, n44107,
    n26052, n26053, n38253, n26054, n26083, n34514, n43803, n28885, n26077,
    n26070, n26066, n26067, n26068, n26072, n26071, n26075, n41129, n26073,
    n26074, n26076, n26088, n26087, n26089, n26098, n26097, n26104, n26102,
    n26101, n26103, n26108, n26106, n26105, n26107, n26128, n26110, n26109,
    n26114, n26112, n26111, n26113, n26122, n26116, n26115, n26120, n26118,
    n26117, n26119, n26121, n26126, n26124, n26123, n26125, n26127, n26129,
    n31983, n26132, n26130, n26131, n26133, n26140, n26147, n26149, n26156,
    n26155, n26161, n26158, n26160, n26166, n26162, n26164, n26163, n26165,
    n26169, n26170, n26176, n26175, n35801, n27870, n26187, n26186, n26188,
    n26190, n26194, n31764, n26215, n26208, n43159, n42699, n26220, n26217,
    n34863, n34859, n36601, n26219, n26213, n35796, n36600, n26218, n26212,
    n26216, n26561, n28067, n26222, n28065, n26221, n40767, n26272, n26229,
    n37654, n26230, n26234, n26231, n26258, n26364, n26247, n26236, n26270,
    n26237, n37039, n26238, n38628, n26266, n26253, n26243, n26241, n36569,
    n26242, n26244, n26246, n26252, n26248, n37612, n26249, n26281, n26265,
    n26375, n26256, n26365, n26255, n26264, n26374, n26262, n26259, n26354,
    n26261, n26263, n26279, n26371, n26269, n26273, n26370, n26267, n26268,
    n26277, n26361, n26275, n26353, n26274, n26276, n26278, n26280, n26284,
    n26287, n26335, n26290, n26289, n26296, n26291, n26294, n26293, n26295,
    n26308, n26297, n26300, n26299, n26306, n26304, n26303, n26305, n26307,
    n26326, n26309, n26314, n26311, n26313, n26316, n26315, n26324, n26320,
    n26318, n26319, n26322, n26321, n26325, n26329, n26333, n36485, n26336,
    n26334, n26342, n26337, n26387, n26344, n26343, n39523, n26357, n26359,
    n26366, n26381, n26372, n26377, n26376, n26378, n26380, n26382, n26386,
    n38376, n26388, n27855, n26420, n26430, n26433, n26452, n26435, n26438,
    n26441, n26442, n26443, n26448, n26451, n26453, n26485, n26454, n26455,
    n38373, n36488, n26473, n26461, n32943, n26465, n26463, n26464, n33569,
    n28119, n26470, n26469, n26467, n26468, n37290, n34880, n26472, n37310,
    n26471, n32942, n26475, n26474, n26480, n36853, n26481, n26482, n38374,
    n26491, n26502, n26504, n31772, n43755, n26556, n26510, n26511, n43886,
    n26517, n26524, n26523, n26532, n26531, n26539, n26538, n40154, n26544,
    n40159, n26554, n26547, n26548, n26549, n43877, n39737, n26553, n26555,
    n26562, n26577, n26563, n26567, n40704, n40695, n26583, n27822, n26584,
    n26597, n29569, n26595, n40803, n31468, n26588, n26589, n26593, n26590,
    n31469, n31679, n26591, n26592, n26594, n26599, n26602, n26601, n26606,
    n26604, n26603, n26605, n26614, n26608, n26607, n26612, n26610, n26609,
    n26611, n26613, n26630, n26616, n26615, n26620, n26618, n26617, n26619,
    n26628, n26622, n26621, n26626, n26624, n26623, n26625, n26627, n26629,
    n26631, n26632, n26635, n26639, n26638, n26643, n26641, n26640, n26642,
    n26670, n26645, n26644, n26649, n26647, n26646, n26648, n26657, n26651,
    n26650, n26655, n26653, n26652, n26654, n26656, n26668, n26661, n26660,
    n26666, n26664, n26663, n26665, n26667, n26669, n26671, n31973, n26674,
    n26672, n26673, n26675, n26682, n26690, n26692, n41125, n41020, n26697,
    n43566, n29613, n26698, n26699, n26710, n26701, n26700, n26709, n26716,
    n26721, n26720, n26942, n26723, n26722, n26725, n26724, n26730, n26728,
    n26727, n26729, n26734, n26732, n26731, n26733, n26753, n26736, n26735,
    n26743, n26739, n26738, n26741, n26740, n26742, n26751, n26745, n26744,
    n26749, n26747, n26746, n26748, n26750, n26752, n26755, n26754, n26759,
    n26757, n26756, n26758, n26767, n26761, n26760, n26765, n26763, n26762,
    n26764, n26766, n26786, n26770, n26769, n26774, n26772, n26771, n26773,
    n26778, n26776, n26775, n26777, n26784, n26782, n26781, n26783, n26785,
    n39670, n26788, n26787, n26797, n26793, n26792, n26795, n26794, n26796,
    n26805, n26799, n26798, n26803, n26801, n26800, n26802, n26804, n26826,
    n26810, n26809, n26812, n26811, n26816, n26814, n26813, n26815, n26824,
    n26822, n26821, n26823, n26825, n26830, n26829, n26836, n26834, n26833,
    n26835, n26847, n26840, n26839, n26845, n26843, n26842, n26844, n26846,
    n26870, n26851, n26850, n26857, n26855, n26854, n26856, n26868, n26861,
    n26860, n26866, n26864, n26863, n26865, n26867, n26869, n43500, n26872,
    n26871, n26876, n26874, n43483, n26873, n26875, n26885, n43495, n26880,
    n26879, n43490, n43509, n26883, n26881, n26882, n26884, n26889, n26887,
    n26886, n26888, n26907, n26890, n26893, n26892, n26897, n26895, n26894,
    n26896, n26905, n26899, n26898, n26903, n26901, n26900, n26902, n26904,
    n26906, n41569, n41568, n42697, n26918, n26915, n26917, n26920, n37269,
    n29511, n26922, n26921, n39701, n26928, n26926, n26925, n26927, n26932,
    n26930, n26929, n26931, n26934, n26933, n36590, n32348, n26936, n31228,
    n26935, n26937, n26941, n26943, n26946, n26945, n26950, n26948, n26947,
    n26949, n26958, n26952, n26951, n26956, n26954, n26953, n26955, n26957,
    n26974, n26960, n26959, n26964, n26962, n26961, n26963, n26972, n26966,
    n26965, n26970, n26968, n26967, n26969, n26971, n26973, n26975, n26976,
    n28484, n26984, n26983, n26988, n26986, n26985, n26987, n27019, n26990,
    n26989, n26994, n26992, n26991, n26993, n27002, n26996, n26995, n27000,
    n26998, n26997, n26999, n27001, n27017, n27008, n27005, n27007, n27015,
    n27013, n27012, n27014, n27016, n27018, n27020, n27025, n31995, n27023,
    n27021, n27022, n27024, n27031, n27039, n27038, n40481, n38144, n39786,
    n27711, n36049, n36040, n27288, n27068, n36047, n27230, n27069, n34042,
    n29442, n36041, n34773, n32515, n27114, n27113, n27121, n27135, n32808,
    n32208, n27252, n27254, n27316, n27284, n27283, n27286, n27285, n27290,
    n27287, n27289, n27298, n27292, n27291, n27296, n27294, n27293, n27295,
    n27297, n27300, n27299, n27305, n27303, n27302, n27304, n27313, n27307,
    n27306, n27311, n27309, n27308, n27310, n27312, n36526, n36666, n36969,
    n27334, n36190, n36230, n39395, n40244, n41541, n28757, n33487, n27403,
    n33501, n32672, n27442, n27441, n27448, n27450, n27455, n27461, n31802,
    n30706, n32475, n29940, n27581, n31801, n41542, n40422, n40141, n27598,
    n36519, n40170, n40166, n40271, n39622, n39624, n40382, n40443, n39386,
    n39451, n40824, n40251, n27641, n41536, n27624, n27793, n27621, n40389,
    n39405, n39398, n40471, n40417, n39780, n40521, n39776, n27622, n41538,
    n27645, n27623, n27633, n40243, n40830, n41539, n32361, n27631, n27635,
    n27634, n27636, n27652, n27651, n27639, n27637, n27638, n27649, n27640,
    n27643, n27642, n27648, n27644, n27646, n27647, n27650, n27657, n27683,
    n27662, n35975, n36665, n36974, n27686, n27688, n36427, n27692, n27691,
    n27693, n27694, n35859, n27698, n27699, n27701, n37107, n37106, n36192,
    n40132, n27703, n36211, n27708, n27714, n27712, n37710, n27716, n36885,
    n37569, n38147, n27723, n27725, n27724, n27726, n27730, n37766, n39422,
    n27735, n27736, n38903, n27739, n38904, n40750, n27740, n41146, n28759,
    n27738, n28099, n41252, n28760, n28098, n40202, n40451, n36227, n27806,
    n27779, n27778, n27780, n31671, n29149, n29561, n27782, n27783, n27794,
    n27807, n27808, n41384, n42025, n41257, n40865, n27819, n41410, n27826,
    n41272, n41185, n28477, n27827, n27832, n27830, n41744, n27828, n27829,
    n27831, n29646, n27835, n27840, n27837, n27839, n27838, n41893, n27849,
    n27842, n27850, n40759, n27864, n31714, n27874, n40760, n27877, n42238,
    n42086, n27881, n27884, n27883, n27886, n28198, n27890, n43913, n27933,
    n28158, n27892, n29199, n27896, n27895, n27903, n27902, n27906, n27909,
    n27908, n27913, n27917, n27916, n40299, n34920, n27926, n32180, n27922,
    n43917, n27924, n28077, n27925, n27931, n28159, n33577, n27928, n43896,
    n40285, n27930, n27932, n27937, n27936, n27939, n27938, n27943, n27941,
    n27940, n27942, n27951, n27945, n27944, n27949, n27947, n27946, n27948,
    n27950, n27967, n27953, n27952, n27957, n27955, n27954, n27956, n27965,
    n27959, n27958, n27963, n27961, n27960, n27962, n27964, n27966, n27968,
    n27969, n27970, n27976, n27975, n27980, n27978, n27977, n27979, n27988,
    n27982, n27981, n27986, n27984, n27983, n27985, n27987, n28004, n27990,
    n27989, n27994, n27992, n27991, n27993, n28002, n27996, n27995, n28000,
    n27998, n27997, n27999, n28001, n28003, n28378, n28006, n28005, n28010,
    n28008, n28007, n28009, n28018, n28012, n28011, n28016, n28014, n28013,
    n28015, n28017, n28034, n28020, n28019, n28024, n28022, n28021, n28023,
    n28032, n28026, n28025, n28030, n28028, n28027, n28029, n28031, n28033,
    n28377, n28035, n28042, n32001, n28040, n28038, n28551, n28055, n28058,
    n28057, n28063, n28064, n28073, n28066, n42105, n28069, n42109, n28068,
    n28070, n41698, n42557, n28071, n28072, n28087, n28083, n28078, n28081,
    n28080, n28082, n28086, n28089, n28094, n28104, n41527, n43774, n43326,
    n43217, n43000, n42473, n42438, n42393, n40626, n42847, n42457, n40648,
    n40294, n41176, n40157, n40574, n40320, n28121, n28120, n36501, n40319,
    n38828, n38829, n40573, n40362, n40363, n39722, n39721, n40948, n38941,
    n39471, n41504, n40293, n40296, n42061, n40647, n40646, n42145, n40671,
    n40670, n42429, n40625, n40624, n42260, n39222, n37716, n42345, n37717,
    n37452, n42856, n39693, n40107, n42960, n39749, n39913, n43546, n40918,
    n41203, n43654, n41719, n41913, n43897, n28161, n28154, n28155, n28157,
    n28160, n41919, n28374, n28164, n39758, n28168, n28166, n28165, n28167,
    n39910, n28172, n28170, n28169, n28171, n40923, n28177, n28176, n28174,
    n28173, n28175, n41209, n29525, n28181, n28179, n28178, n28180, n41725,
    n28185, n28183, n28182, n28184, n41724, n41928, n28190, n28188, n28187,
    n28189, n41471, n29484, n28195, n28193, n28192, n28194, n43878, n37288,
    n40602, n40651, n40675, n40629, n39211, n36384, n37736, n28204, n37273,
    n37469, n28205, n39709, n40121, n40120, n39763, n39928, n28207, n40926,
    n40925, n41874, n41213, n41727, n41726, n28208, n28209, n28369, n28214,
    n39482, n28212, n28215, n28221, n28217, n36390, n28219, n28218, n28220,
    n28224, n28231, n28230, n28238, n28237, n28244, n28243, n28251, n28250,
    n28256, n28263, n28270, n36380, n28276, n28283, n28290, n28297, n28296,
    n28306, n28304, n28303, n29520, n28313, n28311, n28310, n28312, n28320,
    n28318, n28317, n28319, n28328, n28326, n28325, n28327, n40936, n28335,
    n28333, n28332, n28334, n28337, n28342, n28340, n28339, n28341, n28344,
    n28343, n41733, n28350, n28348, n28347, n28349, n28352, n28351, n41941,
    n28358, n28356, n28355, n28357, n28360, n28359, n39571, n28365, n28363,
    n28362, n28364, n28367, n28366, n28376, n28375, n28412, n28417, n28380,
    n28379, n28384, n28382, n28381, n28383, n28392, n28386, n28385, n28390,
    n28388, n28387, n28389, n28391, n28408, n28394, n28393, n28398, n28396,
    n28395, n28397, n28406, n28400, n28399, n28404, n28402, n28401, n28403,
    n28405, n28407, n28416, n28409, n28410, n28411, n28524, n28450, n28449,
    n28419, n28418, n28423, n28421, n28420, n28422, n28431, n28425, n28424,
    n28429, n28427, n28426, n28428, n28430, n28447, n28433, n28432, n28437,
    n28435, n28434, n28436, n28445, n28439, n28438, n28443, n28441, n28440,
    n28442, n28444, n28446, n28603, n28448, n28452, n28602, n28451, n28458,
    n28453, n28456, n28454, n28455, n28457, n28462, n43031, n28467, n28662,
    n28470, n28472, n42501, n28480, n42587, n28486, n28488, n28487, n28489,
    n41989, n42580, n28493, n28506, n28496, n42579, n28560, n41999, n28495,
    n28852, n42372, n28498, n28500, n28499, n28501, n28552, n28513, n28515,
    n28514, n28516, n28521, n28520, n29684, n42186, n41896, n28526, n42403,
    n42161, n28527, n28528, n28532, n28530, n28529, n28531, n28540, n40796,
    n28544, n28558, n28542, n41962, n41963, n43335, n28543, n28546, n42919,
    n28547, n28548, n42364, n42826, n41990, n42675, n42365, n28561, n28562,
    n28565, n28564, n28569, n28567, n28566, n28568, n28601, n28571, n28570,
    n28575, n28573, n28572, n28574, n28583, n28577, n28576, n28581, n28579,
    n28578, n28580, n28582, n28599, n28589, n28588, n28597, n28595, n28594,
    n28596, n28598, n28600, n28605, n28607, n28606, n28611, n28609, n28610,
    n28614, n28658, n28618, n28617, n28622, n28620, n28619, n28621, n28630,
    n28624, n28623, n28628, n28626, n28625, n28627, n28629, n28646, n28632,
    n28631, n28636, n28634, n28633, n28635, n28644, n28638, n28637, n28642,
    n28640, n28639, n28641, n28643, n28645, n28707, n28647, n28653, n28651,
    n28649, n28650, n28652, n28774, n28659, n43377, n28833, n28664, n28670,
    n28667, n28666, n28721, n28677, n28676, n28681, n28679, n28678, n28680,
    n28685, n28683, n28682, n28684, n28705, n28687, n28686, n28691, n28689,
    n28688, n28690, n28699, n28693, n28692, n28697, n28695, n28694, n28696,
    n28698, n28703, n28701, n28700, n28702, n28704, n28807, n28806, n28708,
    n28710, n28709, n28713, n28711, n28712, n28716, n28718, n28717, n42979,
    n42367, n28730, n28733, n42828, n43028, n28736, n28739, n28738, n28740,
    n28750, n41117, n41119, n28770, n41104, n28777, n28776, n28781, n28779,
    n28778, n28780, n28789, n28783, n28782, n28787, n28785, n28784, n28786,
    n28788, n28805, n28791, n28790, n28795, n28793, n28792, n28794, n28803,
    n28797, n28796, n28801, n28799, n28798, n28800, n28802, n28804, n43240,
    n28808, n28815, n28809, n28813, n28811, n28812, n28814, n28818, n43720,
    n28821, n43120, n28824, n28823, n28831, n29632, n28830, n28843, n28837,
    n28836, n28846, n28876, n41988, n28847, n28849, n28850, n28859, n28862,
    n28861, n28863, n29674, n28874, n28868, n28867, n28871, n28881, n28875,
    n28878, n28884, n42488, n43564, n28883, n28892, n28888, n28887, n28890,
    n28889, n28893, n28897, n28898, n28899, n28902, n28900, n28901, n29541,
    n28906, n29750, n29538, n28904, n28903, n28905, n28950, n29092, n29095,
    n28907, n28908, n28937, n28909, n29150, n28910, n28911, n29557, n28930,
    n28912, n29556, n29148, n28913, n28914, n28920, n29560, n28918, n28915,
    n29761, n29151, n29558, n28916, n28917, n28919, n28921, n28926, n29084,
    n29089, n28923, n28922, n28924, n28925, n28927, n28932, n29057, n29178,
    n28929, n28936, n28931, n28933, n28935, n28938, n28939, n28942, n28940,
    n28941, n29164, n28945, n28944, n41672, n28948, n28946, n32843, n28947,
    n41380, n42012, n28949, n29175, n28952, n28951, n28954, n28953, n28956,
    n28955, n28958, n28957, n28959, n28960, n28962, n29093, n29174, n28961,
    n28964, n28963, n28966, n28965, n28968, n28967, n28972, n28970, n28969,
    n28971, n28980, n28974, n28973, n28978, n28976, n28975, n28977, n28979,
    n28996, n28982, n28981, n28986, n28984, n28983, n28985, n28994, n28988,
    n28987, n28992, n28990, n28989, n28991, n28993, n28995, n29075, n29077,
    n29004, n29001, n31686, n28998, n29043, n28997, n28999, n35494, n29000,
    n29002, n29003, n29006, n29005, n29010, n29008, n29007, n29009, n29018,
    n29012, n29011, n29016, n29014, n29013, n29015, n29017, n29034, n29020,
    n29019, n29024, n29022, n29021, n29023, n29032, n29026, n29025, n29030,
    n29028, n29027, n29029, n29031, n29033, n29070, n29072, n29042, n29039,
    n29069, n29036, n29048, n29035, n29037, n35979, n29038, n29040, n29041,
    n29047, n29044, n29061, n29045, n29046, n29052, n29049, n29065, n29050,
    n29051, n29054, n29053, n29056, n29058, n29060, n29059, n29080, n29062,
    n29064, n29063, n29066, n29068, n29067, n29071, n29074, n29073, n29076,
    n29079, n29078, n29083, n29081, n29082, n29088, n29086, n29087, n29090,
    n29091, n29100, n29094, n29097, n29096, n29098, n29099, n29102, n29101,
    n29106, n29104, n29103, n29105, n29114, n29108, n29107, n29112, n29110,
    n29109, n29111, n29113, n29130, n29116, n29115, n29120, n29118, n29117,
    n29119, n29128, n29122, n29121, n29126, n29124, n29123, n29125, n29127,
    n29129, n29233, n29133, n29166, n29131, n29168, n29132, n29135, n29134,
    n29137, n29136, n29139, n29138, n29141, n29140, n29143, n29142, n29145,
    n29144, n29147, n29146, n29159, n29156, n29154, n29152, n29153, n29155,
    n29157, n29158, n29161, n29160, n29163, n29162, n29165, n29235, n29167,
    n29231, n29170, n29169, n29173, n29549, n29172, n29177, n29226, n29176,
    n29180, n29179, n29182, n29181, n29184, n29183, n29186, n29185, n29188,
    n29187, n29190, n29189, n29192, n29191, n29194, n29193, n29196, n29195,
    n29198, n29197, n29201, n29200, n29203, n29202, n29206, n29205, n29208,
    n29207, n29210, n29209, n29212, n29211, n29214, n29213, n29216, n29215,
    n29218, n29217, n29220, n29219, n29223, n29222, n29225, n29224, n29228,
    n29227, n29230, n29229, n29232, n29239, n29234, n29237, n29236, n29238,
    n29240, n29243, n29241, n29242, n29245, n31168, n29244, n29247, n29246,
    n29249, n29248, n29251, n29250, n29253, n29252, n29255, n29254, n29257,
    n29256, n29259, n29258, n29261, n29260, n29263, n29262, n29265, n29264,
    n29267, n29266, n29269, n29268, n29271, n29270, n29273, n29272, n29275,
    n29274, n29277, n29276, n29279, n29278, n29281, n29280, n29283, n29282,
    n29285, n29284, n29287, n29286, n29289, n29288, n29291, n29290, n29293,
    n29292, n29295, n29294, n29297, n29296, n29299, n29298, n29301, n29300,
    n29303, n29302, n29307, n29306, n29313, n29434, n29310, n40723, n29309,
    n29312, n29311, n33900, n29315, n29314, n29317, n29316, n37757, n29319,
    n29318, n29321, n29320, n29326, n29323, n29322, n29325, n29324, n33821,
    n29328, n29327, n29330, n29329, n29332, n35904, n29331, n29334, n29333,
    n29336, n29339, n29335, n29338, n29337, n29341, n29340, n29343, n29342,
    n34547, n29345, n32853, n29344, n29347, n29346, n29352, n29349, n29348,
    n29351, n29350, n33662, n29354, n29353, n29356, n29355, n33646, n29358,
    n29357, n29360, n29359, n37088, n29362, n29361, n29364, n29363, n35542,
    n29366, n29365, n29368, n29367, n29370, n29369, n29372, n29371, n32969,
    n29374, n33074, n29373, n29376, n29375, n29378, n29377, n29380, n29379,
    n29386, n29383, n29382, n29385, n29384, n29388, n29387, n29390, n29389,
    n29403, n29392, n36159, n29391, n29394, n29393, n29396, n29412, n29395,
    n29398, n29397, n29400, n35645, n29399, n29402, n29401, n29405, n29404,
    n29407, n29406, n32968, n29409, n29408, n29411, n29410, n29414, n33757,
    n29413, n29416, n29415, n29418, n33515, n29417, n29420, n29419, n29425,
    n29422, n29435, n29421, n29424, n29423, n29427, n29426, n29429, n29428,
    n29431, n29430, n29433, n29432, n29438, n29437, n29441, n29440, n29443,
    n29444, n29690, n29445, n29446, n29448, n32362, n29447, n30030, n43994,
    n29451, n29450, n29453, n29452, n29455, n29454, n29457, n29456, n29459,
    n29458, n29460, n29464, n29463, n29466, n29465, n29468, n29467, n29470,
    n29469, n29473, n29472, n29475, n29474, n29477, n29476, n29479, n29478,
    n29481, n29480, n29483, n29482, n29486, n29485, n29488, n29487, n29490,
    n29489, n29492, n29491, n29495, n29494, n29497, n29496, n29499, n29498,
    n29501, n29500, n29503, n29502, n29505, n29504, n29508, n29507, n29510,
    n29509, n29513, n29512, n29515, n29514, n29517, n29516, n29519, n29518,
    n29522, n29521, n29524, n29523, n29527, n29526, n29529, n29528, n29531,
    n29530, n29533, n29532, n29535, n29534, n29537, n29536, n29539, n29548,
    n29540, n29542, n29753, n29546, n29718, n29543, n29544, n29754, n29545,
    n29547, n29552, n29551, n29555, n29554, n29564, n29559, n29562, n29563,
    n34518, n29565, n29567, n29566, n34512, n44093, n29571, n29570, n29573,
    n29572, n29576, n29575, n29578, n29577, n37228, n29582, n37508, n29581,
    n29584, n29583, n29586, n29627, n29585, n29588, n29587, n29679, n29590,
    n29589, n29592, n29591, n29622, n29594, n29593, n29596, n29595, n29598,
    n29597, n29600, n29599, n43032, n29602, n29601, n29604, n29603, n29656,
    n29606, n29605, n29608, n29607, n38791, n29610, n29651, n29609, n29612,
    n29611, n29615, n29645, n29614, n29617, n29616, n29619, n29618, n29621,
    n29620, n29624, n29623, n29626, n29625, n29629, n29628, n29631, n29630,
    n29634, n29633, n29636, n29635, n29638, n29637, n29640, n29639, n29642,
    n43565, n29641, n29644, n29643, n29648, n29647, n29650, n29649, n29653,
    n29652, n29655, n29654, n29658, n29657, n29660, n29659, n29662, n29661,
    n29664, n29663, n36991, n29666, n29665, n29668, n29667, n29671, n29670,
    n29673, n29672, n29676, n29675, n29678, n29677, n29681, n29680, n29683,
    n29682, n29686, n29685, n29688, n29687, n36057, n35442, n29689, n29695,
    n29691, n42018, n29692, n30873, n29693, n29694, n29713, n29697, n29696,
    n29699, n29698, n36103, n29701, n34830, n29700, n29703, n29702, n29705,
    n29708, n29704, n29707, n29706, n29710, n29709, n29712, n29711, n29715,
    n29714, n29717, n29716, n29720, n29719, n29723, n29722, n29995, n30048,
    n29870, n29724, n29725, n31370, n29843, n29738, n29731, n30560, n29844,
    n30870, n29727, n29729, n30777, n29728, n29730, n29732, n29737, n29734,
    n41344, n30559, n29733, n29740, n29735, n29736, n43989, n29996, n29739,
    n29742, n29741, n29748, n29744, n29743, n29745, n29746, n29747, n29758,
    n29751, n29757, n29755, n29756, n29765, n29759, n29760, n29762, n29763,
    n29764, n29772, n29769, n29766, n29767, n29768, n29770, n29771, n29774,
    n29773, n29776, n29775, n29778, n29777, n29780, n29779, n29782, n29781,
    n29784, n29783, n29786, n29785, n29788, n29787, n29790, n29789, n29792,
    n29791, n29794, n29793, n29796, n29795, n29798, n29797, n29800, n29799,
    n29802, n29801, n29804, n29803, n29806, n29805, n29808, n29807, n29810,
    n29809, n29812, n29811, n29814, n29813, n29816, n29815, n29818, n29817,
    n29820, n29819, n29822, n29821, n29824, n29823, n29826, n29825, n29828,
    n29827, n29830, n29829, n29832, n29831, n29834, n29833, n29837, n29836,
    n31014, n29838, n29923, n29881, n43993, n29884, n29845, n41382, n30809,
    n29840, n30900, n31045, n41095, n31015, n29839, n29854, n30862, n30812,
    n31018, n29852, n32374, n30705, n31019, n41350, n30894, n30813, n29850,
    n29842, n29848, n30027, n30011, n29846, n29857, n29847, n30814, n29849,
    n29851, n29853, n29927, n30797, n29856, n30800, n29855, n29867, n31040,
    n29865, n30801, n29863, n30049, n29858, n29859, n29861, n30773, n29860,
    n30802, n29862, n29864, n29866, n29897, n30774, n29869, n29868, n29880,
    n29878, n30750, n30778, n29876, n29871, n29872, n29874, n29873, n30779,
    n29875, n29877, n29879, n30597, n30877, n30993, n29883, n30994, n30836,
    n30789, n30857, n30000, n30786, n29882, n29894, n30707, n30832, n29892,
    n29890, n29912, n29885, n29886, n29887, n29888, n30790, n29889, n29891,
    n29893, n29896, n29898, n30761, n29895, n29908, n30764, n29906, n30990,
    n30765, n29904, n29924, n29899, n29911, n29902, n29900, n29901, n30766,
    n29903, n29905, n29907, n29910, n30702, n29909, n29922, n29920, n29918,
    n29915, n29913, n29914, n29916, n30708, n29917, n29919, n29921, n31047,
    n30740, n29926, n30737, n29925, n29937, n29935, n30741, n29933, n29928,
    n29929, n29930, n29931, n30742, n29932, n29934, n29936, n31003, n29939,
    n31006, n29938, n29946, n31002, n29944, n31007, n29942, n29941, n29943,
    n29945, n29948, n29947, n29954, n29952, n29950, n29949, n29951, n29953,
    n29956, n29955, n29962, n29960, n29958, n29957, n29959, n29961, n29964,
    n29963, n29970, n29968, n29966, n29965, n29967, n29969, n29974, n29972,
    n29971, n29973, n29978, n29976, n29975, n29977, n29982, n29980, n29979,
    n29981, n29986, n29984, n29983, n29985, n29990, n29988, n29987, n29989,
    n29994, n29992, n29991, n29993, n30213, n30861, n30029, n30848, n30014,
    n30821, n29999, n29998, n30010, n30008, n30824, n30006, n30001, n30002,
    n30003, n30004, n30825, n30005, n30007, n30009, n30845, n30013, n30012,
    n30024, n30022, n30849, n30020, n30015, n30016, n30017, n30018, n30850,
    n30019, n30021, n30023, n30026, n30858, n30025, n30039, n30037, n30035,
    n30028, n30031, n30033, n30032, n30863, n30034, n30036, n30038, n30041,
    n30040, n30047, n30045, n30043, n30042, n30044, n30046, n30726, n30056,
    n30050, n30558, n30052, n30051, n30730, n30054, n30729, n30053, n30055,
    n30060, n30058, n30057, n30059, n30064, n30062, n30061, n30063, n30068,
    n30066, n30065, n30067, n30070, n30069, n30076, n30074, n30072, n30071,
    n30073, n30075, n30080, n30078, n30077, n30079, n30084, n30082, n30081,
    n30083, n31026, n30086, n31030, n30085, n30092, n31027, n30090, n31031,
    n30088, n30087, n30089, n30091, n30094, n30093, n30100, n30098, n30096,
    n30095, n30097, n30099, n30102, n30101, n30108, n30106, n30104, n30103,
    n30105, n30107, n30110, n30109, n30116, n30114, n30112, n30111, n30113,
    n30115, n30118, n30117, n30124, n30122, n30120, n30119, n30121, n30123,
    n30126, n30125, n30132, n30130, n30128, n30127, n30129, n30131, n30917,
    n30134, n30921, n30133, n30140, n30918, n30138, n30922, n30136, n30135,
    n30137, n30139, n30142, n30141, n30148, n30146, n30144, n30143, n30145,
    n30147, n30150, n30149, n30156, n30154, n30152, n30151, n30153, n30155,
    n30158, n30157, n30164, n30162, n30160, n30159, n30161, n30163, n30168,
    n30166, n30165, n30167, n30172, n30170, n30169, n30171, n30176, n30174,
    n30173, n30175, n30180, n30178, n30177, n30179, n30184, n30182, n30181,
    n30183, n30188, n30186, n30185, n30187, n30192, n30190, n30189, n30191,
    n30196, n30194, n30193, n30195, n30200, n30198, n30197, n30199, n30204,
    n30202, n30201, n30203, n30206, n30205, n30212, n30210, n30208, n30207,
    n30209, n30211, n30833, n30219, n30215, n30214, n30838, n30217, n30216,
    n30218, n30223, n30221, n30220, n30222, n30929, n30225, n30930, n30224,
    n30231, n30933, n30229, n30934, n30227, n30226, n30228, n30230, n30233,
    n30232, n30239, n30237, n30235, n30234, n30236, n30238, n30241, n30240,
    n30247, n30245, n30243, n30242, n30244, n30246, n30249, n30248, n30255,
    n30253, n30251, n30250, n30252, n30254, n30257, n30256, n30263, n30261,
    n30259, n30258, n30260, n30262, n30267, n30265, n30264, n30266, n30271,
    n30269, n30268, n30270, n30273, n30272, n30279, n30277, n30275, n30274,
    n30276, n30278, n31039, n30281, n31041, n30280, n30287, n31044, n30285,
    n31046, n30283, n30282, n30284, n30286, n30289, n30288, n30295, n30293,
    n30291, n30290, n30292, n30294, n30297, n30296, n30303, n30301, n30299,
    n30298, n30300, n30302, n30305, n30304, n30311, n30309, n30307, n30306,
    n30308, n30310, n30313, n30312, n30319, n30317, n30315, n30314, n30316,
    n30318, n30321, n30320, n30327, n30325, n30323, n30322, n30324, n30326,
    n30329, n30328, n30335, n30333, n30331, n30330, n30332, n30334, n30337,
    n30336, n30343, n30341, n30339, n30338, n30340, n30342, n30347, n30345,
    n30344, n30346, n30351, n30349, n30348, n30350, n30355, n30353, n30352,
    n30354, n30359, n30357, n30356, n30358, n30363, n30361, n30360, n30362,
    n30367, n30365, n30364, n30366, n30369, n30368, n30375, n30373, n30371,
    n30370, n30372, n30374, n30379, n30377, n30376, n30378, n30383, n30381,
    n30380, n30382, n30387, n30385, n30384, n30386, n30391, n30389, n30388,
    n30390, n30395, n30393, n30392, n30394, n30399, n30397, n30396, n30398,
    n30401, n30400, n30407, n30405, n30403, n30402, n30404, n30406, n30409,
    n30408, n30415, n30413, n30411, n30410, n30412, n30414, n30417, n30416,
    n30423, n30421, n30419, n30418, n30420, n30422, n30425, n30424, n30431,
    n30429, n30427, n30426, n30428, n30430, n30435, n30433, n30432, n30434,
    n30439, n30437, n30436, n30438, n30977, n30441, n30978, n30440, n30447,
    n30981, n30445, n30982, n30443, n30442, n30444, n30446, n30449, n30448,
    n30455, n30453, n30451, n30450, n30452, n30454, n30457, n30456, n30463,
    n30461, n30459, n30458, n30460, n30462, n30465, n30464, n30471, n30469,
    n30467, n30466, n30468, n30470, n30473, n30472, n30479, n30477, n30475,
    n30474, n30476, n30478, n30481, n30480, n30487, n30485, n30483, n30482,
    n30484, n30486, n30489, n30488, n30495, n30493, n30491, n30490, n30492,
    n30494, n30497, n30496, n30503, n30501, n30499, n30498, n30500, n30502,
    n30507, n30505, n30504, n30506, n30511, n30509, n30508, n30510, n30513,
    n30512, n30519, n30517, n30515, n30514, n30516, n30518, n30521, n30520,
    n30527, n30525, n30523, n30522, n30524, n30526, n30529, n30528, n30535,
    n30533, n30531, n30530, n30532, n30534, n30537, n30536, n30543, n30541,
    n30539, n30538, n30540, n30542, n30545, n30544, n30551, n30549, n30547,
    n30546, n30548, n30550, n30557, n30715, n30553, n30552, n30555, n30718,
    n30554, n30556, n30562, n30599, n30719, n30561, n30566, n30564, n30563,
    n30565, n30570, n30568, n30567, n30569, n30574, n30572, n30571, n30573,
    n30578, n30576, n30575, n30577, n30584, n30580, n30579, n30582, n30581,
    n30583, n30586, n30585, n30588, n30587, n30594, n30592, n30590, n30589,
    n30591, n30593, n30749, n30596, n30595, n30605, n30603, n30753, n30601,
    n30598, n30754, n30600, n30602, n30604, n30607, n30606, n30613, n30611,
    n30609, n30608, n30610, n30612, n30615, n30614, n30621, n30619, n30617,
    n30616, n30618, n30620, n30623, n30622, n30629, n30627, n30625, n30624,
    n30626, n30628, n30631, n30630, n30637, n30635, n30633, n30632, n30634,
    n30636, n30639, n30638, n30645, n30643, n30641, n30640, n30642, n30644,
    n30647, n30646, n30653, n30651, n30649, n30648, n30650, n30652, n30655,
    n30654, n30661, n30659, n30657, n30656, n30658, n30660, n30663, n30662,
    n30669, n30667, n30665, n30664, n30666, n30668, n30671, n30670, n30677,
    n30675, n30673, n30672, n30674, n30676, n30679, n30678, n30685, n30683,
    n30681, n30680, n30682, n30684, n30687, n30686, n30693, n30691, n30689,
    n30688, n30690, n30692, n30695, n30694, n30701, n30699, n30697, n30696,
    n30698, n30700, n30965, n30704, n30966, n30703, n30714, n30969, n30712,
    n30970, n30710, n30709, n30711, n30713, n30717, n30716, n30725, n30723,
    n30721, n30720, n30722, n30724, n30728, n30727, n30736, n30734, n30732,
    n30731, n30733, n30735, n30739, n30738, n30748, n30746, n30744, n30743,
    n30745, n30747, n30752, n30751, n30760, n30758, n30756, n30755, n30757,
    n30759, n30763, n30762, n30772, n30770, n30768, n30767, n30769, n30771,
    n30776, n30775, n30785, n30783, n30781, n30780, n30782, n30784, n30788,
    n30787, n30796, n30794, n30792, n30791, n30793, n30795, n30799, n30798,
    n30808, n30806, n30804, n30803, n30805, n30807, n30811, n30810, n30820,
    n30818, n30816, n30815, n30817, n30819, n30823, n30822, n30831, n30829,
    n30827, n30826, n30828, n30830, n30835, n30834, n30844, n30842, n30840,
    n30839, n30841, n30843, n30847, n30846, n30856, n30854, n30852, n30851,
    n30853, n30855, n30860, n30859, n30869, n30867, n30865, n30864, n30866,
    n30868, n30875, n30989, n30872, n30871, n30885, n30883, n30881, n30899,
    n30876, n30879, n30878, n30995, n30880, n30882, n30884, n30887, n30886,
    n30893, n30891, n30889, n30888, n30890, n30892, n30897, n31038, n30896,
    n30895, n30908, n30906, n30904, n30898, n30902, n30901, n31048, n30903,
    n30905, n30907, n30910, n30909, n30916, n30914, n30912, n30911, n30913,
    n30915, n30920, n30919, n30928, n30926, n30924, n30923, n30925, n30927,
    n30932, n30931, n30940, n30938, n30936, n30935, n30937, n30939, n30942,
    n30941, n30948, n30946, n30944, n30943, n30945, n30947, n30950, n30949,
    n30956, n30954, n30952, n30951, n30953, n30955, n30958, n30957, n30964,
    n30962, n30960, n30959, n30961, n30963, n30968, n30967, n30976, n30974,
    n30972, n30971, n30973, n30975, n30980, n30979, n30988, n30986, n30984,
    n30983, n30985, n30987, n30992, n30991, n31001, n30999, n30997, n30996,
    n30998, n31000, n31005, n31004, n31013, n31011, n31009, n31008, n31010,
    n31012, n31017, n31016, n31025, n31023, n31021, n31020, n31022, n31024,
    n31029, n31028, n31037, n31035, n31033, n31032, n31034, n31036, n31043,
    n31042, n31054, n31052, n31050, n31049, n31051, n31053, n44002, n31200,
    n31062, n31059, n31060, n31061, n31190, n31065, n31064, n31067, n31066,
    n31069, n31068, n31071, n31070, n31073, n31072, n31075, n31074, n31077,
    n31076, n31079, n31078, n31081, n31080, n31083, n31082, n31085, n31084,
    n31087, n31086, n31089, n31088, n31091, n31090, n31093, n31092, n31095,
    n31094, n31097, n31096, n31099, n31098, n31101, n31100, n31103, n31102,
    n31105, n31104, n31107, n31106, n31109, n31108, n31111, n31110, n31113,
    n31112, n31115, n31114, n31117, n31116, n31119, n31118, n31121, n31120,
    n31123, n31122, n31125, n31124, n31127, n31126, n31129, n31128, n31131,
    n31130, n31133, n31132, n31135, n31134, n31137, n31136, n31139, n31138,
    n31141, n31140, n31143, n31142, n31145, n31144, n31147, n31146, n31149,
    n31148, n31151, n31150, n31153, n31152, n31155, n31154, n31157, n31156,
    n31159, n31158, n31161, n31160, n31163, n31162, n31165, n31164, n31167,
    n31166, n31170, n31169, n31172, n31171, n31174, n31173, n31176, n31175,
    n31178, n31177, n31180, n31179, n31182, n31181, n31184, n31183, n31186,
    n31185, n31188, n31187, n31192, n31191, n31195, n31194, n31197, n31201,
    n31199, n31198, n43634, n31224, n31204, n31203, n31207, n31206, n31205,
    n43111, n31253, n31209, n31208, n31211, n31229, n31213, n31212, n31215,
    n31248, n31217, n31216, n41758, n31220, n31219, n31218, n41757, n31233,
    n31222, n31221, n31225, n31227, n31226, n31230, n31232, n31231, n32260,
    n31234, n31236, n31235, n31237, n31240, n31239, n31238, n40056, n32225,
    n31262, n31242, n31241, n31245, n31244, n31243, n43696, n31258, n31247,
    n31246, n31249, n31251, n31250, n31254, n31256, n31255, n31257, n31259,
    n31261, n31260, n31263, n31265, n31264, n31267, n31266, n35317, n31270,
    n31269, n31272, n31271, n31275, n31274, n31278, n31277, n31378, n31279,
    n31281, n31280, n31283, n31282, n31287, n31285, n31284, n39675, n31326,
    n31289, n31288, n31292, n31291, n31290, n42803, n31351, n31294, n31293,
    n31297, n31296, n31295, n37112, n31342, n31299, n31298, n31302, n31301,
    n31300, n41659, n31356, n31304, n31303, n31307, n31306, n31305, n38018,
    n31330, n31309, n31308, n31312, n31311, n31310, n41831, n31334, n31314,
    n31313, n31317, n31316, n31315, n38972, n31338, n31319, n31318, n31323,
    n31321, n31320, n37434, n31347, n31325, n31324, n31327, n31329, n31328,
    n31331, n31333, n31332, n31335, n31337, n31336, n31339, n31341, n31340,
    n31343, n31346, n31345, n31348, n31350, n31349, n31352, n31355, n31354,
    n31357, n34517, n44028, n31363, n31362, n31365, n31364, n31367, n31366,
    n31369, n31368, n31373, n31826, n31532, n32844, n31372, n31375, n31481,
    n31376, n31377, n34496, n31446, n31379, n31381, n31380, n31384, n31383,
    n31386, n31385, n31388, n31387, n31390, n31389, n31392, n31391, n31394,
    n31393, n31396, n31395, n31398, n31397, n31400, n31399, n31402, n31401,
    n31404, n31403, n31406, n31405, n31408, n31407, n31410, n31409, n31412,
    n31411, n31414, n31413, n31416, n31415, n31418, n31417, n31420, n31419,
    n31422, n31421, n31424, n31423, n31426, n31425, n31428, n31427, n31430,
    n31429, n31432, n31431, n31434, n31433, n31436, n31435, n31438, n31437,
    n31441, n31440, n32081, n31445, n31443, n31444, n31461, n31459, n31457,
    n34509, n31455, n31450, n31452, n31453, n31454, n31456, n31458, n34499,
    n31460, n31465, n31463, n31462, n31464, n31467, n31466, n31471, n31470,
    n31472, n31474, n31486, n31473, n31475, n31484, n31476, n31479, n31480,
    n31482, n31483, n31485, n35709, n31490, n35708, n31489, n31491, n31504,
    n31503, n31492, n31497, n31494, n31496, n31501, n31499, n31500, n31502,
    n31506, n31505, n31510, n31508, n31509, n31519, n31518, n31513, n31512,
    n31514, n31515, n31516, n31517, n31521, n31520, n31531, n31523, n31528,
    n31526, n31527, n31711, n31529, n31530, n35697, n31537, n31535, n31533,
    n31621, n31536, n31539, n31538, n32207, n31605, n32204, n31540, n31542,
    n31541, n31543, n31661, n31544, n31545, n31547, n31546, n31548, n31643,
    n31549, n31550, n31552, n31551, n31553, n31592, n31554, n31555, n31557,
    n31556, n31558, n31635, n32280, n31559, n31561, n31560, n34351, n31601,
    n34356, n31562, n31564, n31563, n33222, n31614, n31565, n31566, n31568,
    n31567, n32283, n31651, n32279, n31569, n31571, n31570, n32323, n31584,
    n43952, n31572, n31574, n31573, n31575, n31626, n36280, n31576, n31578,
    n31577, n32834, n31630, n32839, n31579, n31581, n31580, n31582, n31583,
    n31586, n31585, n31597, n31587, n31588, n31590, n31589, n43937, n31591,
    n31594, n31593, n31595, n31596, n31599, n31598, n43942, n31600, n31603,
    n31602, n43972, n31604, n31607, n31606, n31608, n31647, n31609, n31611,
    n31610, n31612, n31613, n31616, n31615, n31617, n31656, n32815, n31618,
    n31620, n31619, n32353, n31639, n32328, n31622, n31624, n31623, n34969,
    n31625, n31628, n31627, n43947, n31629, n31632, n31631, n31634, n31637,
    n31636, n43957, n31638, n31641, n31640, n43962, n31642, n31645, n31644,
    n31646, n31649, n31648, n43983, n31650, n31653, n31652, n31654, n31655,
    n31658, n31657, n43977, n31660, n31664, n31663, n31668, n41359, n31791,
    n31678, n31676, n31669, n31675, n31672, n31673, n31674, n31677, n31680,
    n31693, n31683, n31685, n35468, n31691, n31695, n31689, n31702, n31688,
    n31690, n31692, n34285, n31701, n31694, n31699, n31696, n35470, n31698,
    n31700, n31704, n31703, n31707, n31706, n31709, n31708, n31710, n31712,
    n35738, n31784, n31713, n31720, n31719, n31725, n31724, n31723, n42736,
    n31727, n31726, n31730, n31729, n31728, n43305, n31981, n31732, n31731,
    n31735, n31734, n31733, n43121, n31737, n31736, n31740, n31739, n31738,
    n42043, n32055, n31742, n31741, n31745, n31744, n31743, n42942, n32059,
    n31747, n31746, n31749, n31751, n31750, n31754, n31753, n31752, n42688,
    n32047, n31756, n31755, n31758, n31760, n31759, n31763, n31762, n31761,
    n42029, n32051, n31786, n31783, n31767, n31769, n31776, n31774, n31773,
    n31775, n31781, n31778, n31780, n31782, n35742, n31785, n31789, n33488,
    n31792, n35485, n31798, n35484, n31797, n31800, n31799, n32526, n42052,
    n31811, n35917, n33507, n31813, n31812, n31815, n31814, n31822, n32156,
    n31828, n31827, n31830, n31829, n31832, n31831, n31834, n31833, n31836,
    n31835, n31838, n31837, n31840, n31839, n31842, n31841, n31844, n31843,
    n31846, n31845, n31848, n31847, n31850, n31849, n31852, n31851, n31854,
    n31853, n31856, n31855, n31858, n31857, n31860, n31859, n31862, n31861,
    n31864, n31863, n31866, n31865, n31868, n31867, n31870, n31869, n31872,
    n31871, n31874, n31873, n31876, n31875, n31878, n31877, n31880, n31879,
    n31882, n31881, n31884, n31883, n31886, n31885, n31888, n31887, n31890,
    n31889, n39307, n34071, n31893, n31906, n31897, n31902, n31899, n31900,
    n31901, n32234, n31915, n34523, n31914, n32101, n31917, n31918, n31919,
    n31926, n31924, n31940, n31923, n31925, n34478, n31931, n31929, n35631,
    n31928, n31930, n31932, n31934, n31933, n31935, n32076, n31949, n31944,
    n31942, n31939, n31941, n31943, n34477, n31947, n32097, n31945, n31946,
    n31948, n31950, n31952, n31951, n35916, n33163, n33139, n32255, n31955,
    n31957, n31956, n31959, n31958, n31961, n31964, n31963, n31962, n41049,
    n34228, n32015, n31966, n31965, n31967, n31970, n31969, n31968, n41462,
    n34136, n32023, n31972, n31971, n31976, n31975, n31974, n41040, n34166,
    n32011, n31978, n31977, n31980, n31979, n31982, n31986, n31985, n31984,
    n40550, n34189, n32033, n31988, n31987, n31992, n31991, n31990, n39894,
    n32007, n31994, n31993, n31998, n31997, n31996, n41426, n34606, n32019,
    n32000, n31999, n32004, n32003, n32002, n41688, n34074, n32037, n32006,
    n32005, n32008, n32010, n32009, n32012, n32014, n32013, n32016, n32018,
    n32017, n44068, n32020, n32022, n32021, n44073, n32024, n32026, n32025,
    n32027, n32030, n32029, n32028, n41773, n34151, n32041, n32032, n32031,
    n44086, n32034, n32036, n32035, n32038, n32040, n32039, n44063, n32042,
    n32044, n32043, n44044, n32046, n32045, n32048, n44049, n32050, n32049,
    n32052, n44054, n32054, n32053, n32056, n44039, n32058, n32057, n32060,
    n32064, n32063, n32529, n32068, n32534, n32066, n32065, n32067, n32072,
    n32070, n32069, n32071, n32073, n32074, n32077, n32104, n32078, n32096,
    n34580, n32090, n32079, n32088, n32114, n32113, n32086, n32085, n32091,
    n32087, n32089, n32094, n32092, n32093, n33711, n32095, n32100, n32098,
    n32099, n32102, n32103, n32106, n32105, n39931, n32109, n44029, n32108,
    n32112, n32111, n32115, n32135, n35870, n32117, n32125, n32120, n32122,
    n32137, n32124, n32133, n32126, n32129, n32128, n32130, n32132, n32134,
    n32139, n32138, n32140, n32142, n32141, n32146, n32151, n32150, n32153,
    n32152, n32155, n32154, n32158, n43982, n32157, n32160, n32159, n32162,
    n32161, n32164, n32163, n32166, n32165, n39510, n34901, n32170, n37303,
    n32169, n32171, n32900, n32172, n32174, n32173, n32179, n32178, n32182,
    n32181, n32183, n32185, n32184, n32187, n32186, n32189, n32188, n32192,
    n32191, n32195, n32194, n32824, n32816, n32814, n33090, n32203, n32205,
    n34968, n32498, n32497, n32212, n32210, n35459, n32209, n32211, n37280,
    n32216, n32273, n32215, n32222, n32220, n32218, n32219, n32221, n32224,
    n32223, n32227, n32226, n32229, n32228, n32230, n32231, n32241, n32240,
    n34898, n32244, n32242, n32243, n32246, n32245, n32248, n32247, n32250,
    n32249, n32252, n32257, n43932, n32254, n33480, n33481, n32256, n32259,
    n32258, n32262, n32261, n32266, n41081, n32265, n32270, n32268, n32267,
    n32269, n32278, n32272, n33217, n32274, n33216, n32276, n32275, n32277,
    n32813, n33094, n32822, n32282, n32821, n32281, n32288, n32286, n32285,
    n32287, n32289, n32290, n32292, n32291, n32294, n32293, n32298, n32296,
    n32295, n32297, n32306, n32300, n32299, n32304, n32302, n32301, n32303,
    n32305, n32322, n32308, n32307, n32312, n32310, n32309, n32311, n32320,
    n32314, n32313, n32318, n32316, n32315, n32317, n32319, n32321, n32677,
    n32325, n32324, n32333, n32329, n32327, n32326, n32485, n32357, n32331,
    n32332, n32335, n35500, n32338, n32339, n32343, n32342, n32346, n40775,
    n32350, n32349, n32352, n32351, n32355, n32354, n32360, n32356, n32358,
    n32359, n35670, n32365, n32363, n32364, n41363, n32378, n32375, n32377,
    n32376, n32380, n32379, n32382, n32381, n32386, n32384, n32383, n32385,
    n32394, n32388, n32387, n32392, n32390, n32389, n32391, n32393, n32410,
    n32396, n32395, n32400, n32398, n32397, n32399, n32408, n32402, n32401,
    n32406, n32404, n32403, n32405, n32407, n32409, n32613, n32412, n32411,
    n32416, n32414, n32413, n32415, n32424, n32418, n32417, n32422, n32420,
    n32419, n32421, n32423, n32440, n32426, n32425, n32430, n32428, n32427,
    n32429, n32438, n32432, n32431, n32436, n32434, n32433, n32435, n32437,
    n32439, n32612, n32787, n32442, n32441, n32445, n34768, n32443, n32444,
    n32447, n32446, n32451, n32449, n32448, n32450, n32471, n32453, n32452,
    n32457, n32455, n32454, n32456, n32465, n32459, n32458, n32463, n32461,
    n32460, n32462, n32464, n32469, n32467, n32466, n32468, n32470, n32786,
    n40542, n32474, n32473, n32493, n32491, n32476, n32986, n32477, n32478,
    n32487, n35694, n32480, n32479, n34967, n32482, n32481, n32483, n32484,
    n32565, n32486, n32607, n32488, n32490, n32492, n32496, n32495, n32513,
    n32516, n32500, n32503, n32502, n32505, n32504, n32510, n32507, n32508,
    n35740, n32512, n32511, n32514, n32523, n32521, n32517, n32519, n32518,
    n32520, n32522, n32525, n35407, n43930, n32524, n32528, n32527, n32538,
    n32531, n32530, n32536, n32533, n32535, n32537, n32543, n32539, n32541,
    n32542, n32544, n32564, n32548, n32624, n32562, n32626, n44022, n32551,
    n32555, n34286, n32553, n32554, n32560, n32557, n32558, n32559, n32561,
    n32563, n32567, n32985, n33268, n32568, n32569, n32573, n32571, n32570,
    n32572, n32605, n32575, n32574, n32579, n32577, n32576, n32578, n32603,
    n32581, n32580, n32585, n32583, n32582, n32584, n32593, n32587, n32586,
    n32591, n32589, n32588, n32590, n32592, n32601, n32595, n32594, n32599,
    n32597, n32596, n32598, n32600, n32602, n35550, n32604, n32617, n32609,
    n32611, n32610, n32615, n39740, n32614, n32616, n32619, n32618, n32621,
    n32620, n32623, n32622, n32628, n32625, n32627, n32636, n32634, n32632,
    n32633, n32635, n32638, n32637, n32640, n32639, n32642, n32641, n32646,
    n32644, n32643, n32645, n32654, n32648, n32647, n32652, n32650, n32649,
    n32651, n32653, n32670, n32656, n32655, n32660, n32658, n32657, n32659,
    n32668, n32662, n32661, n32666, n32664, n32663, n32665, n32667, n32669,
    n33221, n32676, n32673, n32674, n33066, n32750, n32675, n32683, n32679,
    n32681, n32714, n32682, n32685, n32684, n32689, n32687, n32686, n32688,
    n32697, n32691, n32690, n32695, n32693, n32692, n32694, n32696, n32713,
    n32699, n32698, n32703, n32701, n32700, n32702, n32711, n32705, n32704,
    n32709, n32707, n32706, n32708, n32710, n32712, n32833, n32719, n32715,
    n32717, n32718, n32721, n32720, n32725, n32723, n32722, n32724, n32733,
    n32727, n32726, n32731, n32729, n32728, n32730, n32732, n32749, n32735,
    n32734, n32739, n32737, n32736, n32738, n32747, n32741, n32740, n32745,
    n32743, n32742, n32744, n32746, n32748, n34350, n32755, n32751, n32753,
    n32754, n32791, n32757, n32756, n32761, n32759, n32758, n32760, n32769,
    n32763, n32762, n32767, n32765, n32764, n32766, n32768, n32785, n32771,
    n32770, n32775, n32773, n32772, n32774, n32783, n32777, n32776, n32781,
    n32779, n32778, n32780, n32782, n32784, n33169, n33168, n40809, n32789,
    n32788, n32790, n32797, n32793, n32795, n33206, n32796, n32802, n32801,
    n32804, n32803, n32806, n32805, n32812, n32810, n32809, n32811, n32820,
    n32818, n32817, n32819, n32823, n32832, n32825, n32830, n32828, n32827,
    n32829, n32831, n32836, n32835, n32842, n32837, n32840, n33225, n32841,
    n35918, n33925, n33872, n33873, n33765, n33764, n33766, n33621, n33739,
    n36176, n37324, n40544, n32851, n32866, n32847, n34626, n35642, n32850,
    n32879, n32852, n33870, n33106, n33770, n33516, n32967, n32960, n33116,
    n33705, n33647, n33661, n33856, n34546, n32854, n33970, n32855, n32856,
    n33155, n33819, n33594, n34625, n32872, n32862, n33923, n33891, n32864,
    n39426, n32863, n32877, n41325, n32869, n35945, n32875, n32873, n33892,
    n32874, n32876, n32878, n32888, n37758, n33945, n32975, n35995, n35997,
    n32976, n35842, n32882, n37578, n33835, n33602, n33601, n33814, n32884,
    n41092, n38910, n35939, n41401, n32885, n33894, n39425, n32886, n35942,
    n32887, n40311, n32899, n32897, n32898, n32903, n32901, n32902, n32904,
    n32906, n32905, n32908, n32907, n32912, n32910, n32909, n32911, n32920,
    n32914, n32913, n32918, n32916, n32915, n32917, n32919, n32936, n32922,
    n32921, n32926, n32924, n32923, n32925, n32934, n32928, n32927, n32932,
    n32930, n32929, n32931, n32933, n32935, n34842, n32941, n32937, n32939,
    n33260, n32940, n34869, n32947, n34853, n32946, n32951, n32949, n32948,
    n32950, n32955, n35720, n32953, n32952, n32954, n32956, n32957, n32959,
    n32958, n32961, n33073, n32965, n32963, n32962, n32964, n32982, n34990,
    n32972, n33619, n32970, n32971, n32973, n32980, n33944, n32974, n33866,
    n33758, n33529, n33759, n33615, n33077, n36411, n33947, n33867, n33761,
    n32977, n33080, n32978, n32979, n32981, n32984, n32983, n34013, n32988,
    n32987, n32989, n33023, n33021, n33141, n32991, n32990, n32995, n32993,
    n32992, n32994, n32999, n32997, n32996, n32998, n33019, n33001, n33000,
    n33005, n33003, n33002, n33004, n33013, n33007, n33006, n33011, n33009,
    n33008, n33010, n33012, n33017, n33015, n33014, n33016, n33018, n37322,
    n33020, n33022, n33025, n33024, n33060, n33058, n33027, n33026, n33030,
    n33028, n33029, n33032, n33031, n33036, n33034, n33033, n33035, n33056,
    n33038, n33037, n33042, n33040, n33039, n33041, n33050, n33044, n33043,
    n33048, n33046, n33045, n33047, n33049, n33054, n33052, n33051, n33053,
    n33055, n36400, n33057, n33059, n33065, n33061, n33266, n33063, n33064,
    n33069, n33068, n33070, n33072, n33071, n33087, n33076, n33075, n33672,
    n33131, n33085, n36412, n33078, n33079, n33119, n33117, n36460, n33081,
    n33082, n33083, n33084, n33086, n33089, n33088, n33092, n33091, n33093,
    n33097, n33096, n33098, n33102, n33100, n33099, n33101, n33103, n33105,
    n33104, n33110, n33108, n33871, n33888, n33107, n33109, n33115, n33111,
    n33112, n36915, n33113, n33114, n33135, n33118, n35849, n36436, n33120,
    n33121, n33122, n33130, n33123, n33128, n33126, n33125, n33127, n33129,
    n33133, n33132, n33134, n33137, n33136, n33138, n33162, n33164, n33145,
    n33140, n33143, n33142, n33144, n37584, n33836, n33146, n33147, n33151,
    n33149, n33148, n33150, n33161, n33153, n33152, n33159, n33154, n33822,
    n33156, n33157, n33158, n33160, n33167, n33165, n33166, n33205, n34329,
    n33171, n33170, n33175, n33173, n33172, n33174, n33201, n33177, n33176,
    n33181, n33179, n33178, n33180, n33189, n33183, n33182, n33187, n33185,
    n33184, n33186, n33188, n33199, n33190, n33195, n33193, n33192, n33194,
    n33197, n33196, n33198, n33200, n34328, n41065, n33203, n33202, n33204,
    n33211, n33207, n33209, n33210, n33215, n33213, n33212, n33214, n33220,
    n36003, n36004, n33218, n33219, n33224, n33223, n33229, n33226, n33227,
    n33228, n33231, n33230, n33235, n33233, n33232, n33234, n33243, n33237,
    n33236, n33241, n33239, n33238, n33240, n33242, n33259, n33245, n33244,
    n33249, n33247, n33246, n33248, n33257, n33251, n33250, n33255, n33253,
    n33252, n33254, n33256, n33258, n35458, n33265, n33261, n33263, n34401,
    n33264, n33270, n33267, n33269, n33274, n33272, n33271, n33273, n33308,
    n33276, n33275, n33280, n33278, n33277, n33279, n33306, n33282, n33281,
    n33286, n33284, n33283, n33285, n33294, n33288, n33287, n33292, n33290,
    n33289, n33291, n33293, n33304, n33296, n33295, n33300, n33297, n33299,
    n33302, n33301, n33303, n33305, n36174, n33307, n33312, n33311, n35869,
    n33319, n33316, n33315, n33317, n33318, n33321, n33320, n33322, n33356,
    n33354, n33324, n33323, n33328, n33326, n33325, n33327, n33336, n33330,
    n33329, n33334, n33332, n33331, n33333, n33335, n33352, n33338, n33337,
    n33342, n33340, n33339, n33341, n33350, n33344, n33343, n33348, n33346,
    n33345, n33347, n33349, n33351, n34965, n33353, n33355, n33544, n33359,
    n33358, n33361, n33360, n33363, n33362, n33365, n33364, n33367, n33366,
    n33369, n33368, n33371, n33370, n33373, n33372, n33375, n33374, n33377,
    n33376, n33379, n33378, n33381, n33380, n33383, n33382, n33385, n33384,
    n33387, n33386, n33389, n33388, n33391, n33390, n33393, n33392, n33395,
    n33394, n33397, n33396, n33399, n33398, n33401, n33400, n33403, n33402,
    n33405, n33404, n33407, n33406, n33409, n33408, n33411, n33410, n33413,
    n33412, n33415, n33414, n33417, n33416, n33419, n33418, n33421, n33420,
    n33423, n33422, n33425, n33427, n33426, n33429, n33431, n33430, n33433,
    n33435, n33434, n33437, n33439, n33438, n33441, n33443, n33442, n33445,
    n33447, n33446, n33449, n33451, n33450, n33453, n33455, n33454, n33457,
    n33459, n33458, n33461, n33463, n33462, n33465, n33467, n33466, n33469,
    n33471, n33470, n33473, n33476, n33475, n33478, n33484, n33479, n33482,
    n33483, n33485, n33493, n40743, n35893, n33491, n35902, n36914, n36975,
    n33489, n33490, n33492, n33495, n33494, n33499, n33497, n33930, n33498,
    n33511, n34615, n35613, n33506, n35924, n33503, n33504, n33505, n33509,
    n33508, n33510, n33513, n33512, n33526, n33517, n33521, n33519, n33518,
    n33520, n33522, n33524, n33523, n33525, n33536, n33534, n33528, n35986,
    n33530, n33531, n33532, n33533, n33535, n33541, n33539, n33538, n33540,
    n33543, n33542, n33547, n33546, n33550, n33549, n33552, n33551, n33554,
    n33553, n33558, n33557, n33560, n33559, n33562, n33561, n33565, n35784,
    n33574, n33568, n33566, n35782, n33567, n33572, n33570, n35785, n33571,
    n33573, n33576, n33575, n33578, n33592, n33584, n33581, n33580, n33582,
    n33583, n33590, n33587, n33586, n33588, n33589, n33591, n33593, n34877,
    n33595, n33599, n33597, n33603, n33596, n33598, n33610, n33820, n33600,
    n33608, n33605, n37749, n33604, n38154, n33606, n33607, n33609, n33614,
    n33611, n33612, n33613, n36070, n33616, n33617, n33618, n33635, n33629,
    n33624, n33623, n33625, n33627, n33626, n33628, n33633, n33631, n33632,
    n33634, n33637, n33636, n33653, n33638, n33645, n33640, n33639, n33641,
    n33643, n33642, n33644, n33651, n33649, n33648, n33650, n33652, n33660,
    n33678, n36212, n33654, n33696, n33655, n36181, n33656, n33657, n33658,
    n33659, n33665, n33663, n33664, n33677, n33668, n33667, n33670, n33669,
    n33671, n33675, n33673, n33862, n33674, n33676, n33684, n33679, n33844,
    n36216, n33680, n33681, n33682, n33683, n33687, n33685, n33686, n33704,
    n33690, n33689, n33692, n33691, n33693, n33702, n33694, n33697, n33695,
    n37096, n33698, n33699, n33700, n33701, n33703, n33708, n33706, n33753,
    n33707, n34070, n38058, n33713, n33712, n33729, n33715, n33722, n33723,
    n33728, n33730, n33732, n33735, n33737, n33736, n33752, n33744, n33740,
    n33742, n33743, n33745, n33750, n37090, n35845, n33746, n33747, n33748,
    n33749, n33751, n33755, n33754, n33780, n33760, n36026, n33762, n33763,
    n33776, n33768, n33767, n33769, n33774, n33771, n33773, n33775, n33778,
    n33777, n33779, n33782, n33781, n33788, n33785, n33787, n33790, n33789,
    n35503, n33798, n33796, n33795, n33797, n33800, n33799, n33812, n33808,
    n33806, n33804, n33803, n33805, n33807, n33810, n33809, n33811, n33818,
    n33813, n37760, n33815, n33816, n33817, n33834, n33830, n33828, n33826,
    n33825, n33827, n33829, n33832, n33831, n33833, n33841, n38178, n33837,
    n33838, n33839, n33840, n33843, n34526, n37700, n33845, n33846, n33847,
    n33861, n33855, n33850, n33849, n33851, n33853, n33852, n33854, n33859,
    n33857, n33858, n33860, n33864, n33863, n33865, n36968, n33868, n33869,
    n33887, n33877, n33875, n33874, n33876, n33885, n33883, n33878, n33879,
    n33881, n33880, n33882, n33884, n33886, n33890, n33889, n33893, n33914,
    n40733, n33896, n33897, n33895, n38913, n33898, n33899, n33912, n34624,
    n33901, n33905, n33903, n33902, n33904, n33910, n33908, n33907, n33909,
    n33911, n33913, n33916, n33920, n41172, n33919, n33922, n33921, n33924,
    n33931, n33929, n33927, n33926, n33928, n33942, n35905, n35914, n33932,
    n33940, n33934, n36058, n33938, n33936, n33935, n33937, n33939, n33941,
    n33950, n33943, n35926, n33946, n36670, n33948, n33949, n33952, n33957,
    n33955, n33954, n33956, n33969, n33959, n33958, n33960, n33967, n33961,
    n34976, n34978, n33962, n38037, n33963, n33964, n33965, n33966, n33968,
    n33973, n33971, n34999, n33972, n40055, n34007, n33975, n33974, n33979,
    n33977, n33976, n33978, n33983, n33981, n33980, n33982, n34003, n33985,
    n33984, n33989, n33987, n33986, n33988, n33997, n33991, n33990, n33995,
    n33993, n33992, n33994, n33996, n34001, n33999, n33998, n34000, n34002,
    n39500, n34005, n34004, n34006, n34010, n34008, n34009, n34015, n34012,
    n34014, n34019, n34017, n34016, n34018, n34052, n34021, n34020, n34025,
    n34023, n34022, n34024, n34050, n34027, n34026, n34031, n34029, n34028,
    n34030, n34039, n34033, n34032, n34037, n34035, n34034, n34036, n34038,
    n34048, n34041, n34040, n34044, n34772, n34043, n34046, n34045, n34047,
    n34049, n37918, n34051, n34278, n34054, n34053, n34062, n34056, n34282,
    n34060, n34059, n34061, n34065, n35884, n34064, n34067, n34066, n34069,
    n34068, n34072, n34111, n38050, n34073, n34079, n34077, n35475, n34717,
    n34075, n34089, n34076, n34596, n34078, n34087, n34249, n34081, n34248,
    n34080, n34125, n34736, n38132, n34085, n34083, n34082, n34731, n39888,
    n34084, n34086, n34096, n34092, n34091, n35185, n34093, n34095, n34098,
    n34100, n34099, n34108, n34102, n34101, n34106, n34104, n34103, n34105,
    n34107, n34110, n34109, n39298, n34112, n34118, n34116, n34113, n34114,
    n34126, n34115, n34360, n34117, n34123, n38123, n34121, n39383, n34120,
    n34122, n34133, n34128, n34127, n34129, n34130, n34132, n34135, n34138,
    n34137, n34146, n34140, n34139, n34144, n34142, n34141, n34143, n34145,
    n34148, n34147, n34150, n34153, n34152, n34161, n34155, n34154, n34159,
    n34157, n34156, n34158, n34160, n34163, n34162, n34168, n34167, n34176,
    n34170, n34169, n34174, n34172, n34171, n34173, n34175, n34178, n34177,
    n34180, n34179, n34184, n34182, n34181, n34183, n34186, n34185, n34191,
    n34190, n34199, n34193, n34192, n34197, n34195, n34194, n34196, n34198,
    n34201, n34200, n34203, n34202, n34207, n34205, n34204, n34206, n34209,
    n34208, n34211, n34210, n34215, n34213, n34212, n34214, n34217, n34216,
    n34219, n34218, n34223, n34221, n34220, n34222, n34225, n34224, n34227,
    n34230, n34229, n34238, n34232, n34231, n34236, n34234, n34233, n34235,
    n34237, n34240, n34239, n34245, n34244, n34255, n34247, n34246, n34253,
    n34251, n34250, n34252, n34254, n34257, n34256, n35021, n37474, n35010,
    n34263, n34261, n34409, n34259, n34264, n34260, n35011, n34262, n34274,
    n34266, n34265, n34267, n34268, n34272, n35032, n40037, n34271, n34273,
    n34276, n38889, n34275, n34277, n34297, n34281, n34280, n35364, n34294,
    n34284, n34289, n34288, n34292, n34291, n35365, n34293, n34295, n34296,
    n34333, n34299, n34298, n34303, n34301, n34300, n34302, n34311, n34305,
    n34304, n34309, n34307, n34306, n34308, n34310, n34327, n34313, n34312,
    n34317, n34315, n34314, n34316, n34325, n34319, n34318, n34323, n34321,
    n34320, n34322, n34324, n34326, n34764, n34763, n41388, n34331, n34330,
    n34332, n34338, n34334, n34336, n34806, n34337, n34342, n34341, n36119,
    n34347, n34345, n34346, n34349, n34348, n34353, n34352, n34359, n34354,
    n34357, n34849, n34847, n34358, n34362, n34361, n34367, n34365, n34364,
    n34366, n34369, n34368, n34371, n34370, n34375, n34373, n34372, n34374,
    n34379, n34377, n34376, n34378, n34399, n34381, n34380, n34385, n34383,
    n34382, n34384, n34393, n34387, n34386, n34391, n34389, n34388, n34390,
    n34392, n34397, n34395, n34394, n34396, n34398, n35308, n34407, n34403,
    n34405, n34406, n34408, n38397, n34749, n34415, n34420, n34413, n34411,
    n34410, n34412, n34414, n34419, n34737, n38469, n34417, n38557, n34416,
    n34418, n34427, n34424, n34422, n34423, n34426, n34429, n34428, n34433,
    n34431, n34430, n34432, n34435, n34434, n34437, n34436, n34441, n34439,
    n34438, n34440, n34443, n34442, n34445, n34444, n34449, n34447, n34446,
    n34448, n34451, n34450, n34453, n34452, n34457, n34455, n34454, n34456,
    n34459, n34458, n34461, n34460, n34465, n34463, n34462, n34464, n34467,
    n34466, n34469, n34468, n34473, n34471, n34470, n34472, n34475, n34474,
    n34494, n34483, n34481, n34479, n34480, n34482, n34484, n34488, n34486,
    n34487, n34491, n34490, n34492, n34493, n34506, n34497, n34501, n34500,
    n34504, n34503, n34510, n34516, n34519, n34520, n35622, n34525, n36872,
    n34527, n34528, n34529, n34544, n36874, n34530, n34542, n34533, n34532,
    n34535, n34534, n34540, n34538, n34537, n34539, n34541, n34543, n34549,
    n34983, n34548, n34556, n34554, n34579, n34553, n34555, n34557, n34559,
    n34558, n34561, n34562, n34564, n34563, n34565, n34567, n34566, n34568,
    n34571, n34570, n34572, n34574, n34573, n34577, n34578, n34582, n34581,
    n34583, n34587, n34586, n34589, n34588, n34593, n34591, n34590, n34592,
    n34595, n34594, n34598, n34597, n34603, n34601, n34600, n34602, n34605,
    n34604, n34608, n34607, n34610, n34609, n34613, n34612, n34619, n34614,
    n34617, n35907, n34616, n34618, n34621, n34620, n34623, n34622, n34636,
    n34661, n34628, n34630, n34627, n35523, n34664, n34629, n34634, n34632,
    n34631, n34633, n34635, n34644, n41158, n40725, n34639, n40724, n34640,
    n34642, n34643, n34647, n34648, n34650, n34649, n34654, n41707, n34653,
    n34658, n34657, n34670, n34660, n34663, n34662, n34668, n34666, n34665,
    n34667, n34669, n34676, n34672, n34674, n34675, n34678, n39028, n35152,
    n34681, n35179, n38478, n34680, n34698, n34683, n34692, n34686, n34688,
    n34690, n34689, n34696, n34694, n34693, n35156, n34695, n34697, n34700,
    n39107, n34699, n34702, n34701, n34706, n34704, n34703, n34705, n34708,
    n34707, n34710, n34709, n34714, n34712, n34711, n34713, n34716, n34715,
    n35350, n34724, n34719, n34720, n34722, n34721, n34723, n34735, n34727,
    n34729, n34728, n34733, n39374, n34732, n34734, n34739, n38562, n34738,
    n34741, n34740, n34745, n34743, n34742, n34744, n34747, n34746, n34751,
    n34750, n34756, n34754, n34753, n34755, n34758, n34757, n34762, n34760,
    n34759, n34761, n34805, n35588, n34765, n34770, n34769, n34777, n34771,
    n34775, n34774, n34776, n34781, n34779, n34778, n34780, n34801, n34783,
    n34782, n34787, n34785, n34784, n34786, n34795, n34789, n34788, n34793,
    n34791, n34790, n34792, n34794, n34799, n34797, n34796, n34798, n34800,
    n35587, n41680, n34803, n34802, n34804, n34811, n34807, n34809, n34810,
    n34828, n36104, n34816, n34822, n44014, n34820, n34819, n34821, n34826,
    n34824, n34825, n34827, n34834, n36982, n34832, n34831, n34833, n34839,
    n34837, n34838, n34841, n34840, n34846, n34845, n34852, n34848, n34850,
    n35456, n34851, n34855, n34854, n34873, n34868, n34856, n34857, n34862,
    n34860, n34861, n34866, n34864, n34865, n34867, n34871, n34870, n34872,
    n34875, n34874, n34878, n34893, n34882, n34881, n34883, n34884, n34891,
    n34887, n34886, n34888, n34889, n34890, n34892, n34895, n34894, n34897,
    n34896, n34900, n34899, n34905, n36599, n34904, n34911, n34907, n34908,
    n34910, n34912, n34916, n34915, n34919, n34922, n34921, n34924, n34923,
    n34926, n34925, n34930, n34928, n34927, n34929, n34932, n34931, n34934,
    n34933, n34938, n34936, n34935, n34937, n34940, n34939, n34942, n34941,
    n34946, n34944, n34943, n34945, n34948, n34947, n34950, n34949, n34954,
    n34952, n34951, n34953, n34956, n34955, n34958, n34957, n34962, n34960,
    n34959, n34961, n34964, n34963, n34973, n35309, n34970, n34971, n34972,
    n34975, n34974, n38031, n37011, n34977, n37010, n34980, n34981, n34982,
    n34998, n34984, n34994, n34988, n34987, n34989, n34992, n34991, n34993,
    n34996, n34995, n34997, n35001, n35000, n35003, n35002, n35007, n35005,
    n35004, n35006, n35009, n35008, n35013, n35012, n35018, n35016, n35015,
    n35017, n35020, n35019, n39805, n35022, n35088, n35027, n35025, n35023,
    n35024, n35026, n35031, n39879, n35029, n38894, n35028, n35030, n35039,
    n35036, n35034, n35035, n35037, n35038, n35041, n35040, n35045, n35043,
    n35042, n35044, n35047, n35046, n35049, n35048, n35053, n35051, n35050,
    n35052, n35055, n35054, n35057, n35056, n35061, n35059, n35058, n35060,
    n35063, n35062, n35065, n35064, n35069, n35067, n35066, n35068, n35071,
    n35070, n35073, n35072, n35077, n35075, n35074, n35076, n35079, n35078,
    n35081, n35080, n35085, n35083, n35082, n35084, n35087, n35086, n35091,
    n35090, n35095, n35093, n35092, n35094, n35098, n35097, n35103, n35101,
    n35102, n36120, n35107, n35689, n35105, n35106, n35119, n35111, n35117,
    n35115, n36129, n35114, n35116, n35118, n35121, n35120, n35125, n35123,
    n35122, n35124, n35127, n35126, n35129, n35128, n35133, n35131, n35130,
    n35132, n35135, n35134, n35137, n35136, n35141, n35139, n35138, n35140,
    n35143, n35142, n35145, n35144, n35149, n35147, n35146, n35148, n35151,
    n35150, n35154, n35153, n35160, n35158, n35157, n35159, n35162, n35161,
    n35164, n39938, n35166, n35236, n35171, n35169, n35167, n35168, n35170,
    n35177, n40048, n35175, n39102, n35174, n35176, n35187, n35183, n35181,
    n35182, n35184, n35186, n35189, n35188, n35193, n35191, n35190, n35192,
    n35195, n35194, n35197, n35196, n35201, n35199, n35198, n35200, n35203,
    n35202, n35205, n35204, n35209, n35207, n35206, n35208, n35211, n35210,
    n35213, n35212, n35217, n35215, n35214, n35216, n35219, n35218, n35221,
    n35220, n35225, n35223, n35222, n35224, n35227, n35226, n35229, n35228,
    n35233, n35231, n35230, n35232, n35235, n35234, n35239, n35238, n35243,
    n35241, n35240, n35242, n35246, n35245, n35248, n35247, n35252, n40565,
    n35251, n35257, n35255, n35256, n35260, n35258, n35259, n35264, n40943,
    n37339, n35263, n35266, n35265, n35271, n35269, n35610, n35268, n35270,
    n35272, n35274, n35273, n35276, n35275, n35280, n35278, n35277, n35279,
    n35282, n35281, n35284, n35283, n35288, n35286, n35285, n35287, n35290,
    n35289, n35292, n35291, n35296, n35294, n35293, n35295, n35298, n35297,
    n35300, n35299, n35304, n35302, n35301, n35303, n35306, n35305, n35698,
    n35313, n35311, n35310, n35312, n35315, n35314, n35319, n35318, n35320,
    n35328, n35333, n35337, n35370, n35335, n35336, n35341, n35339, n35338,
    n35340, n35343, n35342, n35347, n35345, n35344, n35346, n35349, n35348,
    n35353, n35352, n35358, n35356, n35355, n35357, n35360, n35359, n35362,
    n35375, n35373, n35369, n35367, n35368, n35371, n35372, n35374, n35383,
    n35379, n35382, n35385, n35384, n35387, n35386, n35391, n35389, n35388,
    n35390, n35418, n35394, n35393, n35398, n35396, n35395, n35397, n35406,
    n35400, n35399, n35404, n35402, n35401, n35403, n35405, n35416, n35410,
    n35409, n35414, n35412, n35411, n35413, n35415, n35417, n35691, n35424,
    n35419, n35422, n35423, n35427, n35428, n35430, n35429, n35434, n35433,
    n36527, n37089, n35441, n35438, n36515, n35440, n35450, n35444, n37753,
    n35448, n36516, n35447, n35449, n35451, n35454, n40731, n41400, n35923,
    n35925, n35910, n35453, n35455, n35457, n35461, n35460, n35464, n35463,
    n35467, n35481, n35469, n35479, n35472, n35471, n35477, n36135, n35476,
    n35478, n35480, n35483, n35482, n35491, n35487, n35486, n35489, n35488,
    n35490, n35499, n35497, n35493, n35492, n35495, n36141, n35496, n35498,
    n35516, n35511, n36107, n35510, n35506, n35504, n35505, n35508, n35507,
    n35509, n35514, n35878, n35513, n35522, n35520, n35519, n35521, n35524,
    n35949, n35547, n41682, n35540, n35526, n35528, n35538, n35530, n35531,
    n40864, n35535, n35533, n35536, n35537, n35539, n35545, n35640, n35544,
    n35549, n35548, n35556, n35552, n35554, n35592, n35558, n35557, n35562,
    n35560, n35559, n35561, n35570, n35564, n35563, n35568, n35566, n35565,
    n35567, n35569, n35586, n35572, n35571, n35576, n35574, n35573, n35575,
    n35584, n35578, n35577, n35582, n35580, n35579, n35581, n35583, n35585,
    n36330, n36329, n41862, n35590, n35589, n35591, n35597, n35593, n35595,
    n35596, n35600, n35605, n35603, n35604, n35607, n35606, n35612, n35611,
    n35615, n35614, n35618, n35671, n35616, n35672, n35617, n35619, n35621,
    n35620, n35625, n35639, n35637, n35628, n35629, n35635, n35632, n35633,
    n35634, n35636, n35638, n35653, n35643, n35943, n35960, n35651, n35649,
    n35647, n35646, n35648, n35650, n35652, n35661, n41096, n41099, n35655,
    n41105, n35657, n35659, n35662, n35906, n35669, n35664, n35665, n35666,
    n35668, n35674, n35673, n35677, n35675, n35676, n35678, n35680, n35679,
    n35688, n35684, n35683, n35686, n35685, n35690, n35693, n35692, n35704,
    n35696, n35702, n35699, n35700, n35701, n35703, n35706, n35705, n35713,
    n35710, n35712, n36358, n35717, n35716, n35736, n35734, n35723, n35727,
    n35724, n35726, n35732, n35730, n35731, n35733, n36497, n35735, n35748,
    n35737, n35739, n35741, n35743, n35746, n35745, n35747, n35779, n35768,
    n35761, n35764, n35760, n35754, n35753, n35758, n35757, n35759, n36531,
    n35762, n35763, n35765, n35767, n35770, n35773, n35775, n35776, n35783,
    n35794, n35789, n35787, n35786, n35788, n35792, n35791, n35793, n35799,
    n35795, n35797, n35798, n35810, n35803, n36360, n35808, n35807, n35809,
    n35818, n35813, n35812, n35814, n35815, n35817, n35827, n35825, n35824,
    n36981, n35826, n35829, n35828, n36263, n35830, n35839, n35837, n35835,
    n35834, n40961, n40969, n36447, n40387, n35841, n35840, n35855, n36068,
    n36434, n35851, n35844, n35843, n37092, n35848, n35846, n40406, n35847,
    n35853, n35850, n37094, n35852, n35854, n35868, n40377, n35857, n35856,
    n35866, n40857, n35860, n35862, n35864, n35863, n40378, n35865, n35867,
    n35872, n35871, n35874, n35873, n35888, n35876, n35882, n35880, n35879,
    n35881, n35886, n35883, n35885, n35890, n35892, n35898, n35895, n35894,
    n35896, n36342, n35897, n35899, n35901, n35900, n35903, n35934, n35909,
    n35908, n35913, n35911, n35912, n35915, n35922, n35920, n35919, n35921,
    n35932, n35928, n35927, n35929, n35931, n35933, n35937, n35936, n35938,
    n41519, n35946, n35957, n35955, n35948, n35953, n36157, n35950, n36171,
    n35952, n35954, n35956, n42130, n35961, n35965, n35966, n35969, n35968,
    n35973, n40620, n35972, n36345, n35978, n36346, n35977, n35985, n41098,
    n35983, n36353, n35981, n35980, n35982, n35984, n40280, n35987, n35994,
    n40260, n40263, n35992, n35990, n40261, n35991, n35993, n36000, n35996,
    n36031, n36034, n35998, n36066, n35999, n36012, n36006, n36005, n36947,
    n36948, n38815, n36946, n36007, n36008, n36010, n36009, n36014, n36013,
    n36016, n36015, n36018, n36017, n40208, n36030, n40201, n36025, n36023,
    n40193, n36024, n36028, n36027, n36029, n36037, n36033, n36032, n36035,
    n36036, n36044, n36056, n36051, n36050, n36053, n36054, n36060, n36059,
    n36062, n36065, n36064, n39638, n36074, n36067, n36069, n36072, n36071,
    n36073, n36085, n36076, n39616, n36083, n36081, n36079, n39618, n36080,
    n36082, n36084, n36098, n36087, n36089, n36121, n36094, n36093, n36096,
    n36095, n36124, n36102, n36100, n36101, n36106, n36105, n36108, n36114,
    n36112, n36111, n36113, n36117, n36127, n36123, n36130, n36132, n36140,
    n36134, n36133, n36138, n36137, n36139, n36142, n36148, n36146, n36145,
    n36147, n36151, n36156, n36155, n36170, n36160, n36166, n36163, n36165,
    n36172, n36180, n36175, n36178, n36189, n40150, n36185, n36183, n36214,
    n36184, n36187, n36186, n36188, n36201, n40144, n36199, n36191, n36194,
    n40134, n36197, n40135, n36196, n36198, n36200, n36204, n36208, n36207,
    n36210, n36209, n36226, n36213, n36215, n37696, n36219, n36217, n40235,
    n36218, n36224, n36221, n37698, n36223, n36225, n36236, n40339, n36228,
    n40214, n36229, n36234, n36231, n40216, n36232, n36233, n36235, n36238,
    n36241, n41481, n36240, n36247, n36244, n36245, n36246, n36252, n36250,
    n36251, n36254, n36256, n36255, n36260, n40368, n36259, n36262, n36261,
    n36268, n36266, n36265, n36267, n36271, n36270, n36275, n36277, n36276,
    n36278, n36337, n36285, n36284, n36335, n36288, n36287, n36293, n36291,
    n36290, n36292, n36305, n36297, n36296, n36303, n36301, n36300, n36302,
    n36304, n36328, n36309, n36308, n36315, n36313, n36312, n36314, n36326,
    n36319, n36318, n36324, n36322, n36321, n36323, n36325, n36327, n36332,
    n36331, n42134, n36334, n36336, n36340, n36339, n36341, n36344, n36343,
    n36350, n36348, n36347, n36349, n36351, n36356, n36354, n36355, n36361,
    n36362, n36372, n36367, n36368, n36369, n36371, n36394, n36378, n36379,
    n36389, n36383, n36381, n36382, n36387, n36386, n36388, n36392, n36391,
    n36397, n36406, n36402, n36404, n36408, n36407, n36410, n36409, n36426,
    n36414, n36413, n36419, n40463, n37748, n36462, n36416, n36465, n36417,
    n36418, n36424, n36421, n36420, n36422, n36423, n36425, n36432, n36428,
    n36430, n40455, n36431, n36435, n36443, n40987, n36437, n36441, n36463,
    n36438, n36440, n36442, n36454, n36470, n36445, n36449, n36471, n36448,
    n36450, n40979, n36452, n37086, n36451, n36453, n36458, n36456, n36455,
    n36457, n40513, n36478, n40519, n36461, n36469, n36464, n36467, n36466,
    n36468, n36476, n36473, n36472, n36474, n40510, n36475, n36477, n36481,
    n36480, n36484, n36604, n36482, n36483, n36496, n36494, n36851, n36491,
    n36495, n36499, n36498, n36505, n36537, n37315, n36503, n36502, n36536,
    n36504, n36506, n36508, n36507, n36510, n36514, n40445, n40247, n36511,
    n36512, n36513, n36524, n40384, n36522, n36518, n36517, n36520, n38598,
    n36521, n36523, n36525, n36530, n36528, n36529, n36535, n36534, n36540,
    n36538, n36539, n36541, n36545, n36544, n36551, n36548, n36549, n36550,
    n36555, n36554, n36577, n39021, n36802, n36803, n36564, n36778, n37132,
    n37610, n36563, n36585, n38235, n36566, n36567, n36583, n36570, n36571,
    n36572, n36576, n36573, n36581, n39233, n36580, n36582, n36584, n36589,
    n39601, n36588, n36598, n36596, n36594, n39606, n36593, n36595, n36597,
    n36611, n36603, n36602, n36841, n36606, n36605, n36609, n36608, n36610,
    n36619, n36617, n36614, n36618, n36623, n36622, n36631, n36629, n36627,
    n39542, n36626, n36628, n36630, n39244, n36647, n37944, n36651, n36636,
    n36639, n36637, n36638, n36641, n36640, n36645, n38773, n39517, n36644,
    n36646, n36658, n36649, n36650, n36655, n36657, n36962, n36917, n36662,
    n36663, n36674, n38724, n36669, n38723, n36668, n36672, n36671, n36675,
    n38735, n39153, n36681, n39156, n36679, n36678, n36687, n36685, n36684,
    n36686, n36690, n36689, n36700, n39201, n36698, n36696, n36695, n36699,
    n36702, n36701, n36708, n36706, n36704, n36703, n36707, n36710, n36709,
    n36716, n36714, n36712, n36711, n36715, n36718, n36717, n36724, n36722,
    n36720, n36719, n36721, n36723, n36726, n36725, n36732, n36730, n36728,
    n36727, n36731, n36743, n36733, n36734, n36735, n36739, n36741, n36740,
    n36742, n36753, n36751, n36747, n36748, n36750, n36752, n36757, n36755,
    n40886, n36754, n36756, n36761, n36759, n36758, n36760, n36765, n36763,
    n36762, n36764, n36769, n36767, n36766, n36768, n36773, n36771, n36770,
    n36772, n36777, n36775, n36774, n36776, n36781, n39268, n36780, n36791,
    n39271, n36789, n36787, n38678, n36786, n36790, n36798, n36797, n36811,
    n39285, n36809, n36807, n38669, n36806, n36810, n36815, n36813, n36812,
    n36814, n36819, n36817, n36816, n36818, n36821, n36820, n36827, n36825,
    n36823, n36822, n36824, n36826, n40354, n36837, n40559, n36832, n36953,
    n36833, n36835, n36834, n36836, n36839, n36838, n36843, n39658, n36842,
    n36850, n36845, n37558, n36844, n36848, n36847, n36849, n36865, n36856,
    n36855, n36858, n36863, n36864, n37706, n36870, n36884, n39392, n36881,
    n36879, n36875, n36877, n36876, n37012, n36878, n36880, n36882, n39418,
    n36883, n36888, n36886, n36899, n36892, n36897, n36896, n39559, n36898,
    n36912, n36903, n36902, n36910, n37496, n36907, n40183, n36926, n36923,
    n36916, n36964, n36919, n36921, n36920, n36922, n36924, n40189, n36925,
    n36929, n40180, n36928, n36933, n36931, n41311, n36930, n36932, n36937,
    n36935, n36934, n36936, n36941, n36939, n36938, n36945, n36943, n36942,
    n36944, n36959, n36949, n36951, n36950, n36952, n36954, n36956, n36961,
    n36960, n36965, n36980, n38590, n36972, n38593, n36971, n36977, n38592,
    n36976, n36979, n36989, n37238, n36985, n36983, n36984, n36987, n36986,
    n36988, n36999, n36997, n36995, n36994, n36996, n36998, n37005, n37008,
    n37020, n37013, n38033, n37015, n39459, n37014, n37018, n38035, n37017,
    n37019, n37029, n37027, n37022, n38142, n38208, n37032, n37030, n37076,
    n37031, n37051, n37034, n37035, n37036, n37049, n37040, n37041, n37042,
    n37047, n37046, n37050, n37053, n37052, n37059, n37057, n37055, n37054,
    n37058, n37061, n37060, n37067, n37065, n37063, n37062, n37066, n37069,
    n37068, n37075, n37073, n37071, n37070, n37074, n37078, n37077, n37084,
    n37082, n37080, n37079, n37083, n40962, n37105, n37087, n37103, n40956,
    n38155, n37091, n37093, n37100, n37095, n37098, n37097, n37099, n37101,
    n37102, n37104, n37111, n37109, n37108, n37110, n37114, n37113, n37118,
    n37116, n37115, n37117, n37129, n37122, n37127, n37125, n37126, n39193,
    n37134, n39123, n37202, n37133, n37153, n37135, n37136, n37137, n37151,
    n37140, n37141, n37142, n37146, n37149, n37148, n37155, n37154, n37161,
    n37159, n37157, n37156, n37163, n37162, n37169, n37167, n37165, n37164,
    n37171, n37170, n37177, n37175, n37173, n37172, n37179, n37178, n37185,
    n37183, n37181, n37180, n37187, n37186, n37193, n37191, n37189, n37188,
    n37195, n37194, n37201, n37199, n37197, n37196, n37204, n37203, n37212,
    n37210, n37208, n37207, n37216, n37217, n44008, n37222, n37221, n37223,
    n37225, n37224, n37232, n37226, n37229, n37230, n37231, n37233, n37236,
    n37240, n37239, n37255, n37253, n37244, n37249, n37247, n37248, n37250,
    n37257, n37256, n37263, n37258, n37259, n37261, n37260, n37262, n37268,
    n37266, n37276, n37284, n37282, n37281, n37283, n37301, n37299, n37287,
    n37295, n37293, n37291, n37292, n37294, n37297, n37296, n37298, n37300,
    n37307, n37305, n37304, n37306, n37321, n37319, n37309, n37308, n37314,
    n37312, n37311, n37313, n37317, n37316, n37318, n37320, n37328, n37323,
    n37326, n37921, n37331, n37330, n37333, n37332, n37334, n37336, n37335,
    n37337, n37347, n37345, n37343, n37340, n37341, n37342, n37344, n37346,
    n37348, n37350, n37354, n37353, n37358, n37357, n37375, n37371, n37369,
    n37361, n37609, n38778, n37381, n37377, n37378, n37380, n37387, n37385,
    n37389, n37388, n37395, n37393, n37397, n37396, n37405, n37401, n37400,
    n37403, n37402, n37413, n37409, n37408, n37411, n37410, n37415, n37422,
    n37418, n37417, n37420, n37419, n37431, n37427, n37426, n37429, n37428,
    n37432, n37436, n37435, n37440, n37438, n37437, n37439, n37449, n37443,
    n37447, n37446, n37451, n37450, n37458, n37453, n37454, n37456, n37455,
    n37457, n37463, n37462, n37465, n42723, n37471, n37480, n38057, n39819,
    n38062, n37478, n37477, n37479, n37484, n37482, n37481, n37483, n37495,
    n39956, n37497, n37506, n37504, n37510, n37522, n37514, n37512, n37511,
    n37513, n37515, n37518, n37517, n37528, n37524, n37523, n37526, n37525,
    n39646, n37534, n37533, n37538, n37546, n37541, n37540, n37544, n37543,
    n37548, n37553, n37552, n37554, n37565, n37559, n37560, n37562, n37566,
    n40470, n37576, n37582, n37579, n37581, n37580, n38156, n37586, n38157,
    n37583, n37585, n37587, n37592, n37603, n37599, n37598, n37601, n37600,
    n39548, n37607, n38323, n37611, n37613, n37614, n37617, n37616, n37619,
    n37618, n37622, n37632, n37636, n37649, n37647, n37646, n37661, n37659,
    n37652, n37653, n37655, n37656, n37658, n37660, n37663, n37662, n37669,
    n37667, n37665, n37664, n37666, n37668, n37671, n37670, n37677, n37675,
    n37673, n37672, n37674, n37676, n37679, n37678, n37685, n37683, n37681,
    n37680, n37682, n37684, n37687, n37686, n37693, n37691, n37689, n37688,
    n37690, n37692, n37695, n37697, n37705, n37699, n37703, n37701, n40348,
    n37702, n37704, n37708, n37707, n37712, n37709, n37711, n37715, n37714,
    n37719, n37718, n37734, n37722, n37720, n37721, n37724, n37723, n37737,
    n37741, n37740, n37742, n37746, n37770, n37751, n37750, n37752, n38918,
    n37755, n37756, n37764, n40237, n37762, n38917, n37759, n37761, n37763,
    n37768, n37771, n37773, n37775, n37785, n37781, n37780, n37786, n37793,
    n37789, n37788, n37794, n37802, n37798, n37797, n37803, n37812, n37807,
    n37806, n37813, n37820, n37816, n37815, n37821, n37824, n37823, n37826,
    n37829, n37828, n37833, n37832, n37843, n37838, n37837, n37844, n37847,
    n37849, n37865, n37863, n38324, n37950, n37866, n37869, n37875, n37867,
    n37871, n37872, n37874, n37881, n37879, n37883, n37882, n37889, n37887,
    n37891, n37890, n37897, n37895, n37899, n37898, n37907, n37903, n37902,
    n37905, n37904, n37908, n37915, n37911, n37910, n37913, n37912, n37916,
    n37924, n37920, n39503, n37923, n37928, n37926, n37930, n37929, n37940,
    n37936, n37935, n37938, n37937, n37943, n37942, n37960, n37958, n37961,
    n37964, n37954, n37970, n37962, n37966, n37967, n37969, n37974, n37973,
    n37980, n37978, n37975, n37982, n37981, n37988, n37986, n37983, n37990,
    n37989, n37996, n37994, n37991, n37998, n37997, n38004, n38002, n37999,
    n38006, n38005, n38012, n38010, n38007, n38026, n38017, n38022, n38020,
    n38019, n38021, n38024, n38023, n38025, n38046, n38032, n38034, n38041,
    n38036, n38039, n38038, n38040, n38042, n40434, n38122, n38052, n38051,
    n38071, n38055, n38060, n38067, n38065, n38072, n38075, n38074, n38079,
    n38080, n38083, n38082, n38087, n38088, n38091, n38090, n38095, n38096,
    n38099, n38098, n38103, n38104, n38107, n38106, n38111, n38112, n38115,
    n38114, n38119, n38120, n38125, n38124, n38131, n38133, n38137, n38136,
    n38180, n38141, n38166, n38145, n38146, n38162, n38179, n38158, n38171,
    n38159, n38160, n39803, n38161, n38163, n38187, n40533, n38183, n40540,
    n38181, n38182, n38184, n38196, n38192, n38191, n38193, n38204, n38200,
    n38199, n38201, n38216, n38211, n38210, n38213, n38234, n38230, n38225,
    n38224, n38226, n38227, n39019, n38229, n38231, n38240, n38250, n38246,
    n38245, n38247, n38255, n38254, n38264, n38257, n38259, n38258, n38260,
    n38262, n38261, n38263, n38268, n38265, n38274, n38270, n38269, n38271,
    n38278, n38617, n38293, n39278, n38289, n38284, n38283, n38285, n38286,
    n38288, n38290, n38299, n38312, n38308, n38307, n38309, n38318, n38332,
    n38317, n38344, n38335, n38326, n38327, n39603, n38342, n38333, n38338,
    n38339, n38346, n38345, n38352, n38350, n38347, n38354, n38353, n38360,
    n38358, n38355, n38362, n38361, n38368, n38366, n38363, n38371, n39653,
    n38369, n38370, n38382, n38375, n39652, n38380, n38378, n38387, n38386,
    n38391, n38390, n38660, n38392, n38393, n38468, n38399, n38398, n38417,
    n38400, n38404, n38405, n38408, n39957, n39954, n38413, n38418, n38421,
    n38420, n38425, n38426, n38429, n38428, n38433, n38434, n38437, n38436,
    n38441, n38442, n38445, n38444, n38449, n38450, n38453, n38452, n38457,
    n38458, n38461, n38460, n38465, n38466, n38471, n38470, n38477, n38479,
    n38483, n38552, n38488, n39029, n38486, n38485, n38487, n38501, n38496,
    n39041, n38498, n38503, n38502, n38505, n38504, n38509, n38506, n38511,
    n38510, n38513, n38512, n38517, n38514, n38519, n38518, n38521, n38520,
    n38525, n38522, n38527, n38526, n38529, n38528, n38533, n38530, n38535,
    n38534, n38537, n38536, n38541, n38538, n38543, n38542, n38545, n38544,
    n38549, n38546, n38551, n38550, n38555, n38554, n38561, n38558, n38564,
    n38563, n38568, n38566, n38570, n38576, n38574, n38578, n38584, n38582,
    n38586, n38591, n38611, n40262, n38608, n38606, n38596, n38604, n38601,
    n40175, n38600, n38597, n38599, n38722, n38602, n38603, n38607, n38624,
    n38613, n38627, n38622, n38621, n38633, n38629, n38630, n38632, n38634,
    n38637, n38639, n38646, n38644, n38658, n38656, n38647, n38649, n38651,
    n38654, n38653, n38655, n39641, n38657, n38666, n38663, n38668, n38667,
    n38675, n38673, n38671, n38670, n38677, n38676, n38684, n38682, n38680,
    n38679, n38686, n38685, n38693, n38691, n38689, n38688, n38695, n38694,
    n38702, n38700, n38698, n38697, n38705, n38704, n38712, n38710, n38708,
    n38707, n38714, n38713, n38721, n38719, n38717, n38716, n38730, n38726,
    n38725, n38728, n38727, n38729, n38734, n38733, n38736, n38742, n38738,
    n38737, n38739, n38750, n38746, n38745, n38747, n38758, n38754, n38753,
    n38755, n38766, n38762, n38761, n38763, n38777, n38772, n38771, n38774,
    n38782, n38789, n38784, n38783, n38785, n38787, n38786, n38788, n38797,
    n38795, n38793, n38800, n39558, n38805, n38811, n38809, n38819, n38817,
    n38816, n38818, n38827, n38825, n38823, n38822, n38824, n38826, n38830,
    n38831, n38832, n38834, n38837, n38836, n38841, n38838, n38842, n38845,
    n38844, n38849, n38846, n38850, n38853, n38852, n38857, n38854, n38858,
    n38861, n38860, n38865, n38862, n38866, n38869, n38868, n38873, n38870,
    n38874, n38877, n38876, n38881, n38878, n38882, n38887, n38886, n38893,
    n38890, n38895, n38900, n38899, n38908, n38912, n39427, n38911, n38916,
    n38914, n40845, n38915, n38920, n39428, n38919, n38921, n38926, n38937,
    n38932, n38931, n38935, n38934, n38942, n38943, n38957, n38953, n38944,
    n38949, n38947, n38946, n38948, n38951, n38950, n38952, n38955, n38954,
    n38958, n38963, n38961, n38965, n38964, n38971, n38976, n38974, n38973,
    n38975, n38978, n38977, n38979, n38986, n38984, n38988, n38987, n38992,
    n38991, n38998, n38996, n38993, n39000, n38999, n39006, n39004, n39001,
    n39008, n39007, n39014, n39012, n39009, n39018, n39017, n39027, n39025,
    n39022, n39034, n39032, n39031, n39033, n39046, n39043, n39047, n39050,
    n39049, n39054, n39051, n39055, n39058, n39057, n39062, n39059, n39063,
    n39066, n39065, n39070, n39067, n39071, n39074, n39073, n39078, n39075,
    n39079, n39082, n39081, n39086, n39083, n39087, n39090, n39089, n39094,
    n39091, n39095, n39100, n39099, n39106, n39103, n39108, n39115, n39117,
    n39116, n39118, n39191, n39122, n39121, n39132, n39128, n39131, n39135,
    n39138, n39137, n39144, n39140, n39146, n39145, n39152, n39148, n39155,
    n39154, n39162, n39160, n39158, n39164, n39163, n39170, n39166, n39172,
    n39171, n39178, n39174, n39180, n39179, n39186, n39182, n39190, n39189,
    n39199, n39195, n39205, n39207, n39206, n39213, n39212, n39215, n39214,
    n39216, n39220, n39218, n39217, n39219, n39229, n39227, n39225, n39221,
    n39223, n39224, n39226, n39232, n39231, n39239, n39237, n39234, n39243,
    n39242, n39250, n39248, n39245, n39253, n39252, n39259, n39257, n39254,
    n39261, n39260, n39267, n39265, n39262, n39270, n39269, n39277, n39275,
    n39272, n39282, n39281, n39292, n39290, n39287, n39294, n39373, n39300,
    n39299, n39322, n39306, n39305, n39308, n39314, n39816, n39312, n39820,
    n39318, n39317, n39319, n39323, n39326, n39325, n39330, n39327, n39331,
    n39334, n39333, n39338, n39335, n39339, n39342, n39341, n39346, n39343,
    n39347, n39350, n39349, n39354, n39351, n39355, n39358, n39357, n39362,
    n39359, n39363, n39366, n39365, n39370, n39367, n39371, n39376, n39375,
    n39382, n39379, n39384, n40222, n40212, n39391, n39403, n39402, n39406,
    n39397, n39396, n39400, n40126, n39399, n40124, n40226, n39407, n39408,
    n39416, n41017, n39436, n39421, n39432, n39430, n39429, n39431, n39433,
    n39458, n39441, n39443, n39463, n39462, n39465, n39464, n39466, n39468,
    n39467, n39469, n39479, n39477, n39475, n39472, n39473, n39474, n39476,
    n39478, n39484, n39483, n39486, n39485, n39487, n39489, n39488, n39490,
    n39499, n39497, n39495, n39492, n39493, n39494, n39496, n39498, n39506,
    n39501, n39512, n39513, n39521, n39519, n39518, n39520, n39539, n39533,
    n39537, n39536, n39538, n39547, n39545, n39544, n39546, n39553, n39551,
    n39550, n39552, n39554, n39556, n39568, n39566, n39561, n39570, n39582,
    n39572, n39577, n39575, n39574, n39576, n39580, n39579, n39581, n39584,
    n39644, n39591, n39597, n39595, n39611, n39605, n39604, n39608, n39637,
    n39617, n39634, n39632, n39619, n39621, n39630, n39623, n39628, n39625,
    n40444, n40267, n39626, n40505, n40446, n39627, n39629, n39639, n39642,
    n39650, n39647, n39666, n39662, n39655, n39654, n39660, n39657, n39659,
    n39661, n39664, n39663, n39674, n39679, n39677, n39676, n39678, n39681,
    n39680, n39682, n39687, n39686, n39690, n39692, n39691, n39697, n39694,
    n39695, n39696, n39699, n39698, n39706, n39705, n39711, n39714, n39720,
    n39718, n39719, n39726, n39724, n39723, n39725, n39729, n39728, n39731,
    n39730, n39736, n39734, n39733, n39735, n39739, n39738, n39746, n39742,
    n39748, n39747, n39755, n39750, n39751, n39753, n39752, n39760, n43225,
    n39766, n39778, n39777, n39779, n40240, n40523, n39781, n39784, n40821,
    n39782, n39783, n39793, n39787, n39791, n39800, n39801, n39878, n39807,
    n39806, n39827, n39812, n39813, n39823, n39822, n39824, n39828, n39831,
    n39830, n39835, n39832, n39836, n39839, n39838, n39843, n39840, n39844,
    n39847, n39846, n39851, n39848, n39852, n39855, n39854, n39859, n39856,
    n39860, n39863, n39862, n39867, n39864, n39868, n39871, n39870, n39875,
    n39872, n39876, n39881, n39880, n39887, n39884, n39889, n39893, n39899,
    n39900, n39897, n39898, n39906, n39902, n39904, n39903, n39905, n39908,
    n39912, n39911, n39919, n39914, n39915, n39917, n39916, n39918, n39924,
    n39923, n39933, n39932, n39949, n40036, n39941, n39940, n39966, n39950,
    n39961, n39960, n39963, n39968, n39972, n39971, n39977, n39974, n39979,
    n39983, n39982, n39988, n39985, n39990, n39994, n39993, n39999, n39996,
    n40001, n40005, n40004, n40010, n40007, n40012, n40016, n40015, n40021,
    n40018, n40023, n40027, n40026, n40032, n40029, n40034, n40040, n40039,
    n40047, n40044, n40050, n40060, n40058, n40057, n40059, n40062, n40061,
    n40063, n40068, n40087, n40077, n40075, n40074, n42982, n40076, n40083,
    n40082, n40084, n40090, n40487, n40104, n40102, n40095, n40106, n40105,
    n40111, n40108, n40109, n40110, n40113, n40112, n40117, n40116, n40122,
    n40149, n40965, n40131, n40967, n40129, n40128, n40393, n40130, n40133,
    n40139, n40137, n40136, n40138, n40143, n40140, n40145, n40165, n40163,
    n40156, n40155, n40161, n40158, n40160, n40162, n40188, n40171, n40169,
    n40174, n40172, n40173, n40178, n40176, n40177, n40181, n40184, n40187,
    n40190, n40207, n40192, n40198, n40195, n40197, n40199, n40203, n40206,
    n40209, n40338, n40220, n40329, n40218, n40330, n40217, n40219, n40228,
    n40224, n40223, n40225, n40227, n40230, n40233, n40238, n40259, n40250,
    n40246, n40832, n41004, n40252, n40279, n40265, n40264, n40276, n40266,
    n40268, n40274, n40272, n40273, n40281, n40284, n40283, n40287, n40286,
    n40288, n40292, n40290, n40289, n40291, n40305, n40295, n40297, n40303,
    n40301, n40300, n40302, n40304, n40310, n40308, n40307, n40309, n40318,
    n40316, n40314, n40313, n40315, n40317, n40321, n40322, n40323, n40326,
    n40328, n40333, n40332, n40334, n40337, n40336, n40340, n40342, n40343,
    n40346, n40353, n40351, n40352, n40361, n40359, n40357, n40356, n40358,
    n40360, n40364, n40365, n40366, n40370, n40369, n40380, n40379, n40381,
    n40399, n40386, n40383, n40385, n40499, n40397, n40396, n40392, n40390,
    n40391, n40394, n40413, n40416, n40419, n40420, n40424, n40423, n40473,
    n40426, n40432, n40438, n40437, n40440, n40439, n40450, n40498, n40448,
    n40447, n40449, n40453, n40452, n40454, n40457, n40456, n40458, n40461,
    n40472, n40477, n40474, n40489, n40488, n40492, n40491, n40495, n40518,
    n40502, n40501, n40507, n40504, n40506, n40990, n40988, n40509, n40512,
    n40511, n40514, n40522, n40525, n40548, n40543, n41058, n40552, n40551,
    n40556, n40554, n40553, n40555, n40557, n40563, n40561, n40560, n40562,
    n40564, n40569, n40567, n40566, n40568, n40571, n40575, n40576, n40577,
    n40581, n40599, n40595, n40583, n40591, n40584, n40585, n40589, n40588,
    n40590, n40593, n40592, n40594, n40597, n40596, n40600, n40619, n40615,
    n40603, n40611, n40604, n40605, n40609, n40608, n40610, n40613, n40612,
    n40614, n40617, n40616, n40621, n40642, n40638, n40623, n40634, n40628,
    n40627, n40632, n40631, n40633, n40636, n40635, n40637, n40640, n40639,
    n40643, n40664, n40660, n40645, n40656, n40650, n40649, n40654, n40653,
    n40655, n40658, n40657, n40659, n40662, n40661, n40665, n40688, n40684,
    n40667, n40680, n40674, n40673, n40678, n40677, n40679, n40682, n40681,
    n40683, n40686, n40685, n40689, n40690, n40701, n40699, n40694, n40697,
    n40696, n40698, n40702, n40722, n40705, n40720, n40714, n40712, n40710,
    n40711, n40713, n40730, n40728, n40870, n40727, n40729, n40742, n40737,
    n40735, n40736, n40871, n40739, n40740, n40741, n40756, n40749, n40764,
    n40761, n40763, n40942, n40944, n40774, n40768, n41069, n40772, n41068,
    n40771, n40773, n40777, n40776, n40779, n40778, n40780, n40792, n40785,
    n40788, n40787, n40790, n40789, n40794, n40801, n40799, n40800, n40808,
    n40814, n40811, n41390, n40822, n40826, n40825, n40827, n40837, n40828,
    n40829, n40834, n40831, n40833, n40835, n40849, n40867, n41260, n40866,
    n40868, n40878, n41157, n40874, n41159, n40873, n40876, n40875, n40877,
    n40890, n40885, n40884, n40888, n40887, n40903, n40898, n40897, n40901,
    n40900, n40905, n40915, n40910, n40909, n40913, n40912, n40917, n40919,
    n40920, n40940, n40922, n40924, n43196, n40930, n40928, n40927, n40929,
    n40931, n40938, n40947, n40945, n40946, n40951, n40949, n40950, n40952,
    n40957, n40978, n40975, n40966, n40971, n40970, n40984, n40996, n40989,
    n40991, n40995, n41001, n41000, n41007, n41038, n41021, n41036, n41032,
    n41028, n41026, n41027, n41029, n41042, n41041, n41046, n41044, n41043,
    n41045, n41047, n41057, n41051, n41050, n41055, n41053, n41052, n41054,
    n41056, n41061, n41060, n41062, n41066, n41071, n41070, n41075, n41074,
    n41090, n41080, n41086, n41082, n41178, n41084, n41083, n41085, n41094,
    n41097, n41103, n41404, n41102, n41101, n41417, n41110, n41108, n41418,
    n41106, n41107, n41109, n41116, n41144, n41126, n41142, n41138, n41134,
    n41132, n41133, n41135, n42341, n41163, n41161, n41160, n41162, n41164,
    n41184, n41175, n41174, n41180, n41177, n41179, n41181, n41188, n41193,
    n41189, n41190, n41192, n41202, n41277, n41195, n41198, n41197, n41199,
    n41205, n41207, n41228, n41210, n41220, n41218, n41216, n41215, n41217,
    n41219, n41226, n41247, n41241, n41251, n41261, n41262, n41267, n41266,
    n41274, n41270, n41273, n41282, n41288, n41285, n41292, n41291, n41293,
    n41300, n41297, n41304, n41303, n41305, n41315, n41313, n41312, n41323,
    n41321, n41320, n41322, n41379, n41328, n41353, n41334, n41343, n41346,
    n41347, n41360, n41361, n41364, n41366, n41367, n41377, n41376, n41383,
    n41385, n41396, n41392, n41405, n41419, n41406, n41412, n41409, n41517,
    n41523, n41420, n41428, n41427, n41432, n41430, n41429, n41431, n41433,
    n41440, n41446, n41445, n41449, n41447, n41448, n41460, n41452, n41464,
    n41463, n41468, n41466, n41465, n41467, n41469, n41930, n41480, n41478,
    n41476, n41475, n41477, n41479, n43847, n41487, n41485, n41483, n41482,
    n41484, n41486, n41489, n41700, n41494, n41497, n41498, n41500, n41503,
    n41501, n41704, n41502, n41507, n41505, n41506, n41508, n41522, n41521,
    n41524, n41525, n41533, n41551, n41550, n41544, n41570, n41617, n41572,
    n41571, n41576, n41574, n41573, n41575, n41582, n41577, n41580, n41579,
    n41581, n41586, n41584, n41583, n41585, n41610, n41587, n41590, n41589,
    n41596, n41594, n41593, n41595, n41608, n41600, n41599, n41606, n41604,
    n41603, n41605, n41607, n41609, n41787, n41612, n41616, n41618, n41621,
    n41620, n41630, n41623, n41622, n41627, n41625, n41624, n41626, n41628,
    n41629, n41636, n41634, n41632, n41633, n41635, n41655, n41638, n41637,
    n41647, n41640, n41639, n41644, n41642, n41641, n41643, n41645, n41646,
    n41653, n41651, n41649, n41650, n41652, n41654, n41782, n41786, n41658,
    n41663, n41661, n41660, n41662, n41665, n41664, n41666, n41674, n41673,
    n41676, n41686, n41690, n41689, n41694, n41692, n41691, n41693, n41695,
    n41717, n41715, n41701, n41706, n41705, n41709, n41708, n41710, n41720,
    n41721, n41739, n41723, n41722, n41729, n41738, n41740, n41741, n41751,
    n41753, n41752, n41767, n41761, n41760, n41762, n41766, n41768, n41775,
    n41774, n41779, n41777, n41776, n41778, n41780, n41788, n41792, n41791,
    n42755, n41794, n41793, n41803, n41796, n41795, n41800, n41798, n41797,
    n41799, n41801, n41802, n41809, n41807, n41806, n41808, n41828, n41811,
    n41810, n41820, n41813, n41812, n41817, n41815, n41814, n41816, n41818,
    n41819, n41826, n41824, n41823, n41825, n41827, n42753, n41829, n41830,
    n41835, n41833, n41832, n41834, n41837, n41836, n41838, n41843, n41847,
    n41861, n41897, n41849, n41853, n41851, n41850, n41852, n41868, n41870,
    n41892, n41887, n41871, n41885, n41878, n41883, n41881, n41880, n41882,
    n41884, n41890, n41895, n41911, n41909, n41903, n41901, n41900, n41915,
    n41914, n41917, n41918, n41925, n41923, n41922, n41924, n41948, n41929,
    n43756, n41937, n41950, n41961, n41970, n41954, n41957, n41956, n42582,
    n41967, n42967, n41964, n41966, n41975, n41971, n42825, n43337, n41978,
    n43350, n41982, n41980, n41981, n41983, n41984, n41985, n41987, n42544,
    n42921, n41986, n42010, n41993, n41991, n41992, n41994, n41997, n41996,
    n41998, n42000, n42001, n42548, n42005, n42014, n42031, n42030, n42035,
    n42033, n42032, n42034, n42036, n42039, n42038, n42045, n42044, n42049,
    n42047, n42046, n42048, n42050, n42053, n42060, n42080, n42078, n42065,
    n42067, n42068, n42072, n42071, n42074, n42566, n42073, n42075, n42087,
    n42082, n42088, n42101, n42102, n42116, n42141, n42108, n42702, n42106,
    n42107, n42112, n43150, n42300, n42113, n42650, n42114, n42115, n42119,
    n42118, n42124, n42120, n42123, n42648, n42136, n42144, n42142, n42143,
    n42148, n42146, n42147, n42170, n42159, n42154, n42153, n42157, n42155,
    n42156, n42158, n42163, n42162, n42164, n42165, n42167, n42179, n42177,
    n42176, n42187, n42188, n42651, n42192, n42193, n42195, n42194, n42597,
    n42230, n42200, n42210, n42211, n42216, n42217, n42595, n42218, n42221,
    n42220, n42222, n42425, n42223, n42601, n42231, n42291, n42232, n42271,
    n42381, n42239, n42241, n42251, n42261, n42267, n42262, n42265, n42263,
    n42613, n42264, n42266, n42272, n42274, n42273, n42275, n42299, n42286,
    n42290, n42440, n42292, n42302, n42301, n42317, n42306, n42313, n42308,
    n42453, n42311, n42310, n42312, n42328, n42326, n42350, n42698, n42363,
    n42361, n42349, n42357, n42355, n42873, n42356, n42366, n42368, n42370,
    n42369, n42377, n42399, n42384, n42389, n42392, n42390, n42634, n42391,
    n42395, n42394, n42402, n42401, n42421, n42407, n42406, n42419, n42413,
    n42411, n42420, n42428, n42426, n42427, n42430, n42445, n42443, n42441,
    n42442, n42444, n42456, n42454, n42455, n42459, n42458, n42460, n42478,
    n42476, n42474, n42518, n42475, n42497, n42484, n42485, n43043, n42489,
    n42490, n42493, n42502, n42513, n42681, n42506, n42509, n42508, n42521,
    n42523, n42530, n42525, n42884, n42528, n42529, n42531, n42542, n43463,
    n42541, n42540, n42543, n42545, n42972, n43449, n42550, n42559, n42578,
    n42576, n42567, n42570, n42569, n42571, n42581, n42594, n42583, n42591,
    n42596, n42602, n42603, n42605, n42606, n42607, n42615, n42614, n42618,
    n42617, n42636, n42635, n42639, n42638, n42644, n42649, n42655, n42653,
    n42654, n42674, n42663, n42666, n42843, n42667, n42678, n42677, n42686,
    n42690, n42689, n42694, n42692, n42691, n42693, n42695, n43152, n42701,
    n42704, n43147, n42703, n42735, n42993, n42726, n42724, n42858, n42729,
    n42728, n42738, n42737, n42742, n42740, n42739, n42741, n42743, n42752,
    n42751, n43059, n42757, n42756, n42761, n42759, n42758, n42760, n42767,
    n42762, n42765, n42763, n42764, n42766, n42771, n42769, n42768, n42770,
    n42795, n42772, n42775, n42773, n42774, n42781, n42776, n42779, n42777,
    n42778, n42780, n42793, n42785, n42784, n42791, n42789, n42788, n42790,
    n42792, n42794, n43060, n42797, n42798, n43058, n42808, n42806, n42805,
    n42807, n42810, n42809, n42811, n42816, n42819, n42818, n42827, n42831,
    n42830, n42839, n42846, n42844, n42845, n42849, n42848, n42863, n42861,
    n42859, n42860, n42862, n42886, n43010, n42890, n42896, n42996, n42891,
    n42893, n42895, n42918, n42903, n42902, n43206, n42912, n42910, n42954,
    n42920, n42923, n43352, n42925, n42926, n42929, n42928, n42932, n42931,
    n42940, n42944, n42943, n42948, n42946, n42945, n42947, n42949, n42964,
    n42957, n42955, n42956, n42961, n43461, n42970, n43438, n42968, n42969,
    n42984, n42991, n42994, n43005, n43003, n43001, n43017, n43002, n43011,
    n43026, n43020, n43041, n43034, n43345, n43037, n43036, n43045, n43044,
    n43048, n43047, n43049, n43064, n43062, n43063, n43393, n43066, n43065,
    n43070, n43068, n43067, n43069, n43076, n43071, n43074, n43073, n43075,
    n43080, n43078, n43077, n43079, n43108, n43081, n43084, n43083, n43090,
    n43088, n43087, n43089, n43106, n43096, n43095, n43104, n43102, n43101,
    n43103, n43105, n43107, n43391, n43110, n43109, n43115, n43113, n43112,
    n43114, n43116, n43123, n43122, n43127, n43125, n43124, n43126, n43128,
    n43131, n43136, n43140, n43139, n43187, n43149, n43160, n43151, n43157,
    n43153, n43163, n43161, n43162, n43226, n43757, n43166, n43580, n43169,
    n43167, n43168, n43205, n43191, n43197, n43318, n43532, n43214, n43212,
    n43228, n43213, n43218, n43234, n43232, n43227, n43230, n43229, n43231,
    n43285, n43244, n43243, n43250, n43248, n43247, n43249, n43259, n43253,
    n43252, n43257, n43255, n43254, n43256, n43258, n43283, n43263, n43262,
    n43269, n43267, n43266, n43268, n43281, n43273, n43272, n43279, n43277,
    n43276, n43278, n43280, n43282, n43284, n43287, n43292, n43289, n43288,
    n43290, n43291, n43296, n43299, n43301, n43308, n43307, n43312, n43310,
    n43309, n43311, n43313, n43319, n43320, n43327, n43340, n43332, n43334,
    n43336, n43338, n43339, n43357, n43349, n43346, n43355, n43353, n43354,
    n43356, n43360, n43364, n43363, n43388, n43373, n43375, n43381, n43385,
    n43395, n43392, n43397, n43396, n43406, n43399, n43398, n43403, n43401,
    n43400, n43402, n43404, n43405, n43413, n43411, n43410, n43412, n43432,
    n43415, n43414, n43424, n43417, n43416, n43421, n43419, n43418, n43420,
    n43422, n43423, n43430, n43428, n43427, n43429, n43431, n43433, n43435,
    n43440, n43439, n43445, n43446, n43450, n43451, n43452, n43460, n43454,
    n43458, n43457, n43459, n43468, n43465, n43464, n43466, n43467, n43708,
    n43470, n43471, n43473, n43478, n43477, n43494, n43480, n43479, n43492,
    n43482, n43481, n43488, n43486, n43485, n43487, n43489, n43491, n43493,
    n43520, n43498, n43497, n43511, n43502, n43501, n43507, n43505, n43504,
    n43506, n43508, n43510, n43518, n43516, n43513, n43515, n43517, n43519,
    n43521, n43526, n43541, n43585, n43542, n43553, n43556, n43555, n43563,
    n43557, n43561, n43560, n43562, n43789, n43568, n43574, n43576, n43579,
    n43596, n43588, n43601, n43600, n43746, n43658, n43608, n43665, n43610,
    n43624, n43615, n43614, n43759, n43620, n43616, n43618, n43619, n43622,
    n43646, n43621, n43623, n43632, n43631, n43642, n43636, n43635, n43637,
    n43647, n43648, n43655, n43688, n43664, n43666, n43760, n43674, n43673,
    n43675, n43677, n43778, n43676, n43679, n43678, n43680, n43683, n43692,
    n43691, n43706, n43704, n43700, n43699, n43701, n43710, n43715, n43714,
    n43724, n43723, n43726, n43730, n43733, n43736, n43742, n43740, n43739,
    n43745, n43892, n43810, n43752, n43827, n43825, n43851, n43758, n43879,
    n43761, n43762, n43764, n43815, n43763, n43765, n43768, n43787, n43779,
    n43780, n43790, n43793, n43792, n43801, n43799, n43798, n43805, n43824,
    n43816, n43817, n43831, n43873, n43839, n43846, n43841, n43869, n43845,
    n43860, n43848, n43881, n43849, n43856, n43852, n43854, n43855, n43858,
    n43918, n43857, n43859, n43862, n43863, n43865, n43875, n43874, n43890,
    n43885, n43883, n43900, n43882, n43884, n43906, n43910, n43901, n43902,
    n43908, n43929, n43923, n43919, n43920, n43926, n43928, n43936, n43934,
    n43935, n43941, n43939, n43938, n43940, n43946, n43944, n43943, n43945,
    n43951, n43949, n43948, n43950, n43956, n43954, n43953, n43955, n43961,
    n43959, n43958, n43960, n43966, n43964, n43963, n43965, n43971, n43969,
    n43968, n43970, n43976, n43974, n43973, n43975, n43981, n43979, n43978,
    n43980, n43988, n43986, n43985, n43987, n43999, n43991, n43997, n43995,
    n43996, n43998, n44001, n44006, n44004, n44005, n44010, n44009, n44011,
    n44018, n44016, n44015, n44017, n44027, n44025, n44024, n44026, n44033,
    n44031, n44030, n44032, n44038, n44036, n44035, n44037, n44043, n44041,
    n44040, n44042, n44048, n44046, n44045, n44047, n44053, n44051, n44050,
    n44052, n44058, n44056, n44055, n44057, n44062, n44060, n44059, n44061,
    n44067, n44065, n44064, n44066, n44072, n44070, n44069, n44071, n44077,
    n44075, n44074, n44076, n44081, n44079, n44078, n44080, n44085, n44083,
    n44082, n44084, n44090, n44088, n44087, n44089, n44097, n44095, n44094,
    n44096, n44101, n44103, n44104, n44110, n44108, n44109;
  assign n43927 = ~n43923 | ~n43922;
  assign n43914 = ~n43846 | ~n43845;
  assign n33474 = ~n31820 & ~n31819;
  assign n43525 = ~n32150 & ~n32149;
  assign n32110 = ~n31717 | ~n31716;
  assign n43813 = n34909 & n39531;
  assign n42971 = ~n42548 & ~n42547;
  assign n41949 = ~n42501 | ~P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n42242 = ~n26503 | ~n26502;
  assign n36904 = ~n25966 | ~n25965;
  assign n27875 = ~n26499 & ~n28061;
  assign n39578 = ~n26527;
  assign n26498 = ~n27853 & ~n43835;
  assign n43462 = ~n22933;
  assign n27853 = n27860 ^ n27858;
  assign n34270 = ~n22916;
  assign n26432 = n26391 ^ n26390;
  assign n24787 = ~n34576 | ~n25932;
  assign n23673 = ~n40306 | ~n31816;
  assign n40080 = n24165;
  assign n40081 = ~n31382 | ~n31721;
  assign n39615 = n27247 | n27246;
  assign n25897 = ~n24715 | ~n24714;
  assign n24715 = ~n24623;
  assign n37965 = ~n26266 & ~n26253;
  assign n37279 = ~n23677 | ~n23683;
  assign n32334 = ~n24445 | ~n24444;
  assign n24337 = ~n24336 & ~n24335;
  assign n24434 = ~n35165 & ~n31936;
  assign n34552 = ~n24340 ^ n24339;
  assign n23607 = ~n23605 | ~n23604;
  assign n35392 = ~n33502 & ~n27058;
  assign n36320 = ~n27071 & ~n36049;
  assign n22903 = ~n36316;
  assign n32337 = ~n26044 & ~n31721;
  assign n22914 = n36295;
  assign n22919 = n36306;
  assign n36317 = ~n27095;
  assign n37289 = ~n23084 & ~n23083;
  assign n31721 = ~n34187;
  assign n43061 = ~n23053 & ~n23052;
  assign n23523 = ~n23724 | ~n23322;
  assign n39892 = ~n32238;
  assign n23575 = ~n36795;
  assign n36795 = ~n23489 & ~n23488;
  assign n22947 = n23818 & n23817;
  assign n25634 = ~n23464;
  assign n23481 = ~n23045 & ~n26878;
  assign n22911 = ~n43098;
  assign n23463 = ~n43098 & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n28587 = ~n32119 | ~n33727;
  assign n32127 = ~n23772 & ~n24795;
  assign n43408 = ~n35755 | ~n35718;
  assign n35715 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n26853 = ~n22927 & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n33727 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n32119 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n22928 = P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n35755 = ~n26153 & ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n32506 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n26153 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n24706 = ~n24122 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n43098 = ~n35755 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n43100 = ~n35728 | ~n26153;
  assign n26838 = ~n26877 & ~n35715;
  assign n43514 = ~n23720 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n24610 = ~n24562 | ~n24561;
  assign n24500 = ~n24479 & ~n24478;
  assign n23649 = ~n26513 & ~n23648;
  assign n22923 = n36299;
  assign n22913 = n36289;
  assign n28507 = ~n42501;
  assign n26044 = ~n24216 | ~n24117;
  assign n43054 = ~n42752 | ~n42751;
  assign n33556 = ~n32798 | ~n28079;
  assign n31779 = ~n31524 | ~n31493;
  assign n34569 = n32334 ^ n34258;
  assign n41718 = ~n24767 | ~n24766;
  assign n23053 = ~n23036 | ~n23035;
  assign n43750 = ~n43667 & ~n43666;
  assign n39522 = ~P2_STATE2_REG_3__SCAN_IN;
  assign n41894 = ~n43033 | ~n26052;
  assign n42175 = ~n41894 | ~n26064;
  assign n31718 = n32110 | n31721;
  assign n26579 = ~n26567 | ~n26566;
  assign n40693 = ~n43358 | ~n26588;
  assign n40350 = n28160 | n36363;
  assign n23415 = ~n22943 | ~n22931;
  assign n32149 = ~P2_STATE2_REG_0__SCAN_IN | ~n23539;
  assign n32798 = ~n32800 & ~n32799;
  assign n42708 = ~n42624 | ~n42522;
  assign n39531 = ~n28158 | ~n27892;
  assign n29436 = ~n28928 | ~n29308;
  assign n44019 = ~n43300 | ~n32238;
  assign n43694 = ~n43522 ^ n43521;
  assign n41264 = ~n41568 | ~n26912;
  assign n33548 = ~P2_STATE2_REG_0__SCAN_IN & ~n33545;
  assign n31662 = ~n31826 | ~n31534;
  assign n42336 = ~n41257;
  assign n43358 = ~n26585 | ~n34498;
  assign n33545 = n31822 & n31821;
  assign n43181 = ~n42993;
  assign n43823 = ~n43822 | ~n43821;
  assign n42939 = ~n42938 & ~n42937;
  assign n43554 = ~n43548 & ~n43547;
  assign n43370 = ~n43366 & ~n43365;
  assign n42838 = ~n42837 & ~n42836;
  assign n43595 = ~n43594 & ~n43593;
  assign n43772 = ~n43771 & ~n43770;
  assign n42987 = ~n42986 & ~n42985;
  assign n42685 = ~n42684 & ~n42683;
  assign n43821 = ~n43820 & ~n43819;
  assign n42684 = ~n42679 & ~n43341;
  assign n43771 = ~n43812 & ~n43755;
  assign n42986 = ~n43359 & ~n43341;
  assign n42837 = ~n42832 & ~n43341;
  assign n43594 = ~n43590 | ~n43589;
  assign n43366 = ~n43359 & ~n43358;
  assign n43548 = ~n43545 | ~n43544;
  assign n43656 = ~n43653 & ~n43652;
  assign n42593 = ~n42592 & ~n42591;
  assign n43786 = ~n43785 & ~n43784;
  assign n42938 = ~n42933 & ~n43341;
  assign n42496 = ~n42495 & ~n42494;
  assign n28563 = ~n28557 | ~n28556;
  assign n43652 = ~n43651 | ~n43650;
  assign n43053 = ~n43050 & ~n43049;
  assign n43545 = ~n43581 | ~n43913;
  assign n43629 = ~n43628 | ~n43627;
  assign n43590 = ~n43581 | ~n43876;
  assign n43784 = ~n43783 | ~n43782;
  assign n43687 = ~n43686 & ~n43685;
  assign n42555 = ~n42554 & ~n42553;
  assign n43145 = ~n43142 & ~n43141;
  assign n43030 = ~n43028 & ~n43027;
  assign n28734 = n28733 & n28732;
  assign n43686 = n43776 & n43876;
  assign n43628 = ~n43644 | ~n43876;
  assign n42376 = ~n42375 & ~n42374;
  assign n42504 = ~n42503 & ~n42502;
  assign n28556 = ~n28555 & ~n28554;
  assign n42495 = ~n43042 & ~n43341;
  assign n42590 = ~n42585 & ~n43341;
  assign n42554 = ~n43135 & ~n43341;
  assign n43221 = ~n43219 & ~n43218;
  assign n43822 = ~n43810 | ~n43809;
  assign n43025 = ~n43024 & ~n43023;
  assign n43219 = ~n43216 | ~n43215;
  assign n43237 = ~n43236 | ~n43235;
  assign n42824 = ~n42821 & ~n42820;
  assign n43538 = ~n43535 | ~n43534;
  assign n43773 = ~n43810 | ~n43748;
  assign n42976 = ~n42974 | ~n42973;
  assign n42503 = ~n42499 & ~n42498;
  assign n28856 = ~n28851 | ~n28850;
  assign n28555 = ~n28549 & ~n43341;
  assign n41974 = ~n41973 & ~n41972;
  assign n42009 = ~n42008 & ~n42007;
  assign n42375 = ~n42371 & ~n43341;
  assign n43534 = ~n43533 | ~n43549;
  assign n43630 = ~n43643 & ~n43893;
  assign n43008 = ~n43007 | ~n43006;
  assign n43535 = ~n43531 | ~n43530;
  assign n43236 = ~n43223 | ~n43876;
  assign n43328 = ~n43325 & ~n43324;
  assign n41973 = ~n41968 & ~n43341;
  assign n42499 = ~n28482 | ~n28481;
  assign n43023 = ~n43022 | ~n43021;
  assign n43894 = ~n43906 & ~n43893;
  assign n43907 = ~n43906 & ~n43924;
  assign n43436 = ~n43633 | ~n43523;
  assign n42008 = ~n42815 & ~n43341;
  assign n43204 = ~n43203 & ~n43202;
  assign n43653 = ~n43643 & ~n43924;
  assign n28851 = ~n28848 | ~n28847;
  assign n28855 = ~n28854 & ~n43027;
  assign n43747 = ~n43744 & ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n42535 = ~n42534 & ~n42533;
  assign n28482 = ~n28479 | ~n43462;
  assign n42481 = ~n42480 & ~n42479;
  assign n43324 = ~n43323 | ~n43322;
  assign n43531 = ~n43532 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n43609 = ~n43608 | ~n43660;
  assign n43533 = ~n43532;
  assign n42963 = ~n42962 & ~n42961;
  assign n42973 = ~n42972 | ~n22933;
  assign n43202 = ~n43201 | ~n43200;
  assign n43785 = ~n43775 & ~n43924;
  assign n43007 = ~n43014 | ~n43913;
  assign n42917 = ~n42916 & ~n42915;
  assign n43119 = ~n43130 | ~n43693;
  assign n41750 = ~n41749 | ~n41748;
  assign n43134 = ~n43130 | ~n43523;
  assign n42915 = ~n42914 | ~n42913;
  assign n43602 = ~n43598 | ~n43661;
  assign n42962 = ~n42959 | ~n42958;
  assign n43744 = ~n43746 & ~n43743;
  assign n42480 = ~n42515 & ~n43811;
  assign n28479 = ~n28478 | ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n28509 = ~n28506 & ~n28505;
  assign n42814 = ~n42885 | ~n43693;
  assign n43593 = ~n43592 & ~n43591;
  assign n42889 = ~n42885 | ~n43523;
  assign n43210 = ~n43208 | ~n43207;
  assign n42673 = ~n42672 & ~n42671;
  assign n41748 = ~n41747 & ~n41746;
  assign n43129 = ~n43143 | ~n32242;
  assign n42734 = ~n42733 & ~n42732;
  assign n28481 = ~n28507 | ~n28480;
  assign n43144 = ~n43143 | ~n43367;
  assign n43325 = ~n43315 & ~n43924;
  assign n43203 = ~n43315 & ~n43893;
  assign n41281 = ~n41280 & ~n41279;
  assign n42999 = ~n42995 | ~n42994;
  assign n42643 = ~n42631 | ~n42630;
  assign n42853 = ~n42840 & ~n43924;
  assign n42622 = ~n42610 | ~n42609;
  assign n43143 = ~n43120;
  assign n42472 = ~n42471 | ~n42470;
  assign n42732 = ~n42731 | ~n42730;
  assign n41747 = ~n41742 & ~n43341;
  assign n43208 = ~n43206;
  assign n43304 = ~n43368 | ~n43297;
  assign n42883 = ~n42882 | ~n42881;
  assign n42995 = ~n42991 | ~n42990;
  assign n41280 = ~n41275 & ~n43341;
  assign n28829 = ~n43120 & ~n44019;
  assign n42866 = ~n42865 | ~n42864;
  assign n42867 = ~n42854 & ~n43924;
  assign n43369 = ~n43368 | ~n43367;
  assign n43314 = ~n43368 | ~n32242;
  assign n42229 = ~n42228 & ~n42227;
  assign n42610 = ~n42623 | ~n42603;
  assign n43220 = ~n43222 | ~n43809;
  assign n42362 = ~n42361 & ~n42360;
  assign n42577 = n42576 & n42575;
  assign n41275 = ~n41193 | ~n41192;
  assign n43368 = ~n43571;
  assign n42631 = ~n42623 | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n42744 = ~n42822 | ~n32242;
  assign n42881 = ~n42880 & ~n42879;
  assign n42316 = ~n42315 & ~n42314;
  assign n42298 = ~n42297 & ~n42296;
  assign n42823 = ~n42822 | ~n43367;
  assign n42471 = ~n42468 | ~n42713;
  assign n42951 = ~n42898 | ~n43550;
  assign n43238 = n43222 & n43748;
  assign n43591 = ~n43551 & ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n42609 = ~n42608 | ~n42607;
  assign n42468 = ~n42469 | ~n42466;
  assign n42463 = ~n42450 & ~n43924;
  assign n42898 = ~n42897 | ~n42906;
  assign n43170 = ~n43550;
  assign n43052 = ~n43051 | ~n43367;
  assign n42879 = ~n42878 | ~n42877;
  assign n43009 = ~n43013 & ~n43924;
  assign n42575 = ~n42574 & ~n42573;
  assign n42434 = ~n42433 | ~n42432;
  assign n41716 = ~n41715 & ~n41714;
  assign n42449 = ~n42436 & ~n43924;
  assign n42360 = ~n42359 | ~n42358;
  assign n42661 = ~n42659 | ~n42658;
  assign n42448 = ~n42447 | ~n42446;
  assign n42623 = ~n42599 & ~n42598;
  assign n42950 = ~n43051 | ~n32242;
  assign n42470 = ~n42469 | ~n42717;
  assign n42296 = ~n42295 | ~n42294;
  assign n42710 = ~n42706 | ~n42992;
  assign n42630 = ~n42629 | ~n42628;
  assign n42435 = ~n42422 & ~n43924;
  assign n42227 = ~n42226 | ~n42225;
  assign n42169 = ~n42168 & ~n42167;
  assign n42450 = ~n42304 | ~n42656;
  assign n42599 = ~n42604 & ~n43893;
  assign n42380 = ~n42379 | ~n43809;
  assign n42422 = ~n42196 | ~n42378;
  assign n42079 = ~n42078 & ~n42077;
  assign n42659 = ~n42657 | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n42436 = ~n42277 | ~n42343;
  assign n42706 = ~n42705 | ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n42469 = ~n42465 | ~n42464;
  assign n42234 = ~n42604 & ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n42037 = ~n42028 | ~n32242;
  assign n41841 = ~n41842 | ~n43693;
  assign n42574 = ~n42563 & ~n42562;
  assign n42482 = ~n42514 | ~n43809;
  assign n42629 = ~n42627 | ~n42626;
  assign n28865 = ~n28864 | ~n28863;
  assign n28842 = ~n28841 | ~n28840;
  assign n43051 = ~n42941;
  assign n43040 = ~n43039 & ~n43038;
  assign n41714 = ~n41713 | ~n41712;
  assign n42869 = ~n42344 | ~n42708;
  assign n42152 = ~n42138 | ~n43809;
  assign n41510 = ~n41509 & ~n41508;
  assign n42127 = ~n42126 & ~n42125;
  assign n42627 = ~n42625 | ~n42652;
  assign n42418 = ~n42417 | ~n42416;
  assign n42196 = ~n42660 | ~n42215;
  assign n40807 = ~n40806 & ~n40805;
  assign n42573 = ~n42572 | ~n42571;
  assign n28503 = ~n28502 | ~n28501;
  assign n42604 = ~n42378 & ~n42628;
  assign n28840 = ~n28839 & ~n28838;
  assign n42277 = ~n42276 | ~n42282;
  assign n42304 = ~n42561 | ~n42303;
  assign n41712 = ~n41711 & ~n41710;
  assign n42151 = ~n42150 & ~n42149;
  assign n42344 = ~n42343 | ~n42350;
  assign n42647 = ~n42687 | ~n43297;
  assign n42077 = ~n42076 | ~n42075;
  assign n28864 = ~n42687 | ~n43367;
  assign n28475 = ~n43031 & ~n44019;
  assign n42852 = ~n42851 | ~n42850;
  assign n42213 = ~n42208 | ~n42207;
  assign n42150 = ~n42139 & ~n43811;
  assign n27935 = ~n27874 & ~n28074;
  assign n42343 = ~n42624 | ~n42524;
  assign n28085 = ~n28075 & ~n28074;
  assign n42562 = ~n42059 & ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n41509 = ~n41702 & ~n43811;
  assign n42671 = ~n42670 | ~n42669;
  assign n28502 = ~n41687 | ~n43367;
  assign n41891 = ~n41890 & ~n41889;
  assign n28742 = ~n28741 | ~n28740;
  assign n42687 = ~n28858;
  assign n26576 = ~n26575 | ~n26574;
  assign n28537 = ~n28536 | ~n28535;
  assign n41656 = ~n41619 | ~n41618;
  assign n42416 = ~n42415 & ~n42414;
  assign n42660 = ~n42624 | ~n42214;
  assign n41860 = ~n41859 & ~n41858;
  assign n41947 = ~n41946 & ~n41945;
  assign n41765 = ~n41755 & ~n41754;
  assign n42656 = ~n42624 | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n41615 = ~n41755 & ~n33538;
  assign n39567 = ~n39566 & ~n39565;
  assign n43922 = ~n43921 & ~n43920;
  assign n43528 = ~n43527 | ~n43526;
  assign n41687 = ~n42409;
  assign n28535 = ~n28534 & ~n28533;
  assign n41511 = ~n41489 | ~n41700;
  assign n42190 = n42189 & n42188;
  assign n28741 = ~n42042 | ~n43367;
  assign n42041 = ~n42042 | ~n43297;
  assign n41089 = ~n41088 & ~n41087;
  assign n43889 = ~n43888 & ~n43887;
  assign n42642 = ~n42641 & ~n42640;
  assign n26574 = ~n26573 & ~n26572;
  assign n42398 = ~n42397 & ~n42396;
  assign n41945 = ~n41944 | ~n41943;
  assign n41858 = ~n41857 | ~n41856;
  assign n43904 = ~n43903 & ~n43902;
  assign n42207 = ~n42206 | ~n42658;
  assign n43770 = ~n43769 | ~n43768;
  assign n42208 = ~n42205 | ~n42662;
  assign n41713 = ~n41701 | ~n41700;
  assign n43921 = ~n43916 & ~n43915;
  assign n41856 = ~n41855 & ~n41854;
  assign n39649 = ~n39648 & ~n39647;
  assign n42462 = ~n42461 | ~n42460;
  assign n41263 = ~n41258 | ~n41257;
  assign n43887 = ~n43899 & ~n43886;
  assign n40103 = ~n40102 & ~n40101;
  assign n25990 = ~n25989 | ~n25988;
  assign n42189 = n42183 & n42182;
  assign n42621 = ~n42620 & ~n42619;
  assign n42042 = ~n28735;
  assign n43639 = ~n43638 & ~n43637;
  assign n41499 = ~n41494 | ~n41493;
  assign n26560 = ~n40769 | ~n26559;
  assign n43903 = ~n43899 & ~n43915;
  assign n43769 = ~n43766 & ~n43765;
  assign n42397 = ~n42632 & ~n43811;
  assign n39565 = ~n39564 | ~n39563;
  assign n28084 = ~n28083 | ~n28082;
  assign n28835 = ~n28463 & ~n28462;
  assign n28518 = ~n28517 | ~n28516;
  assign n27821 = ~n27818 & ~n42336;
  assign n28074 = ~n41699 & ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n42069 = ~n42065 | ~n42064;
  assign n43861 = ~n43916 & ~n43886;
  assign n42409 = ~n28046 | ~n28045;
  assign n42205 = ~n42664 | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n42103 = ~n42098 | ~n42097;
  assign n26912 = ~n26911 | ~n26910;
  assign n40954 = ~n40953 & ~n40952;
  assign n27934 = ~n27933 | ~n27932;
  assign n40782 = ~n40781 & ~n40780;
  assign n41889 = ~n43916 & ~n41888;
  assign n42512 = ~n42511 & ~n42510;
  assign n41944 = ~n41939 & ~n41938;
  assign n42314 = ~n42313 | ~n42312;
  assign n42270 = ~n42269 & ~n42268;
  assign n41087 = ~n41086 | ~n41085;
  assign n41183 = ~n41182 | ~n41181;
  assign n28373 = ~n28372 | ~n28371;
  assign n27818 = ~n27756 & ~n27755;
  assign n39564 = n39562 & n39561;
  assign n25988 = ~n25987 & ~n25986;
  assign n43133 = ~n43132 | ~n43131;
  assign n41910 = n41909 & n41908;
  assign n41699 = n41488 & P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n28517 = ~n41772 | ~n43367;
  assign n43638 = ~n43756 & ~n43695;
  assign n41227 = ~n41226 & ~n41225;
  assign n43916 = ~n39582 ^ n39581;
  assign n41493 = ~n41492 | ~n41491;
  assign n40101 = ~n40100 | ~n40099;
  assign n43703 = ~n43702 & ~n43701;
  assign n43819 = ~n43818 | ~n43817;
  assign n43899 = ~n43524;
  assign n43782 = ~n43781 & ~n43780;
  assign n42269 = ~n42611 & ~n43811;
  assign n38813 = ~n38806 & ~n38805;
  assign n43627 = ~n43626 & ~n43625;
  assign n43888 = ~n43885 | ~n43884;
  assign n41258 = ~n41256 | ~n41255;
  assign n28463 = ~n28525 | ~n28524;
  assign n27848 = ~n27847 | ~n27846;
  assign n42064 = ~n42063 | ~n42081;
  assign n26559 = ~n26558 & ~n26557;
  assign n28372 = ~n28225 & ~n28224;
  assign n41771 = ~n41772 | ~n43297;
  assign n40953 = ~n40942 & ~n43811;
  assign n39648 = ~n39645 | ~n39644;
  assign n42098 = ~n42095 | ~n42305;
  assign n42097 = ~n42096 | ~n42303;
  assign n42182 = ~n42181 & ~n42180;
  assign n43434 = ~n43814 & ~n35967;
  assign n41423 = ~n41422 | ~n41421;
  assign n41256 = ~n41249 | ~n41248;
  assign n41736 = ~n41735 | ~n41734;
  assign n43626 = ~n43624 | ~n43623;
  assign n42203 = ~n42307 | ~n42199;
  assign n41943 = ~n43814 | ~n41942;
  assign n43818 = ~n43814 | ~n43813;
  assign n43685 = ~n43684 | ~n43683;
  assign n41908 = n41907 & n41906;
  assign n38665 = ~n38664 & ~n38663;
  assign n42813 = ~n42812 & ~n42811;
  assign n28491 = ~n28490 | ~n28489;
  assign n39713 = ~n39673 & ~n39672;
  assign n42063 = ~n42062 | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n27846 = ~n27845 & ~n27844;
  assign n28772 = ~n28769 & ~n42336;
  assign n43702 = ~n43878 & ~n43695;
  assign n27755 = ~n27754 | ~n27753;
  assign n26908 = ~n41566 ^ n41564;
  assign n42388 = ~n42386 & ~n42385;
  assign n42281 = ~n42279 | ~n42278;
  assign n28525 = ~n28044 & ~n28043;
  assign n41960 = ~n41959 & ~n41958;
  assign n41567 = ~n41566 | ~n41565;
  assign n42505 = ~n27031 | ~n27030;
  assign n41492 = ~n41490 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n39930 = ~n39926 & ~n39925;
  assign n41735 = ~n41731 & ~n41730;
  assign n28490 = ~n41461 | ~n43367;
  assign n42386 = ~n42384 & ~n42383;
  assign n43684 = ~n43681 & ~n43680;
  assign n39669 = ~n39666 & ~n39665;
  assign n41169 = ~n41167 & ~n41166;
  assign n42342 = ~n42340 & ~n42339;
  assign n41422 = ~n41416 & ~n41415;
  assign n40939 = ~n40938 & ~n40937;
  assign n42812 = ~n43611 & ~n43695;
  assign n39560 = ~n38803 & ~n39588;
  assign n43200 = ~n43199 & ~n43198;
  assign n27753 = ~n27752 & ~n27751;
  assign n41906 = ~n41905 & ~n41904;
  assign n43118 = ~n43117 & ~n43116;
  assign n40766 = ~n41079 & ~n40761;
  assign n28106 = ~n28103 & ~n42336;
  assign n41443 = ~n41461 | ~n43297;
  assign n26707 = ~n26706 | ~n26705;
  assign n43650 = ~n43649 & ~n43648;
  assign n28769 = ~n28768 & ~n28767;
  assign n38664 = ~n38661 | ~n38660;
  assign n42888 = ~n42887 | ~n42886;
  assign n41248 = ~n41247 | ~n41246;
  assign n41459 = ~n41458 & ~n41457;
  assign n40879 = ~n40878 & ~n40877;
  assign n42340 = ~n42336 & ~n42335;
  assign n41166 = ~n41165 | ~n41164;
  assign n43199 = ~n43197 | ~n43318;
  assign n28767 = ~n28766 | ~n28765;
  assign n39925 = ~n39924 | ~n39923;
  assign n43322 = ~n43321 & ~n43320;
  assign n41416 = ~n41399 & ~n41531;
  assign n26705 = ~n26704 & ~n26703;
  assign n27887 = ~n42086 | ~n42083;
  assign n41953 = ~n26682 | ~n26681;
  assign n41037 = ~n41036 & ~n41035;
  assign n28103 = ~n28102 & ~n28101;
  assign n40765 = ~n40764 & ~n40763;
  assign n40153 = ~n42382 & ~n26504;
  assign n41079 = ~n40764 | ~n40762;
  assign n41201 = ~n41200 & ~n41199;
  assign n40097 = ~n40095 & ~n40094;
  assign n42093 = ~n42086 | ~n42244;
  assign n39590 = ~n39588 & ~n39587;
  assign n41840 = ~n41839 & ~n41838;
  assign n43117 = ~n43672 & ~n43695;
  assign n41246 = ~n41245 & ~n41244;
  assign n40955 = ~n40941 | ~n43809;
  assign n41845 = ~n41844 | ~n41843;
  assign n38803 = ~n38801 & ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n28101 = ~n41532 & ~n42318;
  assign n39769 = ~n39768 & ~n39767;
  assign n26719 = ~n26713 & ~n44019;
  assign n42335 = ~n42334 & ~n42333;
  assign n37567 = ~n37565 & ~n37564;
  assign n40123 = ~n40119 & ~n40118;
  assign n43589 = ~n43588 & ~n43587;
  assign n25490 = ~n38016 | ~n25489;
  assign n38135 = n38016 & n38015;
  assign n41035 = ~n41034 | ~n41033;
  assign n43544 = ~n43543 & ~n43542;
  assign n38381 = ~n38380 & ~n38379;
  assign n27029 = ~n28485 | ~n28484;
  assign n41457 = ~n41456 | ~n41455;
  assign n41839 = ~n43196 & ~n43695;
  assign n41165 = ~n41155 & ~n41154;
  assign n41244 = ~n41243 | ~n41242;
  assign n37448 = ~n37447 & ~n37446;
  assign n37128 = ~n37127 & ~n37126;
  assign n38801 = ~n38802;
  assign n41678 = ~n41677 | ~n41676;
  assign n28765 = ~n28764 & ~n28763;
  assign n43235 = ~n43234 & ~n43233;
  assign n40846 = ~n40844 & ~n40843;
  assign n41614 = ~n41613 & ~n41612;
  assign n27833 = ~n27832 | ~n27831;
  assign n41123 = ~n41112 & ~n41111;
  assign n39588 = ~n38802 & ~n39558;
  assign n41668 = ~n41667 & ~n41666;
  assign n28763 = ~n41091 & ~n42318;
  assign n40844 = ~n40842 & ~n42336;
  assign n43215 = ~n43214 & ~n43213;
  assign n38802 = ~n39586 | ~n38800;
  assign n40869 = ~n40863 & ~n41237;
  assign n43233 = ~n43232 | ~n43231;
  assign n41194 = ~n26140 | ~n26139;
  assign n41112 = ~n41091 & ~n41531;
  assign n41268 = ~n41267 & ~n41266;
  assign n40118 = ~n40117 | ~n40116;
  assign n41155 = ~n41531 & ~n42319;
  assign n41764 = ~n41763 | ~n41762;
  assign n41255 = ~n41254 | ~n41253;
  assign n40721 = ~n40720 & ~n40719;
  assign n41143 = ~n41142 & ~n41141;
  assign n26681 = ~n26680 | ~n26679;
  assign n41224 = ~n40936 & ~n28338;
  assign n42334 = ~n42319 & ~n42318;
  assign n41033 = ~n41032 & ~n41031;
  assign n39712 = ~n39708 & ~n39707;
  assign n39767 = ~n39766 | ~n39765;
  assign n37738 = ~n37734 & ~n37733;
  assign n39707 = ~n39706 | ~n39705;
  assign n26596 = ~n26595 | ~n26594;
  assign n41031 = ~n41030 | ~n41029;
  assign n41141 = ~n41140 | ~n41139;
  assign n37505 = ~n37504 & ~n37503;
  assign n43587 = ~n43586 | ~n43585;
  assign n42913 = ~n42912 & ~n42911;
  assign n37563 = ~n37561 & ~n37560;
  assign n27744 = ~n28098 | ~n41513;
  assign n40719 = ~n40718 | ~n40717;
  assign n43006 = n43005 & n43004;
  assign n36911 = ~n36910 & ~n36909;
  assign n40842 = ~n40841 & ~n40840;
  assign n41254 = ~n41237 & ~n42318;
  assign n41667 = ~n41657 & ~n43695;
  assign n42958 = ~n42957 & ~n42956;
  assign n40863 = ~n40858 | ~n40857;
  assign n41562 = ~n41561 & ~n41560;
  assign n37352 = ~n37122 | ~n37121;
  assign n37827 = ~n37443 | ~n38014;
  assign n41611 = ~n43224;
  assign n41763 = ~n43225 | ~n41756;
  assign n41561 = ~n42336 & ~n41559;
  assign n40840 = ~n40839 | ~n40838;
  assign n39185 = ~n39184 & ~n39183;
  assign n39161 = ~n39160 & ~n39159;
  assign n39198 = ~n39197 & ~n39196;
  assign n40858 = ~n40856 | ~n40855;
  assign n38267 = ~n38266 & ~n38265;
  assign n39143 = ~n39142 & ~n39141;
  assign n39169 = ~n39168 & ~n39167;
  assign n41237 = ~n40862 & ~n40861;
  assign n39177 = ~n39176 & ~n39175;
  assign n39151 = ~n39150 & ~n39149;
  assign n39136 = ~n39134 & ~n39133;
  assign n41152 = ~n41151 | ~n41150;
  assign n41139 = ~n41138 & ~n41137;
  assign n40717 = ~n40716 & ~n40715;
  assign n37473 = ~n37463 | ~n37462;
  assign n37733 = ~n37732 | ~n37731;
  assign n43004 = ~n43003 & ~n43002;
  assign n42730 = ~n42729 & ~n42728;
  assign n38997 = ~n38996 & ~n38995;
  assign n42864 = ~n42863 & ~n42862;
  assign n39026 = ~n39025 & ~n39024;
  assign n39013 = ~n39012 & ~n39011;
  assign n38990 = ~n38986 & ~n38985;
  assign n26139 = ~n26138 | ~n26137;
  assign n36909 = ~n36908 | ~n36907;
  assign n40700 = ~n40699 & ~n40698;
  assign n38640 = ~n38638 & ~n38637;
  assign n39005 = ~n39004 & ~n39003;
  assign n43021 = ~n43020 & ~n43019;
  assign n38967 = ~n38963 & ~n38962;
  assign n26712 = ~n26138 & ~n26137;
  assign n38395 = ~n38394 & ~n38393;
  assign n39011 = ~n39010 | ~n39009;
  assign n39133 = ~n39132 | ~n39131;
  assign n39614 = ~n39611 & ~n39610;
  assign n39238 = ~n39237 & ~n39236;
  assign n39024 = ~n39023 | ~n39022;
  assign n40839 = ~n40819 & ~n40818;
  assign n39291 = ~n39290 & ~n39289;
  assign n38252 = ~n38250 & ~n38249;
  assign n41559 = ~n41558 & ~n41557;
  assign n39183 = ~n39182 | ~n39181;
  assign n39196 = ~n39195 | ~n39194;
  assign n39258 = ~n39257 & ~n39256;
  assign n38928 = ~n38922 & ~n38921;
  assign n39249 = ~n39248 & ~n39247;
  assign n39159 = ~n39158 | ~n39157;
  assign n36131 = ~n36127 & ~n36126;
  assign n38962 = ~n38961 | ~n38960;
  assign n37732 = ~n37730 & ~n37729;
  assign n39003 = ~n39002 | ~n39001;
  assign n37278 = ~n37268 | ~n37267;
  assign n39141 = ~n39140 | ~n39139;
  assign n39167 = ~n39166 | ~n39165;
  assign n38985 = ~n38984 | ~n38983;
  assign n40862 = ~n40860 & ~n41250;
  assign n39175 = ~n39174 | ~n39173;
  assign n40755 = ~n40754 & ~n40753;
  assign n39149 = ~n39148 | ~n39147;
  assign n40791 = ~n40790 | ~n40789;
  assign n42533 = ~n42532 | ~n42531;
  assign n37557 = ~n36858 | ~n36857;
  assign n26082 = ~n26081 | ~n26080;
  assign n24761 = ~n24760 | ~n24759;
  assign n39209 = ~n39205 & ~n39204;
  assign n41137 = ~n41136 | ~n41135;
  assign n39762 = ~n39761 & ~n39760;
  assign n36099 = ~n36098 & ~n36097;
  assign n39266 = ~n39265 & ~n39264;
  assign n37009 = ~n37007 | ~n37006;
  assign n38244 = ~n38234 & ~n38233;
  assign n38995 = ~n38994 | ~n38993;
  assign n39935 = ~n40707 & ~n39934;
  assign n39276 = ~n39275 & ~n39274;
  assign n42477 = ~n42476 & ~n42475;
  assign n37472 = ~n37471 | ~n37470;
  assign n38752 = ~n38750 & ~n38749;
  assign n41557 = ~n41556 & ~n42318;
  assign n37845 = ~n37843 & ~n37842;
  assign n40819 = ~n42318 & ~n40816;
  assign n37932 = ~n37928 & ~n37927;
  assign n38760 = ~n38758 & ~n38757;
  assign n41238 = ~n28759;
  assign n37747 = ~n37745 & ~n37744;
  assign n26086 = ~n41130;
  assign n37877 = ~n37865 & ~n37864;
  assign n37254 = ~n37253 & ~n37252;
  assign n37234 = ~n37218 & ~n37217;
  assign n39610 = ~n39609 | ~n39608;
  assign n26939 = ~n26938 | ~n26937;
  assign n38303 = ~n38293 & ~n38292;
  assign n40065 = ~n40064 & ~n40063;
  assign n38206 = ~n38204 & ~n38203;
  assign n37893 = ~n37889 & ~n37888;
  assign n37787 = ~n37785 & ~n37784;
  assign n37804 = ~n37802 & ~n37801;
  assign n38315 = ~n38312 & ~n38311;
  assign n37007 = ~n37005 & ~n37004;
  assign n37885 = ~n37881 & ~n37880;
  assign n37633 = ~n37631 & ~n37630;
  assign n38003 = ~n38002 & ~n38001;
  assign n37901 = ~n37897 & ~n37896;
  assign n38243 = ~P2_INSTQUEUE_REG_2__0__SCAN_IN | ~n39020;
  assign n39289 = ~n39288 | ~n39287;
  assign n26501 = ~n26500 & ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n38812 = ~n38811 & ~n38810;
  assign n39236 = ~n39235 | ~n39234;
  assign n37972 = ~n37960 & ~n37959;
  assign n38780 = ~n38777 & ~n38776;
  assign n37987 = ~n37986 & ~n37985;
  assign n38233 = ~n38232 | ~n38231;
  assign n38901 = ~n38900 & ~n38899;
  assign n37120 = ~n36547 | ~n36546;
  assign n38249 = ~n38248 | ~n38247;
  assign n39256 = ~n39255 | ~n39254;
  assign n27743 = ~n41252;
  assign n38198 = ~n38196 & ~n38195;
  assign n38922 = ~n41531 & ~n40816;
  assign n39247 = ~n39246 | ~n39245;
  assign n39264 = ~n39263 | ~n39262;
  assign n39274 = ~n39273 | ~n39272;
  assign n38219 = ~n38216 & ~n38215;
  assign n40753 = ~n41531 & ~n41556;
  assign n37979 = ~n37978 & ~n37977;
  assign n38011 = ~n38010 & ~n38009;
  assign n42911 = ~n42910 | ~n42954;
  assign n37351 = ~n37349 & ~n37348;
  assign n38276 = ~n38274 & ~n38273;
  assign n40496 = ~n40495 & ~n40494;
  assign n28761 = ~n28759 | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n24759 = ~n24758 & ~n24757;
  assign n26092 = ~n25993 & ~n25992;
  assign n38768 = ~n38766 & ~n38765;
  assign n37814 = ~n37812 & ~n37811;
  assign n26080 = ~n26079 & ~n26078;
  assign n39204 = ~n39203 | ~n39202;
  assign n38251 = ~P2_INSTQUEUE_REG_2__1__SCAN_IN | ~n39020;
  assign n40853 = ~n40861 | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n42532 = ~n42521 & ~n42520;
  assign n40860 = ~n41252 & ~n40859;
  assign n39684 = ~n39683 & ~n39682;
  assign n37822 = ~n37820 & ~n37819;
  assign n37795 = ~n37793 & ~n37792;
  assign n38744 = ~n38742 & ~n38741;
  assign n37995 = ~n37994 & ~n37993;
  assign n38302 = ~P2_INSTQUEUE_REG_10__5__SCAN_IN | ~n39284;
  assign n38571 = ~n38570 & ~n38569;
  assign n38796 = ~n38795 & ~n38794;
  assign n38765 = ~n38764 | ~n38763;
  assign n36125 = ~n36123 & ~n36122;
  assign n38215 = ~n38214 | ~n38213;
  assign n38388 = ~n25067 & ~n25066;
  assign n39192 = ~n39130 | ~n39531;
  assign n38981 = ~n38980 & ~n38979;
  assign n38572 = ~n38568 & ~n38567;
  assign n37842 = ~n37841 | ~n37840;
  assign n38001 = ~n38000 | ~n37999;
  assign n38273 = ~n38272 | ~n38271;
  assign n37864 = ~n37863 | ~n37862;
  assign n43019 = ~n43018 | ~n43017;
  assign n37985 = ~n37984 | ~n37983;
  assign n38311 = ~n38310 | ~n38309;
  assign n38203 = ~n38202 | ~n38201;
  assign n39598 = ~n39597 & ~n39596;
  assign n38292 = ~n38291 | ~n38290;
  assign n38776 = ~n38775 | ~n38774;
  assign n37801 = ~n37800 | ~n37799;
  assign n37004 = ~n37003 | ~n37002;
  assign n37252 = ~n37251 | ~n37250;
  assign n36547 = ~n36203 & ~n36202;
  assign n27863 = ~n27862 | ~P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n37744 = ~n37743 | ~n37742;
  assign n26938 = ~n42909 | ~n41756;
  assign n37277 = ~n37276 | ~n37275;
  assign n38757 = ~n38756 | ~n38755;
  assign n38248 = ~n38246 & ~n38245;
  assign n37888 = ~n37887 | ~n37886;
  assign n39609 = ~n39605 & ~n39604;
  assign n37959 = ~n37958 | ~n37957;
  assign n37631 = ~n37619 | ~n37618;
  assign n25993 = ~n26085 | ~n26084;
  assign n37927 = ~n37926 | ~n37925;
  assign n38741 = ~n38740 | ~n38739;
  assign n37880 = ~n37879 | ~n37878;
  assign n38367 = ~n38366 & ~n38365;
  assign n37811 = ~n37810 | ~n37809;
  assign n38579 = ~n38578 & ~n38577;
  assign n38966 = ~n38965 & ~n38964;
  assign n38580 = ~n38576 & ~n38575;
  assign n38195 = ~n38194 | ~n38193;
  assign n37977 = ~n37976 | ~n37975;
  assign n38587 = ~n38586 & ~n38585;
  assign n42877 = ~n42876 & ~n42875;
  assign n42358 = ~n42357 & ~n42356;
  assign n39683 = n42723 & n41756;
  assign n38588 = ~n38584 & ~n38583;
  assign n37792 = ~n37791 | ~n37790;
  assign n38351 = ~n38350 & ~n38349;
  assign n38009 = ~n38008 | ~n38007;
  assign n40816 = ~n38908 | ~n38907;
  assign n38989 = ~n38988 & ~n38987;
  assign n38749 = ~n38748 | ~n38747;
  assign n38359 = ~n38358 & ~n38357;
  assign n38232 = ~n38230 & ~n38229;
  assign n38343 = ~n38342 & ~n38341;
  assign n37784 = ~n37783 | ~n37782;
  assign n37819 = ~n37818 | ~n37817;
  assign n37896 = ~n37895 | ~n37894;
  assign n26085 = ~n25850 & ~n25849;
  assign n38272 = ~n38270 & ~n38269;
  assign n37383 = ~n37371 & ~n37370;
  assign n37971 = ~n37970 & ~n37969;
  assign n37391 = ~n37387 & ~n37386;
  assign n36852 = ~n36854 | ~n36489;
  assign n38740 = ~n38738 & ~n38737;
  assign n40054 = ~n43016;
  assign n38310 = ~n38308 & ~n38307;
  assign n37530 = ~n37528 & ~n37527;
  assign n27862 = ~n40757;
  assign n37200 = ~n37199 & ~n37198;
  assign n38692 = ~n38691 & ~n38690;
  assign n37931 = ~n37930 & ~n37929;
  assign n37407 = ~n37405 & ~n37404;
  assign n37892 = ~n37891 & ~n37890;
  assign n37211 = ~n37210 & ~n37209;
  assign n37152 = ~n37151 & ~n37150;
  assign n37390 = ~n37389 & ~n37388;
  assign n39208 = ~n39207 & ~n39206;
  assign n42293 = ~n42290 & ~n42289;
  assign n36279 = ~n36277 & ~n36276;
  assign n40485 = ~n40483 & ~n40482;
  assign n37251 = ~n37245 & ~n37244;
  assign n37900 = ~n37899 & ~n37898;
  assign n37595 = ~n37591 & ~n37590;
  assign n37606 = ~n37603 & ~n37602;
  assign n38291 = ~n38289 & ~n38288;
  assign n37425 = ~n37422 & ~n37421;
  assign n38202 = ~n38200 & ~n38199;
  assign n38242 = ~n38241 | ~n39016;
  assign n38775 = ~n38772 & ~n38771;
  assign n39130 = ~n39129 | ~n39188;
  assign n38711 = ~n38710 & ~n38709;
  assign n38756 = ~n38754 & ~n38753;
  assign n37800 = ~n37798 & ~n37797;
  assign n37382 = ~n37381 & ~n37380;
  assign n37841 = ~n37838 & ~n37837;
  assign n37399 = ~n37395 & ~n37394;
  assign n40752 = ~n40751 | ~n40750;
  assign n38940 = ~n38937 & ~n38936;
  assign n38194 = ~n38192 & ~n38191;
  assign n38583 = ~n38582 | ~n38581;
  assign n37818 = ~n37816 & ~n37815;
  assign n37876 = ~n37875 & ~n37874;
  assign n38720 = ~n38719 & ~n38718;
  assign n38214 = ~n38211 & ~n38210;
  assign n37743 = ~n37741 & ~n37740;
  assign n37398 = ~n37397 & ~n37396;
  assign n37192 = ~n37191 & ~n37190;
  assign n37791 = ~n37789 & ~n37788;
  assign n38674 = ~n38673 & ~n38672;
  assign n37884 = ~n37883 & ~n37882;
  assign n38748 = ~n38746 & ~n38745;
  assign n37168 = ~n37167 & ~n37166;
  assign n37176 = ~n37175 & ~n37174;
  assign n38764 = ~n38762 & ~n38761;
  assign n37184 = ~n37183 & ~n37182;
  assign n38683 = ~n38682 & ~n38681;
  assign n37783 = ~n37781 & ~n37780;
  assign n38701 = ~n38700 & ~n38699;
  assign n37160 = ~n37159 & ~n37158;
  assign n37810 = ~n37807 & ~n37806;
  assign n38170 = ~n38166 & ~n38165;
  assign n37850 = ~n37848 & ~n37847;
  assign n43872 = ~n43871 | ~n43870;
  assign n41018 = ~n41016 & ~n41015;
  assign n37386 = ~n37385 | ~n37384;
  assign n37555 = ~n37553 & ~n37552;
  assign n37745 = ~n37836 & ~n37739;
  assign n40757 = n27867 ^ n42353;
  assign n43844 = ~n43843 & ~n43868;
  assign n38313 = ~n37956 | ~n39531;
  assign n42619 = ~n42618 | ~n42617;
  assign n25066 = ~n25065 & ~n25064;
  assign n38301 = ~n38300 | ~n39279;
  assign n39804 = ~n39802 & ~n39801;
  assign n35363 = ~n36090 | ~n35334;
  assign n27737 = ~n27739 & ~n42337;
  assign n37590 = ~n37589 | ~n40484;
  assign n43474 = ~n43444 & ~n43443;
  assign n40086 = ~n43802 | ~n44021;
  assign n40751 = ~n27739;
  assign n39439 = ~n39436 & ~n39435;
  assign n43804 = ~n43803 | ~n43802;
  assign n37521 = ~n37520 & ~n37519;
  assign n38241 = ~n38240 | ~n38239;
  assign n37370 = ~n37369 | ~n37368;
  assign n36399 = ~n36394 & ~n36393;
  assign n36854 = ~n36487 | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n39129 = ~n39128 | ~n39127;
  assign n37394 = ~n37393 | ~n37392;
  assign n28162 = ~n39701 | ~n39700;
  assign n40483 = ~n42336 & ~n40469;
  assign n42517 = ~n37466 & ~n37272;
  assign n37467 = ~n37466 & ~n37465;
  assign n38027 = ~n38026 & ~n38025;
  assign n38807 = ~n37216 & ~n37215;
  assign n43838 = ~n43840 & ~n43842;
  assign n43843 = ~n43842;
  assign n43871 = ~n43840;
  assign n42432 = ~n42431 & ~n42430;
  assign n37589 = ~n37588 & ~n37587;
  assign n38209 = ~n37873 & ~n37872;
  assign n43868 = ~n43870;
  assign n38770 = ~n37379 & ~n37378;
  assign n37861 = ~n37860 & ~n37859;
  assign n26483 = ~n36488 | ~n26476;
  assign n38165 = ~n38164 | ~n38163;
  assign n41015 = ~n42336 & ~n41014;
  assign n42985 = ~n42984 | ~n43361;
  assign n37956 = ~n37955 & ~n37954;
  assign n38306 = ~n37968 & ~n37967;
  assign n39802 = ~n42336 & ~n39799;
  assign n37835 = ~n37615 & ~n37614;
  assign n37836 = ~n37628 & ~n37627;
  assign n38300 = ~n38299 | ~n38298;
  assign n25797 = ~n25796 | ~n25795;
  assign n42225 = ~n42224 & ~n42223;
  assign n39283 = ~n38287 & ~n38286;
  assign n40541 = ~n40539 & ~n40538;
  assign n38228 = ~n38236 & ~n38224;
  assign n39120 = ~n39124 & ~n39116;
  assign n39435 = ~n39434 | ~n39433;
  assign n40469 = ~n40468 & ~n40467;
  assign n43802 = ~n43442;
  assign n38328 = ~n38325 & ~n38335;
  assign n43303 = ~n43302 & ~n43301;
  assign n26339 = ~n26336;
  assign n38190 = ~n38187 & ~n38186;
  assign n39612 = ~n38338 | ~n38337;
  assign n40538 = ~n42336 & ~n40537;
  assign n40002 = ~n39999 & ~n39998;
  assign n37272 = ~n37271 & ~n37270;
  assign n37001 = ~n36275 & ~n36274;
  assign n43302 = ~n43569 & ~n43298;
  assign n37873 = ~n37868 & ~n37867;
  assign n37379 = ~n37374 & ~n37373;
  assign n39991 = ~n39988 & ~n39987;
  assign n40467 = ~n40466 & ~n42318;
  assign n38236 = ~n38223 | ~n39508;
  assign n37860 = ~n37866 & ~n37868;
  assign n40013 = ~n40010 & ~n40009;
  assign n39980 = ~n39977 & ~n39976;
  assign n40435 = ~n40433 & ~n40432;
  assign n40051 = ~n40047 & ~n40046;
  assign n38287 = ~n38295 & ~n38283;
  assign n39969 = ~n39966 & ~n39965;
  assign n36090 = ~n35331 | ~n35330;
  assign n37423 = ~n37044 | ~n39531;
  assign n41014 = ~n41013 & ~n41012;
  assign n42287 = ~n36377 & ~n36376;
  assign n37955 = ~n37963 & ~n37961;
  assign n39799 = ~n39798 & ~n39797;
  assign n37215 = ~n37214 & ~n37213;
  assign n42850 = ~n42849 & ~n42848;
  assign n43573 = ~n43570 & ~n43569;
  assign n37968 = ~n37963 & ~n37962;
  assign n40024 = ~n40021 & ~n40020;
  assign n40035 = ~n40032 & ~n40031;
  assign n38337 = ~n38336 | ~n38335;
  assign n41886 = ~n41885 | ~n41884;
  assign n39124 = ~n39112 | ~n39508;
  assign n43870 = ~n43834 | ~n43891;
  assign n26338 = ~n26337;
  assign n39434 = ~n39424 & ~n39423;
  assign n39845 = ~n39843 & ~n39842;
  assign n37588 = ~n40466 & ~n41531;
  assign n38875 = ~n38873 & ~n38872;
  assign n37615 = ~n37621 & ~n37620;
  assign n39877 = ~n39875 & ~n39874;
  assign n39861 = ~n39859 & ~n39858;
  assign n38859 = ~n38857 & ~n38856;
  assign n38164 = ~n38153 & ~n38152;
  assign n39890 = ~n39887 & ~n39886;
  assign n38896 = ~n38893 & ~n38892;
  assign n38843 = ~n38841 & ~n38840;
  assign n38883 = ~n38881 & ~n38880;
  assign n39837 = ~n39835 & ~n39834;
  assign n38186 = ~n38185 | ~n38184;
  assign n39829 = ~n39827 & ~n39826;
  assign n38851 = ~n38849 & ~n38848;
  assign n37628 = ~n37622 & ~n37621;
  assign n39853 = ~n39851 & ~n39850;
  assign n39869 = ~n39867 & ~n39866;
  assign n38867 = ~n38865 & ~n38864;
  assign n43840 = ~n43834 & ~n43891;
  assign n38049 = ~n38046 & ~n38045;
  assign n35331 = ~n36088 & ~n35329;
  assign n37044 = ~n37043 & ~n37042;
  assign n38435 = ~n38433 & ~n38432;
  assign n38089 = ~n38087 & ~n38086;
  assign n38073 = ~n38071 & ~n38070;
  assign n38105 = ~n38103 & ~n38102;
  assign n38427 = ~n38425 & ~n38424;
  assign n38097 = ~n38095 & ~n38094;
  assign n38121 = ~n38119 & ~n38118;
  assign n40537 = ~n40536 & ~n40535;
  assign n38419 = ~n38417 & ~n38416;
  assign n38113 = ~n38111 & ~n38110;
  assign n40433 = ~n42336 & ~n40430;
  assign n38223 = ~n38222 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n26458 = ~n36485 & ~n43835;
  assign n38459 = ~n38457 & ~n38456;
  assign n37963 = ~n37949 | ~n39508;
  assign n39423 = ~n41011 & ~n41531;
  assign n39460 = ~n39458 & ~n39457;
  assign n43834 = ~n43833 | ~n43835;
  assign n39112 = ~n39111 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n28726 = ~n28725 | ~n28724;
  assign n43830 = ~n43829 & ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n37779 = ~n37770 & ~n37769;
  assign n38185 = ~n38177 & ~n38176;
  assign n43671 = ~n43751 | ~n43749;
  assign n38620 = ~n38619 & ~n38618;
  assign n40085 = ~n40079 | ~n40078;
  assign n38930 = ~n38631 & ~n38630;
  assign n41012 = ~n41011 & ~n42318;
  assign n37145 = ~n37144 | ~n38316;
  assign n37205 = ~n37138 & ~n37137;
  assign n37941 = ~n37645 | ~n39531;
  assign n40644 = ~n40642 & ~n40641;
  assign n38045 = ~n38044 | ~n40434;
  assign n42494 = ~n42493 | ~n42492;
  assign n42669 = ~n42668 & ~n42667;
  assign n38336 = ~n39524 & ~n38322;
  assign n38451 = ~n38449 & ~n38448;
  assign n37366 = ~n37373 | ~n37372;
  assign n38443 = ~n38441 & ~n38440;
  assign n38134 = ~n38131 & ~n38130;
  assign n39797 = ~n39796 & ~n42318;
  assign n38480 = ~n38477 & ~n38476;
  assign n37868 = ~n37856 | ~n39508;
  assign n38467 = ~n38465 & ~n38464;
  assign n38081 = ~n38079 & ~n38078;
  assign n38295 = ~n38282 | ~n39508;
  assign n37574 = ~n37573 | ~n38148;
  assign n43751 = ~n43669 | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n36376 = ~n36375 & ~n36374;
  assign n38282 = ~n38281 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n40536 = ~n42318 & ~n40532;
  assign n37043 = ~n37851 & ~n37038;
  assign n37608 = ~n37607 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n37037 = ~n37038 & ~n37034;
  assign n35329 = ~n35328 & ~P1_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n38222 = ~n39015 | ~n38221;
  assign n38618 = ~n38617 & ~n38625;
  assign n39111 = ~n39110 | ~n39187;
  assign n35816 = ~n36370 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n38631 = ~n38626 & ~n38625;
  assign n36118 = ~n36116 & ~n36115;
  assign n43663 = ~n43662 | ~n43661;
  assign n37138 = ~n37143 & ~n38316;
  assign n37144 = ~n37143;
  assign n40257 = ~n40256 | ~n40255;
  assign n37645 = ~n37644 & ~n37643;
  assign n41938 = ~n41937 | ~n41936;
  assign n39419 = ~n39417 & ~n39416;
  assign n42553 = ~n42552 | ~n43137;
  assign n40691 = ~n40688 & ~n40687;
  assign n39457 = ~n42336 & ~n39456;
  assign n43604 = ~n43603;
  assign n39530 = ~n39529 | ~n39528;
  assign n36274 = ~n36273 & ~n36272;
  assign n38322 = ~n38321 & ~n38320;
  assign n37769 = ~n37768 | ~n37767;
  assign n37949 = ~n37948 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n40430 = ~n40429 & ~n40428;
  assign n43836 = ~n41876 | ~n41875;
  assign n28828 = ~n28827 | ~n28826;
  assign n37856 = ~n37855 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n36568 = n37610 & n36574;
  assign n38177 = ~n41531 & ~n40532;
  assign n43826 = ~n43828 & ~n43825;
  assign n27859 = ~n27858;
  assign n36738 = ~n36737 | ~n39113;
  assign n38044 = ~n38043 & ~n38042;
  assign n36575 = ~n36574 | ~n36573;
  assign n40429 = ~n40408 & ~n42318;
  assign n41730 = ~n41729 | ~n41728;
  assign n36749 = ~n36745 & ~n39113;
  assign n39417 = ~n42336 & ~n39415;
  assign n37855 = ~n38208 | ~n37854;
  assign n43190 = ~n43189 & ~n43188;
  assign n38221 = ~n39021;
  assign n43603 = ~n43195 | ~n43194;
  assign n39456 = ~n39455 & ~n39454;
  assign n38320 = ~n39607 & ~n38319;
  assign n36737 = ~n36745;
  assign n37573 = ~n37571 | ~P3_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n38281 = ~n38280 | ~n39278;
  assign n38151 = ~n38150 | ~n38149;
  assign n42633 = ~n37125 | ~n37445;
  assign n40041 = ~n39955 | ~n39954;
  assign n37657 = ~n37652 & ~n37651;
  assign n43669 = ~n43670;
  assign n38933 = ~n38612;
  assign n43749 = ~n43670 | ~n43743;
  assign n28674 = ~n28673 | ~n28672;
  assign n36656 = ~n36655 & ~n36654;
  assign n40601 = ~n40599 & ~n40598;
  assign n39882 = ~n39818 | ~n39817;
  assign n37643 = ~n38220 & ~n37651;
  assign n39514 = ~n39527 & ~n39529;
  assign n42007 = ~n42006 | ~n42817;
  assign n42491 = ~n28723 & ~n28722;
  assign n39602 = ~n38319;
  assign n37948 = ~n38612 | ~n38305;
  assign n37028 = ~n37027 & ~n37026;
  assign n42333 = ~n42332 | ~n42331;
  assign n35321 = ~n35319 & ~n35318;
  assign n37365 = ~n38321 & ~n37364;
  assign n38888 = ~n39818 | ~n37493;
  assign n38043 = ~n41531 & ~n40408;
  assign n36574 = ~n36565 & ~n39524;
  assign n36370 = ~n36358 | ~n35780;
  assign n36088 = ~n35327 & ~n35366;
  assign n43662 = ~n43660 | ~n43659;
  assign n40078 = ~n40077 | ~n40076;
  assign n39110 = ~n39193;
  assign n27732 = ~n37766 | ~n37765;
  assign n37026 = ~n37025 | ~n37024;
  assign n41307 = ~n39543;
  assign n39377 = ~n39313 | ~n39312;
  assign n41221 = ~n41220 | ~n41219;
  assign n39415 = ~n39414 & ~n39413;
  assign n42665 = ~n35380 & ~n35379;
  assign n38616 = ~P2_STATEBS16_REG_SCAN_IN | ~n38615;
  assign n39527 = ~n39510 & ~n39509;
  assign n35780 = ~P2_STATE2_REG_1__SCAN_IN & ~n35806;
  assign n40622 = ~n40619 & ~n40618;
  assign n36206 = ~n35971 | ~n35970;
  assign n39817 = ~n39816 & ~n39815;
  assign n42332 = ~n42329 | ~P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n25115 = ~n36253;
  assign n41563 = ~n41554 | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n39955 = ~n39953 & ~n39952;
  assign n43670 = ~n43668 | ~n43835;
  assign n37493 = ~n38059 & ~n37492;
  assign n36654 = ~n36653 & ~n37944;
  assign n42980 = ~n42979 & ~n42978;
  assign n38305 = ~n36634 | ~n38279;
  assign n36565 = ~n38321 & ~n36577;
  assign n37033 = ~P2_STATEBS16_REG_SCAN_IN | ~n37045;
  assign n37571 = ~n38030 & ~n40431;
  assign n38126 = ~n38061 | ~n38060;
  assign n28768 = ~n28754 | ~n28753;
  assign n38149 = ~n38173 | ~n40531;
  assign n38174 = ~n38173 & ~n38172;
  assign n42057 = ~n42054 | ~P3_EBX_REG_31__SCAN_IN;
  assign n35327 = ~n35326 & ~n35325;
  assign n43189 = ~n43186 | ~n43185;
  assign n43180 = ~n43179 & ~n43178;
  assign n39455 = ~n39447 | ~n39446;
  assign n38472 = ~n38409 | ~n39954;
  assign n42137 = ~n42133 & ~n42132;
  assign n39101 = ~n39042 | ~n39041;
  assign n43376 = ~n28671 & ~n28721;
  assign n38959 = ~n38957 & ~n38956;
  assign n35326 = ~n35323 & ~n35322;
  assign n39543 = ~n39507 & ~n37947;
  assign n37492 = ~n38884 & ~n37491;
  assign n38497 = ~n38496 & ~n38495;
  assign n42937 = ~n42936 | ~n42935;
  assign n40666 = ~n40664 & ~n40663;
  assign n39042 = ~n39953 & ~n39040;
  assign n42329 = ~n42328 | ~n42327;
  assign n26383 = ~n26360 | ~n26359;
  assign n43179 = ~n43172 & ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n39187 = ~n36744 | ~n38279;
  assign n42056 = ~P3_EBX_REG_30__SCAN_IN | ~n42055;
  assign n37045 = ~n37946 & ~n37637;
  assign n42132 = ~n42131 & ~n42130;
  assign n41867 = ~n41866 | ~n42129;
  assign n42054 = ~n42131 | ~n42053;
  assign n38409 = ~n38407 & ~n38406;
  assign n39413 = ~n39412 | ~n39411;
  assign n43178 = ~n43177 | ~n43176;
  assign n28753 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN | ~n28752;
  assign n36736 = ~P2_STATEBS16_REG_SCAN_IN | ~n36744;
  assign n39313 = ~n39309 & ~n39308;
  assign n38061 = ~n38056 & ~n38055;
  assign n35806 = ~n35779 | ~n35778;
  assign n35832 = ~n24742 & ~n24741;
  assign n43194 = ~n43193 | ~n43599;
  assign n38030 = ~n37570 & ~n37572;
  assign n41933 = ~n41727 | ~n41726;
  assign n42027 = ~n42023 & ~n42022;
  assign n37147 = ~n37131 | ~n37130;
  assign n39015 = ~n37650 | ~n38279;
  assign n37854 = ~n36744 | ~n37947;
  assign n38150 = ~n38172 | ~P3_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n43186 = ~n43183 & ~n43182;
  assign n42646 = n42645 & n42644;
  assign n39952 = ~n39951 | ~n39950;
  assign n24721 = ~n24722;
  assign n24723 = ~n24722 & ~P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n24869 = ~n34812;
  assign n38173 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN & ~n38148;
  assign n43657 = ~n43607 | ~n43835;
  assign n37642 = ~P2_STATEBS16_REG_SCAN_IN | ~n37650;
  assign n39815 = ~n39814 | ~n39813;
  assign n28474 = ~n28473 | ~n28472;
  assign n38407 = ~n38411 & ~n38403;
  assign n26360 = ~n26352 & ~n26351;
  assign n43606 = ~n43192 | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n35323 = ~n34058 | ~n35324;
  assign n43185 = ~n43184 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n42117 = ~n34837 & ~n35378;
  assign n41685 = ~n41684 | ~n41863;
  assign n28671 = n28670 & n28669;
  assign n43188 = ~n43536 & ~n43187;
  assign n38056 = n38063 & n38064;
  assign n41553 = ~n41552 | ~P3_STATE2_REG_2__SCAN_IN;
  assign n42004 = ~n42003 & ~n43027;
  assign n41866 = ~n41864 | ~n41863;
  assign n36744 = ~n23700 & ~n34906;
  assign n39309 = ~n39306 & ~n39305;
  assign n42131 = ~n43930 | ~n42129;
  assign n37131 = ~n23700;
  assign n39951 = ~n39948 | ~n39947;
  assign n35778 = ~n35777 | ~n35776;
  assign n42133 = ~P3_EBX_REG_30__SCAN_IN & ~n42129;
  assign n42327 = ~n42326 & ~n42325;
  assign n42055 = ~P3_EBX_REG_31__SCAN_IN & ~n42129;
  assign n39040 = ~n39097 & ~n39039;
  assign n38495 = ~n38494 | ~n39041;
  assign n41534 = ~n41530 & ~n41529;
  assign n37491 = ~P1_STATE2_REG_3__SCAN_IN & ~n37490;
  assign n28752 = ~n28751 | ~n28750;
  assign n35602 = ~n35432 | ~n35431;
  assign n25978 = ~n40096 & ~n40094;
  assign n43348 = ~n43347 | ~n43346;
  assign n40880 = ~n40852 | ~n40851;
  assign n35517 = ~n33796 | ~n33795;
  assign n25973 = ~n39589 & ~n25972;
  assign n36109 = ~n34345 | ~n34814;
  assign n28102 = ~n28097 & ~n28096;
  assign n38172 = ~n38147 & ~n38146;
  assign n39814 = ~n39811 | ~n39810;
  assign n38148 = ~n37572 | ~n40431;
  assign n36652 = ~n23700 | ~n37130;
  assign n42022 = ~n42021 & ~n42020;
  assign n43177 = ~n43174 & ~n43173;
  assign n25965 = ~n24753 | ~n24752;
  assign n38066 = ~n38065 | ~n38064;
  assign n24741 = ~n24740 & ~P1_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n40349 = ~n40347 & ~n40346;
  assign n34521 = ~n34513 | ~n34512;
  assign n41122 = ~n41121 & ~n41120;
  assign n42309 = ~n33785 | ~n34836;
  assign n36793 = ~n36639 & ~n36638;
  assign n40852 = ~n40849 | ~n41153;
  assign n40096 = ~n25979 | ~n25977;
  assign n42129 = ~n41865 | ~P3_EBX_REG_29__SCAN_IN;
  assign n34063 = ~n33317 | ~n33794;
  assign n38412 = ~n38411 | ~n38410;
  assign n41249 = ~n41234 | ~n41259;
  assign n28097 = ~n28090 & ~n28089;
  assign n34813 = ~n24858 & ~n24857;
  assign n37490 = ~n37489 & ~n37488;
  assign n39589 = ~n38383 | ~n25971;
  assign n25976 = ~n25975 & ~n38385;
  assign n39810 = ~n39946 & ~n39809;
  assign n41529 = ~n41528 | ~n41527;
  assign n37572 = ~n37569 & ~n37568;
  assign n42020 = ~n42019 & ~n42018;
  assign n37859 = ~n37869 & ~n37858;
  assign n34585 = ~n34584;
  assign n39947 = ~n39946 & ~n39945;
  assign n43536 = ~n43171 | ~n43835;
  assign n23700 = ~n23699 ^ n25106;
  assign n24672 = ~n35330 & ~P1_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n42040 = n42039 & n42038;
  assign n40407 = ~n40405 & ~n40404;
  assign n28059 = ~n28058 | ~n28057;
  assign n38064 = ~n39946 & ~n38054;
  assign n40151 = ~n40149 & ~n40148;
  assign n38494 = ~n38493 | ~n38492;
  assign n24720 = ~n24717 | ~n26568;
  assign n43209 = ~n42905 | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n24742 = ~n24739 & ~n24738;
  assign n42568 = ~n33558 | ~n33557;
  assign n25963 = ~n24754 | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n39039 = ~P1_STATE2_REG_3__SCAN_IN & ~n39038;
  assign n35432 = ~n28228 & ~n28227;
  assign n28751 = ~n41245 & ~n28749;
  assign n42374 = ~n42373 | ~n42372;
  assign n42325 = ~n42324 | ~n42323;
  assign n42975 = ~n43448 & ~n42550;
  assign n42836 = ~n42835 | ~n42834;
  assign n28732 = ~n28731 | ~n28853;
  assign n41552 = ~n41551 | ~n42324;
  assign n34131 = ~n34129 & ~n34687;
  assign n42019 = ~n42017 | ~n42016;
  assign n40482 = ~n40481 & ~n40480;
  assign n25110 = ~n25107;
  assign n41995 = ~n43462 | ~n41994;
  assign n39809 = ~n39944 & ~n39808;
  assign n40404 = ~n40403 & ~n40402;
  assign n36152 = ~n36150 & ~n36149;
  assign n34094 = ~n34092 & ~n34687;
  assign n28228 = ~n34652 | ~n34651;
  assign n26402 = ~n26395 & ~n26394;
  assign n24739 = ~n24737 & ~n24736;
  assign n35627 = ~n34511 & ~n34510;
  assign n42021 = ~P3_STATE2_REG_0__SCAN_IN & ~n42015;
  assign n42331 = ~n42330 | ~n42337;
  assign n27756 = ~n41398 & ~n41235;
  assign n39945 = ~n39944 & ~n39943;
  assign n40976 = ~n40975 | ~n40974;
  assign n40345 = ~n40344 & ~n40343;
  assign n38054 = ~n39944 & ~n38053;
  assign n40582 = ~n40578 & ~n40577;
  assign n35324 = ~n34057 | ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n39304 = ~n39944 & ~n39303;
  assign n42324 = ~n41550 & ~n41549;
  assign n24754 = ~n43462 | ~n24751;
  assign n28853 = ~n43462 | ~n42828;
  assign n41865 = ~n41683 & ~n41682;
  assign n38493 = ~n38491 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n35155 = ~n34690 | ~n34689;
  assign n41067 = ~n41064 & ~n41063;
  assign n28096 = ~n28095 & ~n28094;
  assign n26369 = ~n26363 | ~n26362;
  assign n28749 = ~n28748 | ~n28747;
  assign n26379 = ~n26373 | ~n26372;
  assign n39038 = ~n39037 & ~n39036;
  assign n41013 = ~n41010 | ~n41009;
  assign n41424 = ~n41398 & ~n41397;
  assign n38410 = ~n39946 & ~n38402;
  assign n26422 = ~n26421 | ~n26420;
  assign n41234 = ~n42330 | ~P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n43173 = ~n42901 | ~n42900;
  assign n40539 = ~n40531 & ~n40530;
  assign n26423 = ~n26419 | ~n26418;
  assign n40094 = n43462 & n38643;
  assign n26580 = ~n26569 | ~n26568;
  assign n28090 = ~n28748;
  assign n26416 = ~n26415 | ~n26414;
  assign n37489 = ~n37487 & ~n39944;
  assign n26417 = ~n26413 | ~n26412;
  assign n26408 = ~n26407 | ~n26406;
  assign n42905 = ~n42907;
  assign n43207 = ~n42907 | ~n42906;
  assign n43530 = ~n43175 | ~n43835;
  assign n41530 = ~n41512 & ~n41513;
  assign n41121 = ~n41117 & ~n41512;
  assign n41528 = ~n41526 & ~n41525;
  assign n26401 = ~n26400 & ~n26399;
  assign n42907 = ~n42904 | ~n43835;
  assign n26395 = ~n26392 & ~n26790;
  assign n39303 = ~n39383 & ~n39374;
  assign n26409 = ~n26405 & ~n26806;
  assign n41549 = ~n41548 | ~n41547;
  assign n38053 = ~n38132 & ~n38123;
  assign n26418 = ~n38296 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n38835 = ~n38833 & ~n38832;
  assign n40754 = ~n41153 & ~n40749;
  assign n26419 = ~n37376 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n26406 = ~n39125 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n26403 = ~n37623 & ~n35254;
  assign n40520 = ~n40518 & ~n40517;
  assign n26400 = ~n26397 & ~n26396;
  assign n42017 = ~n42013 & ~n41671;
  assign n26413 = ~n39523 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n26414 = ~n37139 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n43182 = ~n42997 & ~n42902;
  assign n40402 = ~n40529 & ~n40401;
  assign n26415 = ~n36648 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n34511 = ~n34508 | ~n34507;
  assign n42408 = ~n28056 & ~n28523;
  assign n33733 = ~n34523 | ~n33732;
  assign n38491 = ~n38490 | ~n38489;
  assign n42589 = ~n42588 | ~n42587;
  assign n41009 = ~n41008 | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n34652 = ~n33918 & ~n33917;
  assign n41683 = ~n41393 | ~P3_EBX_REG_27__SCAN_IN;
  assign n42330 = ~n41555 & ~n41233;
  assign n36556 = ~n40325 & ~n37637;
  assign n41064 = ~n41062 & ~n41389;
  assign n35774 = ~n35771 | ~n35770;
  assign n39126 = ~n39125 | ~n39522;
  assign n26349 = ~n26348 & ~n26347;
  assign n42715 = ~n42714 & ~n42713;
  assign n26351 = ~n37623 & ~n43091;
  assign n26356 = ~n39523 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n28554 = ~n28553 | ~n28552;
  assign n26363 = ~n36648 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n26367 = ~n38296 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n26373 = ~n37376 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n39037 = ~n39035 & ~n39944;
  assign n39943 = ~n40037 & ~n40048;
  assign n41770 = n41769 & n41768;
  assign n26421 = ~n37870 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n40327 = ~n40324 & ~n40323;
  assign n38402 = ~n39944 & ~n38401;
  assign n41415 = ~n41414 | ~n41413;
  assign n40428 = ~n40427 & ~n40426;
  assign n41187 = ~n22933 & ~P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n40147 = ~n40146 & ~n40145;
  assign n39808 = ~n39888 & ~n39879;
  assign n40578 = ~n40572 | ~n40571;
  assign n26566 = ~n22933 | ~P1_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n28095 = ~n28092 | ~n28091;
  assign n40974 = ~n40973 | ~n40972;
  assign n40480 = ~n40529 & ~n40479;
  assign n28748 = ~n28744 & ~n28756;
  assign n37487 = ~n38894 & ~n38889;
  assign n27823 = ~n22933 | ~P1_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n41120 = ~n41119 & ~n41118;
  assign n40255 = ~n40254 | ~n40253;
  assign n40468 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN & ~n40534;
  assign n41558 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN & ~n41555;
  assign n28754 = ~n41236 | ~n28744;
  assign n40236 = ~n40234 & ~n40233;
  assign n41526 = ~n41516 & ~n41515;
  assign n40530 = ~n40529 & ~n40528;
  assign n40535 = ~n40534 & ~n40533;
  assign n42015 = ~n42014 & ~n42013;
  assign n34343 = ~n24850 | ~n24849;
  assign n41154 = ~n42337 & ~n41153;
  assign n41387 = ~n41381 | ~P3_STATE2_REG_1__SCAN_IN;
  assign n41512 = ~n41116 & ~n41115;
  assign n34269 = ~n34267 & ~n34687;
  assign n42714 = ~n42718 & ~n42712;
  assign n23664 = ~n23661;
  assign n26394 = ~n26393 & ~n43426;
  assign n40534 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN | ~n40465;
  assign n42997 = ~n42899 | ~n43835;
  assign n43807 = ~n43793 & ~n43792;
  assign n43472 = ~n43447 & ~n43446;
  assign n27350 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN | ~n41114;
  assign n26399 = ~n26398 & ~n26819;
  assign n40427 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN & ~n40465;
  assign n41393 = ~n41390 & ~n41389;
  assign n26348 = ~n26393 & ~n26345;
  assign n26347 = ~n26398 & ~n26346;
  assign n39798 = ~n39795 & ~n39794;
  assign n27040 = ~n27039 | ~n27038;
  assign n42683 = ~n42682 | ~n42681;
  assign n41555 = ~n41232 & ~n41231;
  assign n41153 = n40746 & n40745;
  assign n28744 = ~n41114 & ~n41235;
  assign n34507 = ~n34506 & ~n34505;
  assign n40572 = ~n40569 & ~n40568;
  assign n41413 = n41412 & n41411;
  assign n38401 = ~n38478 & ~n38469;
  assign n26250 = ~n37612 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n24618 = ~n24828 & ~n24745;
  assign n41548 = ~n41544 & ~n41543;
  assign n43444 = ~n43440 & ~n43439;
  assign n41168 = ~n41514 | ~n42337;
  assign n42900 = ~n42990 | ~n42992;
  assign n24840 = ~n24828 & ~n24873;
  assign n39035 = ~n39107 & ~n39102;
  assign n28891 = ~n28890 | ~n28889;
  assign n38296 = ~n26364;
  assign n24716 = ~n24710 | ~n24711;
  assign n37623 = ~n37612;
  assign n42719 = ~n42718 & ~n42717;
  assign n27720 = ~n37710;
  assign n40464 = ~n40462 & ~n40461;
  assign n26362 = ~n37965 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n38927 = ~n38926 & ~n38925;
  assign n39795 = ~n40240 & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n26412 = ~n37965 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n39794 = ~n39793 & ~n40524;
  assign n40232 = ~n40231 & ~n40230;
  assign n23661 = ~n23658 & ~n23657;
  assign n40526 = ~n40525 & ~n40524;
  assign n26292 = ~n37965;
  assign n42990 = ~n42721 | ~n43835;
  assign n42718 = ~n42711 & ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n43447 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN | ~n42965;
  assign n42586 = ~n41439 & ~n41438;
  assign n39454 = ~n40409 & ~P3_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n41006 = ~n40250 & ~n40249;
  assign n40400 = ~n40399 & ~n40398;
  assign n26239 = ~n38628 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n41972 = ~n41971 | ~n41970;
  assign n41236 = ~n41541 & ~n28755;
  assign n40465 = ~n40409 & ~n40421;
  assign n41411 = n41410 & n41409;
  assign n41114 = ~n41541 & ~n41516;
  assign n40478 = ~n40477 & ~n40476;
  assign n41232 = ~n41230 & ~n41229;
  assign n42464 = ~n42712 & ~n42711;
  assign n40516 = ~n40515 & ~n40514;
  assign n37638 = ~n32896 | ~n32895;
  assign n39424 = ~n41002 & ~n39420;
  assign n41229 = ~n41000 | ~n40999;
  assign n40249 = ~n40248 | ~n40247;
  assign n41378 = ~n41377 | ~n41376;
  assign n40818 = ~n41235 & ~n40817;
  assign n42965 = ~n42547 & ~n42537;
  assign n44020 = ~n32632 | ~n32631;
  assign n42712 = n42351 & n42350;
  assign n27751 = ~n41240 & ~n41407;
  assign n43437 = ~n42541 | ~n42540;
  assign n43791 = ~n43568 | ~n43567;
  assign n38925 = ~n41397 & ~n40817;
  assign n40409 = ~n39453 & ~n39452;
  assign n33731 = ~n34502 | ~n33728;
  assign n43012 = ~n42894 & ~n42893;
  assign n35769 = ~n35736 & ~n35735;
  assign n41458 = ~n41452 & ~n41451;
  assign n42717 = ~n42467 | ~n43835;
  assign n24615 = ~n24609 | ~n24611;
  assign n40524 = ~n39792 | ~n39791;
  assign n40475 = ~n40415 & ~n40414;
  assign n39792 = ~n40415 & ~n39789;
  assign n39420 = ~n37774 & ~n37772;
  assign n43567 = ~n43371 & ~n28886;
  assign n39452 = ~n39771 | ~n39774;
  assign n24623 = ~n24614 | ~n24613;
  assign n39442 = ~n39402 & ~n39401;
  assign n38176 = ~n38175 & ~n40533;
  assign n40964 = ~n40396 & ~n40395;
  assign n39414 = ~n39393 & ~n39392;
  assign n41969 = ~n26691 & ~n41437;
  assign n42280 = ~n42257 | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n40460 = ~n40459 & ~n40458;
  assign n42537 = ~P1_INSTADDRPOINTER_REG_26__SCAN_IN | ~n42930;
  assign n40999 = ~n39772 & ~n39771;
  assign n34502 = ~n33726 & ~n33725;
  assign n42466 = ~n42352 | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n28766 = ~n28756 | ~n41239;
  assign n40545 = ~n39743 | ~P3_EBX_REG_23__SCAN_IN;
  assign n42250 = ~n42387 & ~n42383;
  assign n37591 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN & ~n38175;
  assign n28557 = ~n28548 | ~P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n41746 = ~n41745 | ~n41744;
  assign n22916 = n34726;
  assign n41242 = ~n41241 & ~n41259;
  assign n40248 = ~n40246 & ~n40245;
  assign n24816 = ~n24815 | ~n24814;
  assign n24614 = ~n24575;
  assign n28756 = ~n41113 & ~n41240;
  assign n37021 = ~n36870 & ~n37713;
  assign n38790 = ~n37509 & ~n37229;
  assign n42527 = ~n42275 & ~n42700;
  assign n42383 = ~n42249 | ~n42248;
  assign n28869 = ~n28868 | ~n28867;
  assign n28838 = ~n28837 | ~n28836;
  assign n42538 = ~n42966 | ~n41984;
  assign n42346 = ~n42285 | ~n43835;
  assign n42278 = ~n42258 | ~n42601;
  assign n42254 = ~n42253 | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n43371 = ~n28877 & ~n43566;
  assign n43853 = ~n43617 | ~n43616;
  assign n41935 = ~n41214;
  assign n38175 = ~n38142 | ~n40470;
  assign n42892 = ~n42727 | ~n43152;
  assign n42558 = ~n41072 & ~n41073;
  assign n33725 = ~n33724 & ~n33723;
  assign n42592 = ~n42584 & ~n42583;
  assign n39743 = ~n39503 & ~n39502;
  assign n27750 = ~n41113 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n38188 = ~n38168 | ~n38167;
  assign n41902 = ~n41901 & ~n41900;
  assign n40770 = ~n26217 & ~n36846;
  assign n42930 = ~n42826 & ~n42921;
  assign n40414 = ~n40413 | ~n40412;
  assign n38047 = ~n37593 | ~n37592;
  assign n41451 = ~n35512 | ~n27841;
  assign n42178 = ~n42177 & ~n42176;
  assign n42652 = ~n42727;
  assign n41450 = ~n41019 & ~n29613;
  assign n38924 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~n40244;
  assign n40088 = ~n25957 | ~n39640;
  assign n42258 = ~n42256 | ~n43835;
  assign n42727 = ~n42122 | ~n42121;
  assign n24575 = ~n24502 | ~n24501;
  assign n24419 = ~n24418 & ~n24417;
  assign n37085 = ~n35841 & ~n35840;
  assign n28877 = ~n28876 & ~n28875;
  assign n40092 = ~n25961 & ~n25960;
  assign n37637 = ~n37945;
  assign n41942 = ~n41888;
  assign n33724 = ~n34489 & ~P1_STATE2_REG_1__SCAN_IN;
  assign n42966 = ~n41978 & ~n41977;
  assign n41214 = n28216 & n28215;
  assign n42249 = ~n42247 & ~n42246;
  assign n41239 = ~n41545 & ~n28755;
  assign n41373 = ~n41370 & ~n41369;
  assign n39557 = ~n36890 & ~n36889;
  assign n41019 = ~n26697 & ~n43566;
  assign n42171 = ~n41847 & ~n43566;
  assign n43617 = ~n43155 | ~n43154;
  assign n23697 = ~n23673 | ~n23672;
  assign n42584 = ~n41965 & ~n41964;
  assign n41073 = ~n40767 | ~n28064;
  assign n42676 = ~n41977 & ~n28547;
  assign n41124 = ~n40702 & ~n43566;
  assign n42121 = ~n43148 | ~n42702;
  assign n41888 = ~n23085 | ~n28370;
  assign n35361 = ~n34281 & ~n34280;
  assign n42122 = ~n43158 | ~n42120;
  assign n42248 = ~n42240 | ~n42215;
  assign n43559 = ~n42175;
  assign n28216 = ~n28211 | ~n41877;
  assign n38279 = ~n37947;
  assign n41934 = ~n39482;
  assign n41931 = ~n40602;
  assign n39640 = ~n38645 | ~n25953;
  assign n41369 = ~n41368 | ~n41367;
  assign n39785 = ~n39775 | ~n39395;
  assign n41859 = ~n41849 & ~P1_REIP_REG_21__SCAN_IN;
  assign n36542 = ~n36543;
  assign n34489 = ~n33720 | ~n33719;
  assign n41977 = ~n41271 | ~n28543;
  assign n42252 = ~n42243 | ~n43835;
  assign n42385 = ~n42240 & ~n42239;
  assign n41453 = ~n43794;
  assign n41946 = ~n41926 & ~n43808;
  assign n28886 = ~P1_REIP_REG_28__SCAN_IN & ~n28882;
  assign n36173 = ~n36170 & ~n36169;
  assign n43797 = ~n41129;
  assign n37713 = ~n36869 | ~n36868;
  assign n43386 = ~P1_REIP_REG_27__SCAN_IN & ~n43373;
  assign n41965 = ~n41271 | ~n41270;
  assign n36890 = ~n24154 & ~n24153;
  assign n39389 = ~n41542 | ~n40215;
  assign n43788 = ~n42488 & ~n28882;
  assign n40841 = ~n40815 & ~n41240;
  assign n40982 = ~n40960 & ~n40959;
  assign n41368 = ~n41358 | ~n41357;
  assign n42240 = ~n42209 | ~n43835;
  assign n43165 = ~n43159 | ~n42699;
  assign n39635 = ~n39634 & ~n39633;
  assign n34485 = ~n33713 & ~n33712;
  assign n40669 = ~n41869;
  assign n36895 = ~n41979;
  assign n40388 = ~n40969 & ~n40500;
  assign n28882 = ~n28874 | ~n43372;
  assign n41926 = ~n39732;
  assign n36866 = ~n39388 & ~n41397;
  assign n31796 = ~n24801 | ~n24800;
  assign n35172 = ~n34124 | ~n34119;
  assign n23693 = ~n24781 | ~n23692;
  assign n43767 = ~n43886;
  assign n35178 = ~n34124 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n36543 = ~n27891 & ~n23542;
  assign n37325 = ~n36403 | ~P3_EBX_REG_19__SCAN_IN;
  assign n43148 = ~n43159;
  assign n42246 = ~n42198 | ~n42197;
  assign n42400 = ~n41894;
  assign n43158 = ~n42699;
  assign n41271 = ~n28542 & ~n38650;
  assign n43748 = ~n43893;
  assign n43876 = ~n43755;
  assign n32145 = ~n32143;
  assign n27749 = ~n42321 & ~n38923;
  assign n28559 = ~n34279 & ~n43330;
  assign n27713 = n36193 & n27712;
  assign n24801 = ~n34560 | ~n25932;
  assign n41357 = ~n41356 | ~n41355;
  assign n38781 = ~n42185 & ~n37227;
  assign n40883 = ~n38687;
  assign n41283 = ~n39606;
  assign n26254 = ~n26253;
  assign n42198 = ~n42201 | ~n42100;
  assign n40436 = ~n34898;
  assign n23542 = ~n23541 | ~n23540;
  assign n41290 = ~n37808;
  assign n42662 = ~n42204 | ~n43835;
  assign n42539 = ~n42927 | ~n42922;
  assign n42236 = ~n42201 & ~n42200;
  assign n42092 = ~n42235;
  assign n36403 = ~n36177 & ~n36176;
  assign n41302 = ~n38696;
  assign n39934 = ~n32242;
  assign n38553 = ~n38486 | ~n38485;
  assign n38885 = ~n37478 | ~n37477;
  assign n41295 = ~n39201;
  assign n39098 = ~n39032 | ~n39031;
  assign n40894 = ~n38669;
  assign n40907 = ~n39233;
  assign n40906 = ~n38715;
  assign n39549 = ~n38706;
  assign n43372 = ~n42185 & ~n42160;
  assign n39732 = n41206 & n41204;
  assign n41921 = ~n36390;
  assign n41869 = ~n41204 & ~n41919;
  assign n41879 = ~n28196 | ~n37288;
  assign n39535 = ~n39244;
  assign n38650 = ~n32532 | ~n24157;
  assign n43716 = ~n43715 & ~n43714;
  assign n36459 = ~n35857 & ~n35856;
  assign n39240 = ~n39517;
  assign n38703 = ~n39542;
  assign n40500 = ~n36447 | ~n40441;
  assign n39883 = ~n39823 | ~n39822;
  assign n35962 = ~n35959 & ~n35958;
  assign n36167 = ~n36166 & ~n36165;
  assign n34124 = ~n34560;
  assign n39388 = ~n40221 | ~n36230;
  assign n40042 = ~n39961 | ~n39960;
  assign n40881 = ~n39156;
  assign n41318 = ~n38678;
  assign n43331 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN | ~n42924;
  assign n40277 = ~n40276 & ~n40275;
  assign n40186 = ~n40185 & ~n40184;
  assign n41358 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & ~n41339;
  assign n43341 = ~n36906;
  assign n41976 = ~n36891;
  assign n40205 = ~n40204 & ~n40203;
  assign n26550 = ~n26215;
  assign n41204 = ~n41718;
  assign n34287 = ~n42924;
  assign n32341 = ~n34071 & ~n32340;
  assign n39251 = ~n39541;
  assign n42927 = ~n36891 & ~n42924;
  assign n38687 = ~n36683 | ~n36682;
  assign n35959 = ~n35942 & ~n35941;
  assign n41370 = ~n41336 & ~n41335;
  assign n39200 = ~n41296;
  assign n39241 = ~n39516;
  assign n42185 = ~n42405;
  assign n39280 = ~n40899;
  assign n39230 = ~n40911;
  assign n43732 = ~n43734;
  assign n37808 = ~n36587 | ~n36586;
  assign n42802 = ~n43689;
  assign n41356 = ~n41352 | ~n41351;
  assign n43333 = n36891 & n28558;
  assign n23540 = ~n35719 | ~n35805;
  assign n25944 = ~n25984 | ~n25983;
  assign n39378 = ~n39318 | ~n39317;
  assign n33786 = ~n35381;
  assign n32144 = ~n23689 | ~n23688;
  assign n42235 = ~n42091 | ~n42090;
  assign n40242 = ~n39790 & ~n40998;
  assign n42244 = ~n42085 & ~n42084;
  assign n42201 = ~n42099 | ~n43835;
  assign n36177 = ~n35553 | ~P3_EBX_REG_17__SCAN_IN;
  assign n27706 = ~n27709 | ~P3_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n42091 = ~n42089 | ~n42088;
  assign n26057 = ~n34514 & ~n26056;
  assign n41339 = ~n41338 & ~n41337;
  assign n44021 = ~n43298;
  assign n39959 = ~n39030;
  assign n42305 = ~n42094 | ~n43835;
  assign n36955 = ~n36002;
  assign n41296 = ~n36688 & ~n36794;
  assign n39390 = ~n41546 | ~n40213;
  assign n35553 = ~n35421 & ~n35420;
  assign n41756 = ~n43695;
  assign n43693 = ~n41754;
  assign n38411 = ~n38400 & ~n39301;
  assign n42085 = ~n42089 & ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n26051 = ~n35465 | ~n44107;
  assign n24501 = ~n24500;
  assign n22946 = n35790 & n37279;
  assign n39790 = ~n39394 | ~n39775;
  assign n27709 = ~n27705 | ~n40127;
  assign n39036 = ~n39030 & ~n39942;
  assign n37302 = ~n35790;
  assign n34876 = ~n37279;
  assign n24612 = ~n24610;
  assign n35719 = ~n35766;
  assign n43362 = ~n43713;
  assign n40275 = ~n40274 & ~n40273;
  assign n41920 = ~n40350;
  assign n41352 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~n41340;
  assign n41336 = ~n41338;
  assign n39541 = ~n43061 & ~n36794;
  assign n36237 = ~n43937 & ~n35594;
  assign n40899 = ~n36795 & ~n36794;
  assign n42804 = ~n43697;
  assign n36794 = ~n36778;
  assign n43523 = ~n33538;
  assign n26206 = ~n26205 | ~n26204;
  assign n43911 = ~n43896;
  assign n40607 = ~n40652 | ~n40651;
  assign n43698 = ~n41759;
  assign n24766 = ~n41912;
  assign n43697 = ~n41759 | ~n25790;
  assign n25102 = ~n41759 | ~n25101;
  assign n42083 = ~n41496 & ~n27885;
  assign n39030 = ~n35870 | ~n36136;
  assign n35421 = ~n34404 | ~P3_EBX_REG_15__SCAN_IN;
  assign n39394 = ~n39387 & ~n37023;
  assign n43709 = ~n40693;
  assign n27702 = ~n35861 & ~n27695;
  assign n31795 = ~n31684 & ~n24813;
  assign n31960 = ~n31718;
  assign n27705 = ~n35861;
  assign n37476 = ~n34580 | ~n34409;
  assign n35594 = ~P3_EAX_REG_28__SCAN_IN | ~n34808;
  assign n27754 = ~n27654 | ~n27653;
  assign n26064 = ~n26063 & ~n33714;
  assign n40375 = ~n40374 | ~n40373;
  assign n35465 = ~n35473;
  assign n26048 = ~n31382 | ~n35473;
  assign n41338 = ~n41328 & ~n41327;
  assign n36078 = P3_INSTADDRPOINTER_REG_8__SCAN_IN & n36077;
  assign n41335 = ~n41353 & ~n41334;
  assign n44023 = ~n43300;
  assign n43719 = ~n43718;
  assign n36867 = ~n39387 & ~n41408;
  assign n40652 = ~n39481 & ~n39480;
  assign n35940 = ~n41105 | ~n35658;
  assign n31821 = ~n33474;
  assign n43915 = ~n43813;
  assign n39387 = ~n36227 | ~n40221;
  assign n42090 = ~n41495 | ~n27886;
  assign n24129 = ~n24128 | ~n24127;
  assign n36077 = ~n27347 | ~n22937;
  assign n41327 = ~n41371 & ~n41326;
  assign n41496 = ~n41495 & ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n26062 = ~n43712 & ~n33714;
  assign n43707 = ~n43358;
  assign n31684 = ~n31681 & ~n24811;
  assign n34808 = ~n43942 & ~n34335;
  assign n34404 = ~n34401 & ~n34400;
  assign n31722 = ~n32110;
  assign n37486 = ~n38058;
  assign n26204 = ~n26203 & ~n26202;
  assign n24562 = ~n34569 | ~n33710;
  assign n43809 = ~n43924;
  assign n24479 = ~n36136 & ~P1_STATE2_REG_0__SCAN_IN;
  assign n43718 = ~n43296 | ~n43295;
  assign n34495 = ~n31913 | ~n32234;
  assign n38482 = ~n36136 & ~n34409;
  assign n41912 = ~P2_STATE2_REG_0__SCAN_IN & ~n43912;
  assign n35967 = ~n43525;
  assign n39302 = ~n34569 | ~n36136;
  assign n41326 = ~n36056 | ~n36055;
  assign n35658 = ~n41401 | ~n35656;
  assign n26047 = ~n31717;
  assign n41333 = ~n41371 & ~n41329;
  assign n28323 = ~n39756;
  assign n31681 = ~n24803 & ~n43722;
  assign n24401 = ~n24400;
  assign n38334 = ~n39531;
  assign n28338 = ~n40935;
  assign n34335 = ~P3_EAX_REG_26__SCAN_IN | ~n33208;
  assign n28819 = ~n28818 | ~n28817;
  assign n39481 = ~n28199 | ~n28198;
  assign n31913 = ~n31906 & ~n31905;
  assign n40270 = ~n40171 | ~n40167;
  assign n28088 = ~n27651 & ~n27650;
  assign n40373 = ~n40382 | ~n40167;
  assign n44091 = ~n44028;
  assign n40372 = ~n40451;
  assign n33262 = ~n32938 & ~n33739;
  assign n34651 = ~n27914 | ~n27913;
  assign n28199 = ~n27889 & ~n27888;
  assign n40762 = ~n27883 | ~n28062;
  assign n44003 = ~n31818 | ~n28153;
  assign n33917 = n27907 & n27906;
  assign n35601 = n28242 & n28241;
  assign n35431 = ~n28235 | ~n28234;
  assign n33208 = ~n43947 & ~n32794;
  assign n28226 = ~n27921 | ~n27920;
  assign n39453 = ~n39449 & ~n39448;
  assign n28093 = ~n41516 & ~n28758;
  assign n28764 = ~n28758 & ~n41119;
  assign n31820 = n31818 & n31817;
  assign n41245 = ~n28746 | ~n28745;
  assign n25073 = ~n31904;
  assign n36205 = n28255 & n28254;
  assign n35970 = ~n28248 | ~n28247;
  assign n27344 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN | ~n35989;
  assign n37264 = n28295 & n28294;
  assign n41329 = ~n35669 & ~n35668;
  assign n24803 = ~n34551 & ~n24802;
  assign n40935 = ~n28337 | ~n28336;
  assign n27893 = n26543 & n26542;
  assign n35656 = ~n35535 | ~n35534;
  assign n24336 = ~n24333;
  assign n39920 = ~n28330 | ~n28329;
  assign n36257 = ~n26536 | ~n26535;
  assign n41223 = ~n28344 | ~n28343;
  assign n39756 = ~n28322 | ~n28321;
  assign n27923 = ~n31714;
  assign n35261 = ~n27900 | ~n27899;
  assign n41732 = ~n28352 | ~n28351;
  assign n35249 = n26529 & n26528;
  assign n41078 = ~n37329 | ~P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n28315 = ~n28313 & ~n28312;
  assign n28657 = ~n28656 | ~n28655;
  assign n27921 = ~n27919 & ~n27918;
  assign n28308 = ~n28306 & ~n28305;
  assign n27900 = ~n27898 & ~n27897;
  assign n28715 = ~n43046 & ~n43725;
  assign n28235 = ~n28233 & ~n28232;
  assign n26529 = ~n26526 & ~n26525;
  assign n39448 = ~n39405 | ~n39404;
  assign n27907 = ~n27905 & ~n27904;
  assign n24811 = ~n31682 & ~n24810;
  assign n28242 = ~n28240 & ~n28239;
  assign n26543 = ~n26541 & ~n26540;
  assign n28275 = ~n28273 & ~n28272;
  assign n28281 = ~n28279 & ~n28278;
  assign n39727 = ~n26495 & ~n26494;
  assign n31818 = ~n28150 | ~n28149;
  assign n28268 = ~n28266 & ~n28265;
  assign n27889 = ~n27882 | ~n27881;
  assign n28288 = ~n28286 & ~n28285;
  assign n28295 = ~n28293 & ~n28292;
  assign n26536 = ~n26534 & ~n26533;
  assign n28147 = ~n28146 & ~n28145;
  assign n38595 = ~n40168 | ~n39404;
  assign n28261 = ~n28259 & ~n28258;
  assign n34966 = ~n32839 & ~n32838;
  assign n43293 = ~n28816 & ~n28885;
  assign n28301 = ~n28299 & ~n28298;
  assign n28758 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN | ~n41231;
  assign n28746 = ~n27648 & ~n27647;
  assign n35989 = ~n27346 | ~n27345;
  assign n28255 = ~n28253 & ~n28252;
  assign n28248 = ~n28246 & ~n28245;
  assign n27914 = ~n27911 & ~n27910;
  assign n36046 = ~n36039 & ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n28322 = ~n28320 & ~n28319;
  assign n36045 = ~n36044 & ~n36043;
  assign n41342 = ~n35612 & ~n35611;
  assign n31361 = ~n31927 | ~n44102;
  assign n32938 = ~n32752 | ~P3_EBX_REG_11__SCAN_IN;
  assign n32794 = ~P3_EAX_REG_24__SCAN_IN | ~n32792;
  assign n35935 = ~n35945;
  assign n23647 = n26515 ^ n26514;
  assign n23615 = ~n23613;
  assign n41005 = ~n41540 | ~n40125;
  assign n33951 = ~n33116 & ~n33619;
  assign n35532 = ~n41156 | ~n34641;
  assign n28299 = ~n28361 & ~n29511;
  assign n28286 = ~n28361 & ~n29493;
  assign n32792 = ~n32489 & ~n32494;
  assign n23642 = ~n23640 & ~n23639;
  assign n35527 = ~P3_EBX_REG_27__SCAN_IN & ~n34656;
  assign n32752 = ~n32716 & ~n33066;
  assign n31927 = ~n31909;
  assign n40508 = ~n41540 | ~n40442;
  assign n35744 = ~n27873 | ~n27872;
  assign n28279 = ~n28361 & ~n36380;
  assign n28293 = ~n28361 & ~n28289;
  assign n28266 = ~n28361 & ~n28262;
  assign n41345 = ~n35269 | ~n35268;
  assign n41231 = ~n27633 | ~n27632;
  assign n27346 = ~n27341 & ~n36021;
  assign n28150 = ~n31524;
  assign n36043 = ~n36042 | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n28834 = ~n28614 & ~n28613;
  assign n35951 = ~n34626 & ~n33772;
  assign n26202 = ~n26201 | ~n27872;
  assign n32838 = ~P3_EAX_REG_8__SCAN_IN | ~n32330;
  assign n27882 = ~n27879 & ~n27878;
  assign n23613 = ~n23574 & ~n23573;
  assign n28816 = ~n28714 | ~P1_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n31682 = ~n24808 | ~n24807;
  assign n35667 = ~n36038 & ~n35664;
  assign n28107 = ~n28144 & ~n28143;
  assign n26201 = ~n26190 & ~n26189;
  assign n32871 = ~P3_EBX_REG_31__SCAN_IN & ~n32865;
  assign n28043 = n28042 & n28041;
  assign n23622 = ~n23633;
  assign n23629 = ~n23625 | ~n23624;
  assign n35944 = ~n35642;
  assign n28613 = ~n28860 & ~n43725;
  assign n36509 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN & ~n40968;
  assign n36333 = ~n35459;
  assign n28714 = n28654 & P1_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n35462 = ~n34843;
  assign n42322 = ~n42320 & ~n40968;
  assign n32716 = ~n32680 | ~P3_EBX_REG_9__SCAN_IN;
  assign n36038 = ~n40968 & ~n35609;
  assign n24444 = ~n24443;
  assign n34659 = ~n33923 & ~n34625;
  assign n36967 = ~n36871;
  assign n32330 = ~n32328 & ~n32566;
  assign n27879 = ~n26493 | ~n26492;
  assign n31322 = ~n31286;
  assign n31344 = ~n31817;
  assign n27872 = ~n31765 | ~n26431;
  assign n32494 = ~n32606 | ~n32608;
  assign n32680 = ~n32678 & ~n33620;
  assign n34655 = ~P3_EBX_REG_25__SCAN_IN & ~n33906;
  assign n28143 = ~P2_PHYADDRPOINTER_REG_26__SCAN_IN | ~n28108;
  assign n26205 = ~n26181 | ~n23127;
  assign n28041 = ~n28040 & ~n28039;
  assign n36338 = n32475 & n34968;
  assign n36239 = ~n34968 | ~n32472;
  assign n25573 = ~n25572;
  assign n34536 = ~n33075 | ~n33630;
  assign n26189 = ~n23532 | ~n23531;
  assign n26492 = ~n26491 & ~n26490;
  assign n23515 = ~n23514 | ~n31525;
  assign n31817 = ~n31196 | ~n43061;
  assign n32865 = ~n34611;
  assign n36022 = n27339 & n27340;
  assign n36243 = ~n34968;
  assign n36871 = ~n41403 | ~n41520;
  assign n26514 = ~n26518;
  assign n34673 = ~n34671 | ~n40724;
  assign n28654 = n28612 & P1_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n28612 = n28459 & P1_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n40125 = ~n40422 & ~n42320;
  assign n28152 = ~n28151 & ~n32149;
  assign n28039 = ~n28038 | ~n28037;
  assign n32861 = ~n32859 & ~n32858;
  assign n33906 = ~n33801 | ~n40544;
  assign n40872 = ~n36221 & ~n41095;
  assign n36242 = ~n33090 & ~n32489;
  assign n28414 = ~n28737 & ~n43725;
  assign n35930 = ~n35942;
  assign n27340 = ~n27338 & ~n27337;
  assign n33630 = ~n33515 & ~n33514;
  assign n36154 = ~n35947;
  assign n23621 = ~n23618 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n28108 = ~n43539 & ~n28142;
  assign n34340 = ~n33792 | ~n33791;
  assign n24441 = ~n24503 & ~n32083;
  assign n36153 = ~n41325 & ~n32870;
  assign n26181 = ~n27870 | ~n26180;
  assign n23514 = ~n23506 & ~n35802;
  assign n23722 = ~n26207;
  assign n34671 = ~n34638 & ~n34637;
  assign n36490 = ~n26475 | ~n26474;
  assign n24340 = ~n24230 | ~n24229;
  assign n26493 = ~n26488 & ~n26487;
  assign n31196 = ~n31200;
  assign n31202 = ~n31200 & ~n35802;
  assign n41520 = ~n41400;
  assign n32671 = ~n32251 & ~n33527;
  assign n33801 = ~P3_EBX_REG_23__SCAN_IN & ~n33802;
  assign n23588 = ~n23583;
  assign n34638 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN & ~n34979;
  assign n24252 = ~n24435 | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n27337 = ~n40191 & ~n36927;
  assign n26489 = ~n26192 & ~n26191;
  assign n28459 = n28413 & P1_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n36019 = ~n27679 | ~n27678;
  assign n42320 = ~n41537;
  assign n32870 = ~n32869 | ~n33500;
  assign n32372 = ~n32371 & ~n32370;
  assign n34637 = ~n33898 & ~n34979;
  assign n26180 = ~n31057 | ~n36364;
  assign n32849 = ~n32848 | ~n33500;
  assign n35947 = ~P3_STATE2_REG_3__SCAN_IN | ~n33496;
  assign n23717 = ~n23710 | ~n23709;
  assign n31273 = ~n26046 | ~n44102;
  assign n27338 = ~n27335 & ~n27336;
  assign n27973 = ~n42174 & ~n43725;
  assign n36660 = ~n40734 | ~n40731;
  assign n33496 = ~n34626;
  assign n27028 = ~n27027 | ~n27026;
  assign n33310 = ~n32550 | ~n32549;
  assign n28413 = n28036 & P1_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n41403 = ~n41100 | ~n40734;
  assign n33802 = ~n33823 | ~n39502;
  assign n26198 = ~n26197 & ~n26434;
  assign n27679 = ~n36913 | ~P3_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n23265 = ~n23222 | ~n23221;
  assign n33500 = ~n34626 & ~n40527;
  assign n26477 = ~n26448 & ~n26447;
  assign n34979 = ~n41401;
  assign n28109 = ~n28141 & ~n28140;
  assign n32251 = ~n31955 | ~n31954;
  assign n24431 = ~n24430;
  assign n26478 = ~n26457 & ~n26456;
  assign n32550 = ~n24175 | ~n24174;
  assign n31777 = ~n23719 | ~n23085;
  assign n23263 = ~n26445;
  assign n40734 = ~n37753;
  assign n27678 = ~n27677 | ~n27676;
  assign n28036 = P1_PHYADDRPOINTER_REG_22__SCAN_IN & n27972;
  assign n31920 = ~n24148 & ~n24147;
  assign n31911 = ~n34509 & ~n31910;
  assign n41531 = ~n40857;
  assign n32202 = ~n32860 & ~n32197;
  assign n33823 = ~P3_EBX_REG_21__SCAN_IN & ~n33824;
  assign n25554 = ~n25553;
  assign n23596 = ~n23595 & ~n23594;
  assign n28265 = ~n28264 | ~n28263;
  assign n28239 = ~n28238 | ~n28237;
  assign n26331 = ~n26330 & ~n36840;
  assign n23719 = ~n26545;
  assign n28258 = ~n28257 | ~n28256;
  assign n23926 = ~n23922 | ~n23921;
  assign n26679 = ~n26678 | ~n26677;
  assign n31894 = ~n24125 | ~n24142;
  assign n28232 = ~n28231 | ~n28230;
  assign n24174 = ~n24173 | ~n31697;
  assign n26445 = ~n23281 | ~n23282;
  assign n24175 = ~n31794 | ~n40081;
  assign n27918 = ~n27917 | ~n27916;
  assign n27972 = n26982 & P1_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n33824 = ~n33953 | ~n37324;
  assign n26525 = ~n26524 | ~n26523;
  assign n28245 = ~n28244 | ~n28243;
  assign n27617 = ~n27615 & ~n27614;
  assign n31276 = ~n31448 | ~n26045;
  assign n27330 = ~n36970 & ~n36969;
  assign n27910 = ~n27909 | ~n27908;
  assign n23219 = n23180 & n23179;
  assign n32200 = ~n31671 & ~n31665;
  assign n27904 = ~n27903 | ~n27902;
  assign n26533 = ~n26532 | ~n26531;
  assign n23628 = ~n23627 | ~n23626;
  assign n27676 = ~n27675 | ~n27674;
  assign n27813 = ~n32373 | ~n27812;
  assign n28252 = ~n28251 | ~n28250;
  assign n26980 = ~n41899 & ~n43725;
  assign n27897 = ~n27896 | ~n27895;
  assign n28110 = ~n28139 & ~n28138;
  assign n26456 = ~n26444 | ~n26462;
  assign n24204 = ~n24203 & ~n32337;
  assign n23284 = ~n23281;
  assign n41397 = ~n40743;
  assign n26540 = ~n26539 | ~n26538;
  assign n23595 = ~n23593 & ~n37289;
  assign n40744 = ~n36914 & ~n39615;
  assign n24214 = ~n26044 & ~n33710;
  assign n35377 = ~n25765 | ~n25764;
  assign n27615 = ~n27609 | ~n27612;
  assign n23179 = ~n23178 | ~n23177;
  assign n26330 = ~n26228 & ~n26227;
  assign n26711 = n26636 & n26635;
  assign n33953 = ~P3_EBX_REG_19__SCAN_IN & ~n34986;
  assign n43394 = ~n43393 & ~n43392;
  assign n36374 = ~n25785 | ~n25784;
  assign n39700 = ~n26928 | ~n26927;
  assign n39909 = ~n28172 | ~n28171;
  assign n26982 = ~n26979 & ~n26060;
  assign n32196 = ~n31810 & ~n41374;
  assign n40415 = ~n39451 & ~n40442;
  assign n32263 = ~n25723 | ~n25722;
  assign n28163 = ~n26932 | ~n26931;
  assign n23581 = ~n23580 | ~n23579;
  assign n36830 = ~n25592 | ~n25591;
  assign n26457 = ~n26436 | ~n26435;
  assign n24247 = ~n24245 & ~n24244;
  assign n23180 = ~n23135 & ~n23134;
  assign n35443 = ~n33488;
  assign n37270 = ~n26920 | ~n26919;
  assign n26196 = ~n26195 | ~n26437;
  assign n25540 = ~n25538;
  assign n23922 = ~n23915 | ~n23914;
  assign n25541 = ~n25537 & ~n25538;
  assign n37535 = n25026 & n25025;
  assign n33783 = ~n25751 | ~n25750;
  assign n36828 = ~n25630 | ~n25629;
  assign n32344 = ~n25716 | ~n25715;
  assign n23531 = ~n23530 & ~n23529;
  assign n23716 = ~n23715 | ~n23714;
  assign n36970 = ~n27326 & ~n27325;
  assign n32889 = ~n25571 | ~n25570;
  assign n31824 = ~n41324 & ~n31823;
  assign n28079 = ~n25737 | ~n25736;
  assign n26551 = ~n25675 | ~n25674;
  assign n23177 = ~n23176 & ~n23175;
  assign n39759 = ~n28168 & ~n28167;
  assign n24245 = ~n24233 & ~n24232;
  assign n41208 = ~n28181 & ~n28180;
  assign n34902 = ~n25582 & ~n25581;
  assign n27609 = n27608 & n27607;
  assign n25563 = ~n25561 & ~n25560;
  assign n34986 = ~n34985 | ~n36176;
  assign n23178 = ~n23173 | ~n23172;
  assign n27801 = ~n27800 & ~n27799;
  assign n25722 = ~n25721 & ~n25720;
  assign n25764 = ~n25763 & ~n25762;
  assign n37464 = ~n26924 & ~n26923;
  assign n23134 = ~n23133 & ~n23132;
  assign n26913 = ~n25789 & ~n25788;
  assign n25736 = ~n25735 & ~n25734;
  assign n23135 = ~n23176 & ~n26193;
  assign n26979 = ~n26637 | ~P1_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n41472 = ~n28195 & ~n28194;
  assign n35316 = ~n25771 & ~n25770;
  assign n25026 = ~n25022 & ~n25021;
  assign n23914 = ~n23913 | ~n23912;
  assign n27325 = ~n36667 & ~n36666;
  assign n27727 = ~n41147 | ~n27726;
  assign n26137 = ~n26136 | ~n26135;
  assign n31534 = ~n31533 & ~n31532;
  assign n25063 = ~n25060 & ~n22944;
  assign n40442 = ~n40422;
  assign n41927 = ~n28190 & ~n28189;
  assign n25113 = ~n36249 & ~n43091;
  assign n37499 = ~n24949 & ~n22945;
  assign n26459 = ~n26439 | ~n26438;
  assign n37444 = ~n25780 & ~n25779;
  assign n33555 = ~n25744 & ~n25743;
  assign n32799 = ~n25730 & ~n25729;
  assign n23492 = ~n23544;
  assign n31670 = ~n32361 | ~n31532;
  assign n26228 = n32944 & n32945;
  assign n24244 = ~n24243 | ~n24242;
  assign n25839 = ~n25835 | ~n25834;
  assign n23218 = ~n26434 | ~n23564;
  assign n23696 = ~n23695;
  assign n27717 = ~n41147 & ~n27716;
  assign n27733 = ~n41147 | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n25750 = ~n25749 & ~n25748;
  assign n34835 = ~n25757 & ~n25756;
  assign n26227 = P2_INSTADDRPOINTER_REG_2__SCAN_IN & n26226;
  assign n25060 = ~n22942 & ~n25057;
  assign n24949 = ~n22942 & ~n24943;
  assign n26032 = ~n26029 & ~n26028;
  assign n26981 = ~n26978 & ~n26977;
  assign n36667 = ~n35435 & ~n27321;
  assign n28706 = ~n28616 | ~n28615;
  assign n25730 = ~n25728 | ~n25727;
  assign n25546 = ~n32175;
  assign n25744 = ~n25742 | ~n25741;
  assign n34985 = ~P3_EBX_REG_17__SCAN_IN & ~n34531;
  assign n41362 = ~n31790 | ~n31789;
  assign n41147 = ~n41149;
  assign n25022 = ~n22942 & ~n25018;
  assign n27811 = ~n27810 | ~n27809;
  assign n25539 = ~n25530 | ~n25529;
  assign n26637 = ~n26598 & ~n26059;
  assign n25560 = ~n25559 | ~n25558;
  assign n28415 = ~n28412 & ~n28411;
  assign n27974 = ~n27971 & ~n27970;
  assign n27799 = ~n27798 & ~n31371;
  assign n26135 = ~n26134 | ~n26133;
  assign n27037 = ~n27036 | ~n27035;
  assign n27034 = ~n27033 | ~n27032;
  assign n26688 = ~n26687 | ~n26686;
  assign n23912 = ~n23911 | ~n23919;
  assign n26685 = ~n26684 | ~n26683;
  assign n28050 = ~n28049 | ~n28048;
  assign n26145 = ~n26144 | ~n26143;
  assign n28053 = ~n28052 | ~n28051;
  assign n23176 = ~n26437 & ~n23127;
  assign n23273 = n23272 & n23271;
  assign n26036 = ~n26035 | ~n26034;
  assign n41784 = ~n41783 & ~n41782;
  assign n23925 = ~n23924 & ~n23923;
  assign n28468 = ~n28467 | ~n28466;
  assign n23173 = ~n23170 | ~n26466;
  assign n23688 = ~n23687 & ~n23686;
  assign n25942 = ~n25941 | ~n25940;
  assign n23283 = ~n23282;
  assign n25939 = ~n25938 | ~n25937;
  assign n25844 = ~n25843 | ~n25842;
  assign n28471 = ~n28470 | ~n28469;
  assign n25088 = ~n25087 | ~n25086;
  assign n23656 = ~n23678 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n24243 = ~n24240 & ~n24239;
  assign n25085 = ~n25084 | ~n25083;
  assign n24139 = ~n24240;
  assign n25082 = ~n25081 | ~n25080;
  assign n25757 = ~n25755 | ~n25754;
  assign n25771 = ~n25769 | ~n25768;
  assign n25079 = ~n25078 | ~n25077;
  assign n23549 = ~n23548 & ~n31493;
  assign n27734 = ~n41149 | ~n41002;
  assign n24196 = ~n24195 | ~n24194;
  assign n23915 = ~n23924 | ~n23923;
  assign n26507 = ~n31058 & ~n23127;
  assign n24168 = ~n24167 | ~n24166;
  assign n24187 = ~n24186 | ~n24185;
  assign n24216 = ~n24116 & ~n24115;
  assign n24193 = ~n24192 | ~n24191;
  assign n24181 = ~n24180 | ~n24179;
  assign n24178 = ~n24177 | ~n24176;
  assign n42978 = ~n28824 | ~n28823;
  assign n27731 = ~n41149 | ~n40820;
  assign n24184 = ~n24183 | ~n24182;
  assign n36249 = ~n42796 | ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n24190 = ~n24189 | ~n24188;
  assign n23913 = ~n23905 | ~n23904;
  assign n24839 = ~n24838 & ~n24837;
  assign n26226 = ~n26224 | ~n33564;
  assign n26684 = ~n40080 | ~P1_EBX_REG_18__SCAN_IN;
  assign n23911 = ~n23908 & ~n23907;
  assign n23279 = ~n23512 | ~n23278;
  assign n23921 = ~n23920 | ~n23919;
  assign n26144 = ~n40080 | ~P1_EBX_REG_17__SCAN_IN;
  assign n23924 = ~n23902 | ~n23901;
  assign n25074 = ~n25072 & ~n25071;
  assign n26598 = ~n26093 | ~P1_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n23272 = ~n26168 | ~n23278;
  assign n27681 = ~n27680 | ~P3_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n23221 = ~n23278 | ~n26159;
  assign n24826 = ~n24825 & ~n24824;
  assign n26035 = ~n40080 | ~P1_EBX_REG_16__SCAN_IN;
  assign n27324 = ~n27323 & ~P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n25785 = ~n25783 & ~n25782;
  assign n35435 = ~n35437 & ~n35436;
  assign n24713 = ~n24711;
  assign n24116 = ~n24114 | ~n24113;
  assign n25776 = ~n25774 & ~n25773;
  assign n25675 = ~n25673 & ~n25672;
  assign n24177 = ~n40080 | ~P1_EBX_REG_2__SCAN_IN;
  assign n25716 = ~n25714 & ~n25713;
  assign n26487 = ~n26451 | ~n26450;
  assign n25630 = ~n25628 & ~n25627;
  assign n25742 = ~n25740 & ~n25739;
  assign n24167 = ~n40080 | ~P1_EBX_REG_1__SCAN_IN;
  assign n27816 = ~n32367 | ~n27787;
  assign n24095 = ~n31896 | ~n24094;
  assign n31790 = ~n31787 | ~n41542;
  assign n27878 = ~n27877 | ~n27876;
  assign n25769 = ~n25767 & ~n25766;
  assign n25592 = ~n25590 & ~n25589;
  assign n28615 = ~n28603 & ~n28602;
  assign n28112 = ~n28136 & ~n28135;
  assign n24334 = ~n24332 & ~n24331;
  assign n34531 = ~n33848 | ~n35420;
  assign n25578 = ~n25577 | ~n25576;
  assign n25934 = ~n25894 | ~n25893;
  assign n26031 = ~n41025 & ~n43725;
  assign n25530 = ~n25493 | ~n25492;
  assign n42318 = ~n40980;
  assign n25552 = ~n25549 & ~n25548;
  assign n25755 = ~n25753 & ~n25752;
  assign n32175 = ~n25543 | ~n25542;
  assign n25728 = ~n25726 & ~n25725;
  assign n25571 = ~n25569 & ~n25568;
  assign n23687 = ~n23685 & ~n23684;
  assign n23928 = ~n23895 | ~n23894;
  assign n23175 = ~n23174 | ~n23507;
  assign n26466 = ~n23169 | ~n23168;
  assign n23670 = ~n23685 & ~n35718;
  assign n37468 = ~n41873 & ~n28205;
  assign n31907 = ~n24199 & ~n35466;
  assign n24849 = ~n24848 & ~n24847;
  assign n23920 = ~n23918 | ~n23917;
  assign n27669 = ~n27668 | ~P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n24837 = ~n24836 & ~n24835;
  assign n25720 = ~n25719 | ~n25718;
  assign n23559 = ~n23703 | ~n23564;
  assign n23946 = ~n24101 | ~n23945;
  assign n23901 = ~n24655 | ~n24100;
  assign n24824 = ~n24823 | ~n24822;
  assign n24142 = ~n24124 & ~n24234;
  assign n24779 = ~n24777 & ~n24776;
  assign n25072 = ~n25068 | ~n31793;
  assign n40586 = ~n41873 & ~n28202;
  assign n27674 = ~n27673 | ~P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n23594 = ~n23703 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n32082 = ~n24199;
  assign n24800 = ~n24799 & ~n24798;
  assign n23660 = ~n23659;
  assign n31896 = ~n24162 | ~n31895;
  assign n24814 = ~n24794 | ~n24793;
  assign n23558 = ~n26505 & ~n36357;
  assign n25543 = ~n25758 | ~n34885;
  assign n41546 = ~n40202 & ~n39615;
  assign n27888 = ~n41873 & ~n27880;
  assign n40606 = ~n41873 & ~n28201;
  assign n25535 = ~n25534 | ~n25533;
  assign n25529 = ~n25758 | ~n26440;
  assign n41212 = ~n41873 & ~n41213;
  assign n26093 = ~n26058 & ~n41023;
  assign n28604 = ~n43286;
  assign n25557 = ~n26914 & ~n25544;
  assign n23216 = ~n26505 & ~n26327;
  assign n27342 = ~n32515 & ~n27333;
  assign n25581 = ~n25580 | ~n25579;
  assign n33848 = ~P3_EBX_REG_15__SCAN_IN & ~n33666;
  assign n26462 = ~n22939 | ~n26443;
  assign n33564 = ~n33563 | ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n25930 = ~n25929 | ~n25928;
  assign n23278 = ~n33357;
  assign n24331 = ~n24330 | ~n24329;
  assign n28135 = ~P2_PHYADDRPOINTER_REG_16__SCAN_IN | ~n28113;
  assign n39927 = ~n41873 & ~n28207;
  assign n34498 = ~n24201 & ~n24208;
  assign n32177 = ~n26176 | ~n26175;
  assign n23491 = ~n23520 & ~n25544;
  assign n24239 = ~n24238 | ~n24237;
  assign n32367 = ~n31671 & ~n41375;
  assign n35437 = ~n27318 | ~n27317;
  assign n24611 = ~n24608 & ~n24607;
  assign n23565 = ~n23564 | ~n36795;
  assign n27597 = ~n31801 & ~n27795;
  assign n27814 = ~n31801 & ~n31808;
  assign n23543 = ~n25491 & ~n36795;
  assign n27329 = ~n27328 & ~P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n37735 = ~n41873 & ~n28204;
  assign n25713 = ~n26916 & ~n31210;
  assign n27606 = ~n27605 | ~n22936;
  assign n27326 = ~n27322 & ~n38732;
  assign n24911 = n24910 & n24909;
  assign n24731 = ~n24730 & ~n24729;
  assign n24114 = ~n24111 | ~n24110;
  assign n24711 = ~n24709 & ~n24708;
  assign n24986 = n24985 & n24984;
  assign n24172 = ~n24170 & ~n24169;
  assign n39210 = ~n41873 & ~n28203;
  assign n27664 = ~n27663 | ~P3_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n39480 = ~n41873 & ~n28200;
  assign n31787 = ~n31808;
  assign n24947 = ~n24946 | ~n24945;
  assign n26429 = ~n23127 & ~n26428;
  assign n31910 = ~n31448 | ~n31478;
  assign n25893 = ~n25892 | ~n25891;
  assign n40738 = ~n38909 & ~n38910;
  assign n24847 = ~n24846 | ~n24845;
  assign n24708 = ~n24872 & ~n24707;
  assign n24482 = ~n24872 & ~n24480;
  assign n22944 = ~n25059 | ~n25058;
  assign n27802 = ~n32206 & ~n32868;
  assign n31788 = ~n27807 & ~n27806;
  assign n24559 = ~n24872 & ~n28592;
  assign n27787 = ~n27786 | ~n27785;
  assign n26916 = ~n41474;
  assign n23902 = ~n23896 & ~n34097;
  assign n24835 = ~n24834 | ~n24833;
  assign n27629 = ~n27628 & ~n30706;
  assign n23919 = ~n23910 & ~n23909;
  assign n24162 = ~n24092 & ~n24207;
  assign n24657 = ~n24664 | ~n24654;
  assign n35819 = ~n24868 | ~n24867;
  assign n24608 = ~n24872 & ~n24576;
  assign n31525 = ~n31770;
  assign n24857 = ~n24856 | ~n24855;
  assign n24165 = ~n28825 | ~n24235;
  assign n33666 = ~n33688 | ~n34400;
  assign n26058 = ~n26030 | ~P1_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n26385 = ~n23127 & ~n26384;
  assign n27322 = ~n27250 | ~n27249;
  assign n25025 = n25024 & n25023;
  assign n23577 = ~n23576 & ~n23575;
  assign n31808 = ~n27806 | ~n27791;
  assign n24389 = ~n24388 | ~n24387;
  assign n28113 = ~n28134 & ~n28133;
  assign n24166 = ~n40081 | ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n27331 = ~n27327 & ~n38589;
  assign n27612 = ~n27611 | ~n27792;
  assign n31793 = ~n40081;
  assign n24778 = ~n36688 | ~n39522;
  assign n27619 = ~n27626 & ~n27618;
  assign n23449 = ~n23415 | ~n25093;
  assign n24807 = ~n24806 & ~n24805;
  assign n25094 = ~n23730;
  assign n23652 = ~n36688 & ~n36357;
  assign n31895 = ~n24093 & ~n44100;
  assign n23524 = ~n25544 & ~n36779;
  assign n24909 = n24908 & n24907;
  assign n25834 = n25833 & n25832;
  assign n24984 = n24983 & n24982;
  assign n25928 = ~n24872 | ~n24871;
  assign n24794 = ~n24817 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23889 = ~n24405 | ~n23851;
  assign n23703 = ~n25544 | ~n43061;
  assign n26224 = ~n26223 | ~n26440;
  assign n23262 = ~n23085 | ~n26341;
  assign n24332 = ~n24872 & ~n26099;
  assign n31809 = ~n31806 & ~n31805;
  assign n26285 = ~n26225 & ~n23127;
  assign n22904 = ~n23415;
  assign n31498 = ~n37289 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n24654 = ~n24706;
  assign n31806 = ~n31804 | ~n32472;
  assign n33915 = ~n25717;
  assign n27655 = ~n27671 & ~n32208;
  assign n24211 = ~n31721 & ~n24210;
  assign n23503 = ~n36561 | ~n36795;
  assign n25024 = ~n43721 | ~P1_EAX_REG_11__SCAN_IN;
  assign n24817 = ~n24831;
  assign n27785 = ~n27784 | ~n31666;
  assign n24867 = ~n24866 & ~n24865;
  assign n24207 = ~n25069 | ~n34149;
  assign n24161 = ~n25068 | ~n34097;
  assign n23576 = ~n36561 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n24237 = ~n24236 & ~n35474;
  assign n24234 = ~n31715 & ~n32239;
  assign n26178 = ~n26177 & ~P2_STATE2_REG_1__SCAN_IN;
  assign n27332 = ~n27250 & ~n32208;
  assign n24822 = ~n24821 & ~n24820;
  assign n23934 = ~n24706 & ~n24097;
  assign n25838 = ~n40490 & ~n43725;
  assign n33688 = ~P3_EBX_REG_13__SCAN_IN & ~n33741;
  assign n24119 = ~n32239 & ~n24392;
  assign n23447 = ~n23415 | ~n36561;
  assign n24221 = ~n32239 | ~n24392;
  assign n24481 = ~n24871 & ~n24563;
  assign n24111 = ~n24109 | ~n34226;
  assign n27661 = ~n35976 | ~n35975;
  assign n24709 = ~n24733 & ~n24706;
  assign n32206 = ~n32672 & ~n35267;
  assign n26030 = ~n25889 & ~n41128;
  assign n33585 = ~n34885 & ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n27791 = ~n27790 | ~n27789;
  assign n35436 = ~n27319 | ~n27320;
  assign n27866 = ~n42353 & ~n41072;
  assign n24775 = ~n43061 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n25892 = ~n43721 | ~P1_EAX_REG_15__SCAN_IN;
  assign n24560 = ~n24706 & ~n24565;
  assign n27596 = ~n27595 & ~n27594;
  assign n23728 = ~n37289;
  assign n23545 = ~n43061 | ~n37289;
  assign n27628 = ~n27627 | ~n32489;
  assign n23497 = ~n36779 & ~n36795;
  assign n24793 = ~n24792 & ~n24791;
  assign n28133 = ~P2_PHYADDRPOINTER_REG_14__SCAN_IN | ~n28114;
  assign n26225 = ~n34885 | ~n26440;
  assign n24395 = ~n24394 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n36202 = ~n25759;
  assign n27618 = ~n30706 & ~n22935;
  assign n24297 = ~n24477 & ~n24296;
  assign n31511 = ~n32868 | ~n27610;
  assign n24330 = ~n24727 | ~n24489;
  assign n23513 = ~n23511 | ~n23510;
  assign n28114 = ~n28132 & ~n28131;
  assign n31666 = ~n31825 | ~n32198;
  assign n40052 = ~n26826 & ~n26825;
  assign n24396 = ~n24393 & ~n24397;
  assign n35974 = ~n33095 & ~P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n27250 = ~n32826 | ~n32808;
  assign n37119 = ~n25391 & ~n25390;
  assign n24871 = ~n24727;
  assign n27666 = ~n27657;
  assign n27592 = ~n27604 | ~n27803;
  assign n24112 = ~n24802 & ~n24392;
  assign n35267 = ~n32475 & ~n32472;
  assign n32868 = ~n33487 | ~n32860;
  assign n27789 = ~n27788 & ~n27804;
  assign n32199 = ~n41375 & ~n32198;
  assign n27599 = ~n27616 | ~n32475;
  assign n34097 = ~n39891;
  assign n26327 = ~n23215 & ~n23214;
  assign n27775 = ~n27774 & ~n27788;
  assign n27630 = ~n32475 & ~n27626;
  assign n26449 = ~n25623 & ~n25622;
  assign n37754 = ~n38140 & ~n32883;
  assign n43721 = ~n28810;
  assign n26173 = ~n26166 & ~n26165;
  assign n24102 = ~n24100 & ~n24099;
  assign n25932 = ~n24873;
  assign n24831 = ~n39895 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n24236 = ~n24235 | ~n44099;
  assign n25889 = ~n25885 | ~P1_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n31804 = ~n31803 & ~n32489;
  assign n38968 = ~n26753 & ~n26752;
  assign n38013 = ~n25454 & ~n25453;
  assign n22900 = ~n43061;
  assign n41789 = ~n26870 & ~n26869;
  assign n35858 = ~n39615;
  assign n25235 = ~n25234 & ~n25233;
  assign n34134 = ~n24392;
  assign n27658 = ~n32284 | ~n27656;
  assign n25236 = ~n25222 & ~n25221;
  assign n38140 = ~n37575 | ~P3_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n23120 = ~n23119 | ~n23118;
  assign n23445 = ~n23444 | ~n23443;
  assign n23214 = ~n23213 | ~n23212;
  assign n43475 = ~n43432 | ~n43431;
  assign n23511 = ~n26168 & ~n23509;
  assign n25266 = ~n25250 | ~n25249;
  assign n25146 = ~n25129 | ~n25128;
  assign n23166 = ~n23165 & ~n23164;
  assign n27616 = ~n30706 | ~n31801;
  assign n25623 = ~n25604 | ~n25603;
  assign n27604 = ~n32672 & ~n31802;
  assign n32489 = ~n32672;
  assign n27796 = ~n33501 | ~n31801;
  assign n27626 = ~n31802;
  assign n24802 = ~n34149;
  assign n24150 = ~n34164;
  assign n34226 = ~n31891;
  assign n25885 = ~n25837 & ~n25836;
  assign n32848 = ~n33501 & ~n33487;
  assign n34187 = ~n23848;
  assign n25206 = ~n25190 | ~n25189;
  assign n27803 = ~n30706 & ~n32475;
  assign n28131 = ~P2_PHYADDRPOINTER_REG_12__SCAN_IN | ~n28115;
  assign n24393 = ~n24391 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n32860 = ~n33501;
  assign n33738 = ~P3_EBX_REG_11__SCAN_IN & ~n33124;
  assign n25668 = ~n25651 & ~n25650;
  assign n23260 = ~n23241 | ~n23240;
  assign n24135 = ~n31891 | ~n31382;
  assign n23167 = n23152 & n23151;
  assign n25190 = ~n25182 & ~n25181;
  assign n23848 = ~n23847 | ~n22929;
  assign n25651 = ~n25640 | ~n25639;
  assign n23121 = ~n23102 | ~n23101;
  assign n23241 = ~n23237 & ~n23236;
  assign n25205 = ~n25204 | ~n25203;
  assign n23119 = ~n23113 & ~n23112;
  assign n24097 = ~n23936 & ~n23933;
  assign n27180 = ~n27164 & ~n27163;
  assign n23384 = ~n23370 | ~n23369;
  assign n24658 = ~n24606 & ~n24605;
  assign n24980 = ~n24979 & ~n24978;
  assign n31193 = ~U212;
  assign n25265 = ~n25264 | ~n25263;
  assign n23215 = ~n23201 | ~n23200;
  assign n25691 = ~n25684 & ~n25683;
  assign n25296 = ~n25295 & ~n25294;
  assign n28115 = ~n42070 & ~n28130;
  assign n25667 = ~n25666 & ~n25665;
  assign n25527 = ~n25526 & ~n25525;
  assign n23259 = ~n23258 | ~n23257;
  assign n25297 = ~n25282 & ~n25281;
  assign n25128 = ~n25127 & ~n25126;
  assign n27781 = ~n27771 & ~n27764;
  assign n24943 = ~n24942 & ~n24941;
  assign n34149 = ~n24091 & ~n24090;
  assign n23165 = ~n23161 | ~n23160;
  assign n23213 = ~n23209 & ~n23208;
  assign n25175 = ~n25174 & ~n25173;
  assign n25709 = ~n25708 | ~n25707;
  assign n37575 = ~n37016 & ~n32882;
  assign n25604 = ~n25600 & ~n25599;
  assign n24392 = ~n23888 | ~n22940;
  assign n41790 = ~n26907 | ~n26906;
  assign n25622 = ~n25621 | ~n25620;
  assign n27659 = ~n27315 & ~n27314;
  assign n25145 = ~n25144 | ~n25143;
  assign n23787 = ~n23786;
  assign n27773 = ~n27769 | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n25250 = ~n25242 & ~n25241;
  assign n24905 = ~n24904 & ~n24903;
  assign n27213 = ~n27197 | ~n27196;
  assign n27143 = ~n27127 | ~n27126;
  assign n27764 = ~n27763 & ~n27762;
  assign n23240 = ~n23239 & ~n23238;
  assign n23236 = ~n23235 | ~n23234;
  assign n24568 = ~n24558 | ~n24557;
  assign n27499 = ~n27498 | ~n27497;
  assign n27769 = ~n27768 | ~n27770;
  assign n27281 = ~n27265 | ~n27264;
  assign n27142 = ~n27141 | ~n27140;
  assign n28130 = ~P2_PHYADDRPOINTER_REG_10__SCAN_IN | ~n27929;
  assign n27470 = ~n27454 | ~n27453;
  assign n27590 = ~n27574 | ~n27573;
  assign n37016 = ~n36873 | ~P3_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n23257 = ~n23256 & ~n23255;
  assign n24653 = ~n24637 | ~n24636;
  assign n24704 = ~n24703 | ~n24702;
  assign n24475 = ~n24474 | ~n24473;
  assign n23258 = ~n23250 & ~n23249;
  assign n24476 = ~n24460 | ~n24459;
  assign n23300 = ~n23299 | ~n23298;
  assign n24605 = ~n24604 | ~n24603;
  assign n25189 = ~n25188 & ~n25187;
  assign n23102 = ~n23094 & ~n23093;
  assign n25640 = ~n25633 & ~n25632;
  assign n25620 = ~n25619 & ~n25618;
  assign n23101 = ~n23100 & ~n23099;
  assign n25621 = ~n25613 & ~n25612;
  assign n23113 = ~n23109 | ~n23108;
  assign n25264 = ~n25258 & ~n25257;
  assign n25684 = ~n25680 | ~n25679;
  assign n23432 = ~n23424 & ~n23423;
  assign n25249 = ~n25248 & ~n25247;
  assign n24328 = ~n24312 | ~n24311;
  assign n27197 = ~n27189 & ~n27188;
  assign n25708 = ~n25700 & ~n25699;
  assign n25666 = ~n25662 | ~n25661;
  assign n25707 = ~n25706 & ~n25705;
  assign n24606 = ~n24590 | ~n24589;
  assign n24327 = ~n24326 | ~n24325;
  assign n25204 = ~n25196 & ~n25195;
  assign n27078 = ~n27077 | ~n27076;
  assign n23152 = ~n23144 & ~n23143;
  assign n25143 = ~n25142 & ~n25141;
  assign n25144 = ~n25140 & ~n25139;
  assign n23151 = ~n23150 & ~n23149;
  assign n23474 = ~n23462 & ~n23461;
  assign n25129 = ~n25121 & ~n25120;
  assign n27112 = ~n27093 | ~n27092;
  assign n25161 = ~n25160 & ~n25159;
  assign n24652 = ~n24651 | ~n24650;
  assign n25600 = ~n25596 | ~n25595;
  assign n25203 = ~n25202 & ~n25201;
  assign n25528 = ~n25513 & ~n25512;
  assign n23200 = ~n23199 & ~n23198;
  assign n27163 = ~n27162 | ~n27161;
  assign n27247 = ~n27227 | ~n27226;
  assign n24705 = ~n24689 | ~n24688;
  assign n33067 = ~P3_EBX_REG_9__SCAN_IN & ~n33622;
  assign n25526 = ~n25522 | ~n25521;
  assign U212 = ~n31063 | ~U214;
  assign n23201 = ~n23193 & ~n23192;
  assign n24016 = ~n24000 & ~n23999;
  assign n24689 = ~n24681 & ~n24680;
  assign n23192 = ~n23191 | ~n23190;
  assign n24688 = ~n24687 & ~n24686;
  assign n24703 = ~n24695 & ~n24694;
  assign n23269 = ~n23266 | ~n38277;
  assign n23255 = ~n23254 | ~n23253;
  assign n23256 = ~n23252 | ~n23251;
  assign n23249 = ~n23248 | ~n23247;
  assign n24651 = ~n24643 & ~n24642;
  assign n23461 = ~n23460 | ~n23459;
  assign n23318 = ~n23317 | ~n23316;
  assign n23164 = ~n23163 | ~n23162;
  assign n24636 = ~n24635 & ~n24634;
  assign n23093 = ~n23092 | ~n23091;
  assign n23100 = ~n23096 | ~n23095;
  assign n23099 = ~n23098 | ~n23097;
  assign n23423 = ~n23422 | ~n23421;
  assign n23393 = ~n23392 | ~n23391;
  assign n24603 = ~n24602 & ~n24601;
  assign n27077 = ~n27065 & ~n27064;
  assign n27423 = ~n27422 & ~n27421;
  assign n24325 = ~n24324 & ~n24323;
  assign n27439 = ~n27438 | ~n27437;
  assign n27164 = ~n27150 | ~n27149;
  assign n23785 = ~n23776 & ~n23775;
  assign n27162 = ~n27156 & ~n27155;
  assign n25699 = ~n25698 | ~n25697;
  assign n27454 = ~n27446 & ~n27445;
  assign n25706 = ~n25702 | ~n25701;
  assign n27246 = ~n27245 | ~n27244;
  assign n24295 = ~n24273 & ~n24272;
  assign n24589 = ~n24588 & ~n24587;
  assign n23784 = ~n23783 & ~n23782;
  assign n24386 = ~n24362 & ~n24361;
  assign n27111 = ~n27110 | ~n27109;
  assign n24385 = ~n24384 & ~n24383;
  assign n27092 = ~n27091 & ~n27090;
  assign n27772 = ~n27771 | ~n27770;
  assign n24312 = ~n24304 & ~n24303;
  assign n27763 = ~n27767 & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n27189 = ~n27186 | ~n27185;
  assign n27196 = ~n27195 & ~n27194;
  assign n27762 = ~n27761 | ~n27770;
  assign n24294 = ~n24293 & ~n24292;
  assign n27212 = ~n27211 | ~n27210;
  assign n24326 = ~n24318 & ~n24317;
  assign n27589 = ~n27588 | ~n27587;
  assign n24474 = ~n24466 & ~n24465;
  assign n27558 = ~n27550 & ~n27549;
  assign n24590 = ~n24582 & ~n24581;
  assign n27500 = ~n27484 | ~n27483;
  assign n27264 = ~n27263 & ~n27262;
  assign n25661 = ~n25660 & ~n25659;
  assign n27560 = ~n27544 | ~n27543;
  assign n25665 = ~n25664 | ~n25663;
  assign n27127 = ~n27119 & ~n27118;
  assign n27929 = ~n28129 & ~n28128;
  assign n27394 = ~n27386 & ~n27385;
  assign n24459 = ~n24458 & ~n24457;
  assign n27530 = ~n27514 | ~n27513;
  assign n27378 = ~n27370 & ~n27369;
  assign n27265 = ~n27257 & ~n27256;
  assign n27497 = ~n27496 & ~n27495;
  assign n27528 = ~n27520 & ~n27519;
  assign n24460 = ~n24452 & ~n24451;
  assign n27280 = ~n27279 | ~n27278;
  assign n27141 = ~n27133 & ~n27132;
  assign n25512 = ~n25511 | ~n25510;
  assign n36873 = ~n36222 & ~n33842;
  assign n25522 = ~n25516 & ~n25515;
  assign n27469 = ~n27468 | ~n27467;
  assign n27574 = ~n27566 & ~n27565;
  assign n25650 = ~n25649 | ~n25648;
  assign n24557 = ~n24556 & ~n24555;
  assign n31063 = ~n36558 & ~n23017;
  assign n25525 = ~n25524 | ~n25523;
  assign n24075 = ~n24067 & ~n24066;
  assign n25513 = ~n25503 | ~n25502;
  assign n27179 = n27178 & n27177;
  assign n24558 = ~n24536 & ~n24535;
  assign n23462 = ~n23457 & ~n35715;
  assign n23209 = ~n23205 | ~n23204;
  assign n24293 = ~n24281 | ~n24280;
  assign n23879 = ~n23875 | ~n23874;
  assign n27093 = ~n27085 & ~n27084;
  assign n27064 = ~n27063 | ~n27062;
  assign n27076 = ~n27075 & ~n27074;
  assign n23473 = ~n23472 & ~n23471;
  assign n23118 = ~n23117 & ~n23116;
  assign n25649 = ~n25643 & ~n25642;
  assign n36558 = ~n36557;
  assign n24465 = ~n24464 | ~n24463;
  assign n24582 = ~n24578 | ~n24577;
  assign n25648 = ~n25647 & ~n25646;
  assign n23844 = ~n23840 | ~n23839;
  assign n24066 = ~n24065 | ~n24064;
  assign n28128 = ~P2_PHYADDRPOINTER_REG_8__SCAN_IN | ~n28116;
  assign n24458 = ~n24454 | ~n24453;
  assign n24074 = ~n24073 & ~n24072;
  assign n23846 = ~n23838 & ~n23837;
  assign n25521 = ~n25520 & ~n25519;
  assign n24452 = ~n24448 | ~n24447;
  assign n39901 = ~n39896;
  assign n24555 = ~n24554 | ~n24553;
  assign n24650 = ~n24649 & ~n24648;
  assign n24536 = ~n24524 | ~n24523;
  assign n24088 = ~n24087 & ~n24086;
  assign n27056 = ~n27055 & ~n27054;
  assign n24604 = ~n24596 & ~n24595;
  assign n27057 = ~n27047 & ~n27046;
  assign n24635 = ~n24631 | ~n24630;
  assign n24272 = ~n24271 | ~n24270;
  assign n25603 = ~n25602 & ~n25601;
  assign n24000 = ~n23989 | ~n23988;
  assign n23161 = ~n23157 & ~n23156;
  assign n25618 = ~n25617 | ~n25616;
  assign n24634 = ~n24633 | ~n24632;
  assign n24855 = n24854 & n24853;
  assign n25690 = ~n25689 & ~n25688;
  assign n25700 = ~n25696 | ~n25695;
  assign n25698 = ~n26852 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n25702 = ~n26831 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n23775 = ~n23774 | ~n23773;
  assign n25701 = ~n26837 | ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n25705 = ~n25704 | ~n25703;
  assign n27245 = ~n27237 & ~n27236;
  assign n24273 = ~n24262 | ~n24261;
  assign n24588 = ~n24584 | ~n24583;
  assign n23783 = ~n23779 | ~n23778;
  assign n25503 = ~n25497 & ~n25496;
  assign n24643 = ~n24639 | ~n24638;
  assign n25502 = ~n25501 & ~n25500;
  assign n27219 = ~n27215 | ~n27214;
  assign n25511 = ~n25505 & ~n25504;
  assign n25510 = ~n25509 & ~n25508;
  assign n25639 = ~n25638 & ~n25637;
  assign n24473 = ~n24472 & ~n24471;
  assign n27150 = ~n27148 & ~n27147;
  assign n27437 = ~n27436 & ~n27435;
  assign n23337 = ~n23333 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n27438 = ~n27430 & ~n27429;
  assign n27421 = ~n27420 | ~n27419;
  assign n24324 = ~n24320 | ~n24319;
  assign n36222 = ~n36182 | ~P3_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n23254 = ~n26827 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n24317 = ~n24316 | ~n24315;
  assign n23251 = ~n26837 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n23252 = ~n26831 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n23248 = ~n26852 | ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n27210 = ~n27209 & ~n27208;
  assign n27424 = ~n27416 & ~n27415;
  assign n23394 = ~n23390 & ~n35715;
  assign n27211 = ~n27203 & ~n27202;
  assign n24311 = ~n24310 & ~n24309;
  assign n23250 = ~n23246 | ~n23245;
  assign n27195 = ~n27191 | ~n27190;
  assign n27767 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~n27760;
  assign n27186 = ~n27184 & ~n27183;
  assign n24304 = ~n24300 | ~n24299;
  assign n27133 = ~n27129 | ~n27128;
  assign n27407 = ~n27406 & ~n27405;
  assign n27408 = ~n27400 & ~n27399;
  assign n27565 = ~n27564 | ~n27563;
  assign n27140 = ~n27139 & ~n27138;
  assign n27573 = ~n27572 & ~n27571;
  assign n27126 = ~n27125 & ~n27124;
  assign n27393 = ~n27392 & ~n27391;
  assign n27385 = ~n27384 | ~n27383;
  assign n24512 = ~n24511 | ~n24510;
  assign n27588 = ~n27580 & ~n27579;
  assign n27119 = ~n27116 | ~n27115;
  assign n27587 = ~n27586 & ~n27585;
  assign n27514 = ~n27506 & ~n27505;
  assign n27496 = ~n27492 | ~n27491;
  assign n27513 = ~n27512 & ~n27511;
  assign n27519 = ~n27518 | ~n27517;
  assign n27527 = ~n27526 & ~n27525;
  assign n42522 = ~n42698;
  assign n27498 = ~n27490 & ~n27489;
  assign n27364 = ~n27356 & ~n27355;
  assign n27483 = ~n27482 & ~n27481;
  assign n27363 = ~n27362 & ~n27361;
  assign n27257 = ~n27254 | ~n27253;
  assign n27369 = ~n27368 | ~n27367;
  assign n27377 = ~n27376 & ~n27375;
  assign n27544 = ~n27536 & ~n27535;
  assign n27484 = ~n27476 & ~n27475;
  assign n27543 = ~n27542 & ~n27541;
  assign n27263 = ~n27259 | ~n27258;
  assign n27550 = ~n27546 | ~n27545;
  assign n27177 = ~n27176 & ~n27175;
  assign n27557 = ~n27556 & ~n27555;
  assign n27467 = ~n27466 & ~n27465;
  assign n27468 = ~n27460 & ~n27459;
  assign n23931 = ~n23930 | ~n23929;
  assign n27279 = ~n27271 & ~n27270;
  assign n24680 = ~n24679 | ~n24678;
  assign n27178 = ~n27170 & ~n27169;
  assign n27453 = ~n27452 & ~n27451;
  assign n24702 = ~n24701 & ~n24700;
  assign n27278 = ~n27277 & ~n27276;
  assign n27161 = ~n27160 & ~n27159;
  assign n27155 = ~n27154 & ~n27153;
  assign n27091 = ~n27087 | ~n27086;
  assign n24362 = ~n24350 | ~n24349;
  assign n23306 = ~n23305 | ~n23304;
  assign n23212 = ~n23211 & ~n23210;
  assign n27109 = ~n27108 & ~n27107;
  assign n23268 = ~n23267 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23362 = ~n23358 & ~n35715;
  assign n23431 = ~n23430 & ~n23429;
  assign n24637 = ~n24629 & ~n24628;
  assign n24981 = ~n24944 & ~n37241;
  assign n27110 = ~n27102 & ~n27101;
  assign n23424 = ~n23420 & ~n35715;
  assign n27361 = ~n27360 | ~n27359;
  assign n27585 = ~n27584 | ~n27583;
  assign n27225 = ~n27221 | ~n27220;
  assign n27586 = ~n27582 | ~n27581;
  assign n27218 = ~n27217 | ~n27216;
  assign n27579 = ~n27578 | ~n27577;
  assign n25509 = ~n25507 | ~n25506;
  assign n27506 = ~n27502 | ~n27501;
  assign n27505 = ~n27504 | ~n27503;
  assign n27525 = ~n27524 | ~n27523;
  assign n27370 = ~n27366 | ~n27365;
  assign n27520 = ~n27516 | ~n27515;
  assign n23782 = ~n23781 | ~n23780;
  assign n27362 = ~n27358 | ~n27357;
  assign n27215 = ~n22919 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n27224 = ~n27223 | ~n27222;
  assign n23916 = ~n24098;
  assign n24472 = ~n24468 | ~n24467;
  assign n27511 = ~n27510 | ~n27509;
  assign n27116 = n27114 & n27113;
  assign n27356 = ~n27352 | ~n27351;
  assign n27526 = ~n27522 | ~n27521;
  assign n27512 = ~n27508 | ~n27507;
  assign n27355 = ~n27354 | ~n27353;
  assign n27580 = ~n27576 | ~n27575;
  assign n24471 = ~n24470 | ~n24469;
  assign n27376 = ~n27372 | ~n27371;
  assign n24086 = ~n24085 | ~n24084;
  assign n27436 = ~n27432 | ~n27431;
  assign n24535 = ~n24534 | ~n24533;
  assign n24087 = ~n24083 | ~n24082;
  assign n27435 = ~n27434 | ~n27433;
  assign n24523 = ~n24522 & ~n24521;
  assign n27276 = ~n27275 | ~n27274;
  assign n24524 = ~n24519 & ~n24518;
  assign n27277 = ~n27273 | ~n27272;
  assign n27445 = ~n27444 | ~n27443;
  assign n24079 = ~n43245 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n27270 = ~n27269 | ~n27268;
  assign n24025 = ~n24024 & ~n24023;
  assign n23929 = ~n23893 | ~n23892;
  assign n27271 = ~n27267 | ~n27266;
  assign n27460 = ~n27456 | ~n27455;
  assign n24553 = ~n24552 & ~n24551;
  assign n24081 = ~n24077 | ~n24076;
  assign n27262 = ~n27261 | ~n27260;
  assign n27259 = ~n22919 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n27476 = ~n27472 | ~n27471;
  assign n27475 = ~n27474 | ~n27473;
  assign n27482 = ~n27478 | ~n27477;
  assign n24448 = ~n22907 | ~P1_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n27481 = ~n27480 | ~n27479;
  assign n24556 = ~n24546 | ~n24545;
  assign n27490 = ~n27486 | ~n27485;
  assign n24447 = ~n28775 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n27489 = ~n27488 | ~n27487;
  assign n24451 = ~n24450 | ~n24449;
  assign n24073 = ~n24069 | ~n24068;
  assign n27495 = ~n27494 | ~n27493;
  assign n28116 = ~n28127 & ~n28126;
  assign n24064 = ~n43265 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n27386 = ~n27382 | ~n27381;
  assign n24454 = ~n43245 | ~P1_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n27138 = ~n27137 | ~n27136;
  assign n24457 = ~n24456 | ~n24455;
  assign n27139 = ~n27135 | ~n27134;
  assign n27392 = ~n27388 | ~n27387;
  assign n27391 = ~n27390 | ~n27389;
  assign n27400 = ~n27396 | ~n27395;
  assign n27132 = ~n27131 | ~n27130;
  assign n27399 = ~n27398 | ~n27397;
  assign n27129 = ~n22919 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n24466 = ~n24462 | ~n24461;
  assign n27406 = ~n27402 | ~n27401;
  assign n23843 = ~n23842 | ~n23841;
  assign n27405 = ~n27404 | ~n27403;
  assign n27124 = ~n27123 | ~n27122;
  assign n27566 = ~n27562 | ~n27561;
  assign n27125 = ~n27121 | ~n27120;
  assign n24463 = ~n43265 | ~P1_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n25519 = ~n25518 | ~n25517;
  assign n27571 = ~n27570 | ~n27569;
  assign n27074 = ~n27073 | ~n27072;
  assign n24318 = ~n24314 | ~n24313;
  assign n27208 = ~n27207 | ~n27206;
  assign n27209 = ~n27205 | ~n27204;
  assign n27202 = ~n27201 | ~n27200;
  assign n23878 = ~n23877 | ~n23876;
  assign n27203 = ~n27199 | ~n27198;
  assign n24309 = ~n24308 | ~n24307;
  assign n24310 = ~n24306 | ~n24305;
  assign n27194 = ~n27193 | ~n27192;
  assign n24303 = ~n24302 | ~n24301;
  assign n24281 = ~n24277 & ~n24276;
  assign n27191 = ~n22919 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n24299 = ~n22907 | ~P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n24300 = ~n28775 | ~P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n27184 = ~n33191 & ~n27181;
  assign n24384 = ~n24372 | ~n24371;
  assign n27107 = ~n27106 | ~n27105;
  assign n27085 = ~n27081 | ~n27080;
  assign n27108 = ~n27104 | ~n27103;
  assign n24292 = ~n24291 | ~n24290;
  assign n27102 = ~n27099 | ~n27098;
  assign n27084 = ~n27083 | ~n27082;
  assign n27090 = ~n27089 | ~n27088;
  assign n27087 = ~n22919 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n27375 = ~n27374 | ~n27373;
  assign n24262 = ~n24257 & ~n24256;
  assign n25704 = ~n22906 | ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n27536 = ~n27532 | ~n27531;
  assign n27237 = ~n27234 | ~n27233;
  assign n27535 = ~n27534 | ~n27533;
  assign n25695 = ~n26841 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n27542 = ~n27538 | ~n27537;
  assign n27175 = ~n27174 | ~n27173;
  assign n27541 = ~n27540 | ~n27539;
  assign n27243 = ~n27239 | ~n27238;
  assign n27176 = ~n27172 | ~n27171;
  assign n23776 = ~n23771 | ~n23770;
  assign n25688 = ~n25687 & ~n25686;
  assign n25689 = ~n26820 & ~n25685;
  assign n27549 = ~n27548 | ~n27547;
  assign n27242 = ~n27241 | ~n27240;
  assign n27556 = ~n27552 | ~n27551;
  assign n25683 = ~n25682 | ~n25681;
  assign n25680 = ~n25678 & ~n25677;
  assign n27555 = ~n27554 | ~n27553;
  assign n27169 = ~n27168 | ~n27167;
  assign n27170 = ~n27166 | ~n27165;
  assign n27159 = ~n33298 & ~n27158;
  assign n27160 = ~n33191 & ~n27157;
  assign n29835 = ~U215;
  assign n27156 = ~n27152 & ~n27151;
  assign n27147 = ~n34766 & ~n27146;
  assign n27148 = ~n27145 | ~n27144;
  assign n25596 = ~n25594 & ~n25593;
  assign n24271 = ~n24266 & ~n24265;
  assign n27047 = ~n27043 | ~n27042;
  assign n23815 = ~n23814 | ~n23813;
  assign n27046 = ~n27045 | ~n27044;
  assign n27055 = ~n27051 | ~n27050;
  assign n23756 = ~n23751 & ~n23750;
  assign n24056 = ~n24055 & ~n24054;
  assign n27054 = ~n27053 | ~n27052;
  assign n24323 = ~n24322 | ~n24321;
  assign n24319 = ~n43265 | ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n27065 = ~n27060 | ~n27059;
  assign n27063 = ~n22919 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n24316 = ~n43245 | ~P1_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n27075 = ~n27067 | ~n27066;
  assign n23058 = ~n23057 & ~n23056;
  assign n23205 = ~n23203 & ~n23202;
  assign n23072 = ~n22906 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n24628 = ~n24627 | ~n24626;
  assign n23116 = ~n26820 & ~n23115;
  assign n23457 = ~n23456 & ~n23455;
  assign n23109 = ~n23107 & ~n23106;
  assign n22926 = ~n22925;
  assign n23094 = ~n23090 | ~n23089;
  assign n23472 = ~n23466 | ~n23465;
  assign n23156 = ~n23155 | ~n23154;
  assign n23471 = ~n23470 | ~n23469;
  assign n23476 = ~n22906 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n24944 = ~n24906 | ~P1_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n24642 = ~n24641 | ~n24640;
  assign n23479 = ~n23478 | ~n23477;
  assign n24649 = ~n24645 | ~n24644;
  assign n24648 = ~n24647 | ~n24646;
  assign n25659 = ~n25658 | ~n25657;
  assign n25662 = ~n25655 & ~n25654;
  assign n23989 = ~n23983 & ~n23982;
  assign n23034 = ~n23030 | ~n23029;
  assign n23390 = ~n23389 & ~n23388;
  assign n23024 = ~n23023 & ~n23022;
  assign n23400 = ~n23396 | ~n23395;
  assign n23399 = ~n23398 | ~n23397;
  assign n23341 = ~n22906 | ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n23333 = ~n23332 | ~n23331;
  assign n23327 = ~n23326 | ~n23325;
  assign n23405 = ~n22905 & ~n37805;
  assign n23328 = ~n23324 | ~n23323;
  assign n24681 = ~n24677 | ~n24676;
  assign n23408 = ~n22906 | ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n23420 = ~n23419 & ~n23418;
  assign n23430 = ~n23426 | ~n23425;
  assign n23429 = ~n23428 | ~n23427;
  assign n23988 = ~n23987 & ~n23986;
  assign n23434 = ~n22906 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n23358 = ~n23357 & ~n23356;
  assign n24511 = ~n39311 | ~n24508;
  assign n23368 = ~n23364 | ~n23363;
  assign n23367 = ~n23366 | ~n23365;
  assign n23999 = ~n23998 | ~n23997;
  assign n23253 = ~n26841 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n26827 = ~n25687;
  assign n26837 = ~n26818;
  assign n26831 = ~n25495;
  assign n23305 = ~n23303 & ~n23302;
  assign n26852 = ~n25634;
  assign n23246 = ~n23244 & ~n23243;
  assign n23239 = ~n22905 & ~n42786;
  assign n23237 = ~n23233 | ~n23232;
  assign n27429 = ~n27428 | ~n27427;
  assign n23961 = ~n23957 | ~n23956;
  assign n37853 = ~n41310 & ~n23654;
  assign n30874 = ~n30030;
  assign n36182 = ~n32881 & ~n32880;
  assign n24026 = ~n24020 & ~n24019;
  assign n27416 = ~n27412 | ~n27411;
  assign n27415 = ~n27414 | ~n27413;
  assign n27422 = ~n27418 | ~n27417;
  assign n27430 = ~n27426 | ~n27425;
  assign n24006 = ~n24002 | ~n24001;
  assign n24581 = ~n24580 | ~n24579;
  assign n24005 = ~n24004 | ~n24003;
  assign n23038 = ~n22906 | ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n25637 = ~n25636 | ~n25635;
  assign n23233 = ~n23231 & ~n23230;
  assign n23335 = ~n22924 | ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n24554 = ~n24549 & ~n24548;
  assign n29304 = ~n29305;
  assign n23331 = ~n22911 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n23023 = ~n23021 | ~n23020;
  assign n23032 = ~n23467 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n23029 = ~n23464 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n24261 = ~n24260 & ~n24259;
  assign n24533 = ~n24532 & ~n24531;
  assign n24534 = ~n24529 & ~n24528;
  assign n23030 = ~n23463 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n23026 = ~n22924 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n24629 = ~n24625 | ~n24624;
  assign n24545 = ~n24544 & ~n24543;
  assign n24450 = ~n43246 | ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n24449 = ~n43242 | ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n39311 = ~n34718 | ~n24507;
  assign n28126 = ~P2_PHYADDRPOINTER_REG_6__SCAN_IN | ~n28117;
  assign n24456 = ~n43251 | ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n24462 = ~n43274 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n24461 = ~n43270 | ~P1_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n23016 = ~n23015 & ~n23014;
  assign n24464 = ~n22908 | ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n24468 = ~n43275 | ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n24467 = ~n43264 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n24470 = ~n43261 | ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n26841 = ~n25641;
  assign n43880 = ~n28156;
  assign n23324 = ~n23463 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n39188 = ~n39115 | ~n39114;
  assign n23323 = ~n23464 | ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n23326 = ~n23467 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n25696 = ~n25694 & ~n25693;
  assign n23332 = n23330 & n23329;
  assign n25682 = ~n26858 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n25677 = ~n26791 & ~n43512;
  assign n27471 = ~n22913 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n24322 = ~n22908 | ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n28934 = ~n28930;
  assign n24320 = ~n43270 | ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n24315 = ~n43261 | ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n23893 = ~n23891 | ~n23890;
  assign n24313 = ~n43264 | ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n24314 = ~n43275 | ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n24307 = ~n43242 | ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n27432 = ~n36294 | ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n27427 = ~n22913 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n24308 = ~n43251 | ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n27419 = ~n22914 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n24306 = ~n43274 | ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n24301 = ~n43260 | ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n24302 = ~n43246 | ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n27758 = ~n27765 | ~n27766;
  assign n28775 = ~n24515;
  assign n39279 = ~n38617 | ~n39114;
  assign n27474 = ~n22914 | ~P3_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n42524 = ~n42291 & ~n42282;
  assign n27354 = ~n22914 | ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n27522 = ~n22913 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n27517 = ~n22914 | ~P3_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n27371 = ~n22913 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n27532 = ~n22914 | ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n27534 = ~n22913 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n27575 = ~n22920 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n27576 = ~n22913 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n27567 = ~n22914 | ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n27404 = ~n36320 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n27401 = ~n22914 | ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n27395 = ~n22913 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n24291 = ~n24285 & ~n24284;
  assign n24280 = ~n24279 & ~n24278;
  assign n24439 = ~n37485 | ~n24508;
  assign n24270 = ~n24269 & ~n24268;
  assign n23654 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~n37542;
  assign n35805 = ~n32149;
  assign n41877 = ~n38321 | ~n28197;
  assign n24290 = ~n24289 & ~n24288;
  assign n24020 = ~n24515 & ~n24017;
  assign n27275 = ~n22914 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n27272 = ~n22910 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n27268 = ~n22913 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n24019 = ~n24517 & ~n24018;
  assign n27266 = ~n36320 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n24023 = ~n27011 & ~n24022;
  assign n27267 = ~n22909 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n27261 = ~n36317 | ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n24035 = ~n24030 & ~n24029;
  assign n27253 = ~n22912 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n27136 = ~n22912 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n27134 = ~n22923 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n27130 = ~n22917 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n27131 = ~n22914 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n27128 = ~n22910 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n27122 = ~n36320 | ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n27123 = ~n22909 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n27120 = ~n22913 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n23983 = ~n24515 & ~n23980;
  assign n24906 = ~n24861 & ~n34823;
  assign n23982 = ~n24517 & ~n23981;
  assign n23986 = ~n27011 & ~n23985;
  assign n23998 = ~n23993 & ~n23992;
  assign n27089 = ~n35392 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n27086 = ~n22914 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n23854 = ~n24515 & ~n23853;
  assign n27082 = ~n22913 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n27083 = ~n36310 | ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n27080 = ~n22917 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n23869 = ~n27004 & ~n23866;
  assign n32845 = ~n41145 & ~n42023;
  assign n27072 = ~n22913 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n27067 = ~n36320 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n27062 = ~n22923 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n27059 = ~n36307 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n27060 = ~n22917 | ~P3_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n27052 = ~n22920 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n27053 = ~n35392 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n27050 = ~n36317 | ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n23751 = ~n24515 & ~n27010;
  assign n27044 = ~n22914 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n27045 = ~n36298 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n23750 = ~n24517 & ~n23749;
  assign n27042 = ~n36310 | ~P3_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n23755 = ~n23754 & ~n23753;
  assign n23814 = ~n23810 & ~n23809;
  assign n27043 = ~n36294 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n23766 = ~n23760 & ~n23759;
  assign n23765 = ~n23764 & ~n23763;
  assign n27241 = ~n22920 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n27238 = ~n36307 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n27239 = ~n22914 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n27233 = ~n36320 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n27234 = ~n27232 & ~n27231;
  assign n27222 = ~n35392 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n27223 = ~n22917 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n27220 = ~n36317 | ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n23792 = ~n27004 & ~n24377;
  assign n27216 = ~n22913 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n27217 = ~n36298 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n27214 = ~n22923 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n24065 = ~n22908 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n24069 = ~n43275 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n24068 = ~n43264 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n24072 = ~n24071 | ~n24070;
  assign n23821 = ~n27011 & ~n26096;
  assign n24077 = ~n43251 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n24076 = ~n43246 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n23819 = ~n24517 & ~n24275;
  assign n23820 = ~n24515 & ~n24255;
  assign n24078 = ~n43242 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n24085 = ~n43274 | ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n24546 = ~n24541 & ~n24540;
  assign n24047 = ~n24041 & ~n24040;
  assign n27173 = ~n22920 | ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n27174 = ~n22917 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n27171 = ~n22914 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n27172 = ~n36298 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n27167 = ~n22923 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n27168 = ~n36310 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n27165 = ~n36317 | ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n27149 = ~n36294 | ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n24046 = ~n24045 & ~n24044;
  assign n24057 = ~n24051 & ~n24050;
  assign n24055 = ~n27004 & ~n24052;
  assign n27207 = ~n22913 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n27204 = ~n22917 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n27205 = ~n36298 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n27200 = ~n36320 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n27201 = ~n36307 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n27198 = ~n22923 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n27192 = ~n22914 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n27193 = ~n36317 | ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n27190 = ~n22920 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n23855 = ~n24517 & ~n23852;
  assign n29461 = ~n29058;
  assign n27105 = ~n36307 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n27106 = ~n36298 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n27103 = ~n22923 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n27098 = ~n36320 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n27099 = ~n27097 & ~n27096;
  assign n27088 = ~n22920 | ~P3_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n27728 = ~n39775 | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n23419 = ~n23417 | ~n23416;
  assign n23422 = ~n23458 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n23426 = ~n23463 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n23425 = ~n23464 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n23428 = ~n23467 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n23470 = ~n23467 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n23433 = ~n26832 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n23465 = ~n23464 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n26818 = ~n23463;
  assign n23466 = ~n23463 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n23304 = ~n22911 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n23357 = ~n23354 | ~n23353;
  assign n23456 = ~n23454 | ~n23453;
  assign n43711 = ~n43469 | ~P1_REIP_REG_31__SCAN_IN;
  assign n43367 = ~n43729;
  assign n23360 = ~n22924 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n43361 = ~n43469 | ~P1_REIP_REG_30__SCAN_IN;
  assign n23965 = ~n43251 | ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n23364 = ~n23463 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n23960 = ~n23959 | ~n23958;
  assign n23293 = ~n25645 & ~n43086;
  assign n23956 = ~n43264 | ~P1_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n23460 = ~n22924 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n43137 = ~n43469 | ~P1_REIP_REG_29__SCAN_IN;
  assign n23389 = ~n23387 | ~n23386;
  assign n23392 = ~n23458 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n23064 = ~n23463 | ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n23060 = ~n23458 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n23396 = ~n23463 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n23395 = ~n23464 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n22906 = ~n25645;
  assign n23475 = ~n26832 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n28943 = ~n28937;
  assign n23398 = ~n23467 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n23953 = ~n22908 | ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n23066 = ~n23467 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n23063 = ~n23464 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n23407 = ~n26832 | ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n23057 = ~n23055 | ~n23054;
  assign n23754 = ~n32121 & ~n23752;
  assign n23858 = ~n24527 & ~n23857;
  assign n24249 = ~n29568 & ~n34677;
  assign n28156 = ~n26214 | ~n39508;
  assign n24507 = ~n24506 | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n24469 = ~n22915 | ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n34718 = ~n38481 | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n23880 = ~n22915 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n23753 = ~n24539 & ~n27003;
  assign n24305 = ~n43271 | ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n23868 = ~n32121 & ~n23867;
  assign n23805 = ~n26659 & ~n24368;
  assign n23810 = ~n28585 & ~n24364;
  assign n23864 = ~n28591 & ~n23863;
  assign n23865 = ~n28585 & ~n23862;
  assign n23809 = ~n24539 & ~n24342;
  assign n23825 = ~n26659 & ~n24264;
  assign n24455 = ~n43271 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n23826 = ~n28591 & ~n24267;
  assign n23822 = ~n27009 & ~n24287;
  assign n43246 = ~n32121;
  assign n37485 = ~n24437 & ~n24505;
  assign n39016 = ~n38220 | ~n39114;
  assign n24070 = ~n43271 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n24071 = ~n22915 | ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n43275 = ~n28591;
  assign n23600 = ~n23599 & ~n26214;
  assign n23781 = ~n22915 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n23791 = ~n24527 & ~n24352;
  assign n23796 = ~n24526 & ~n24363;
  assign n24321 = ~n22915 | ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n23763 = ~n24527 & ~n23762;
  assign n22988 = ~n22987 | ~n22986;
  assign n23764 = ~n24526 & ~n23761;
  assign n27236 = ~n27288 & ~n27235;
  assign n23760 = ~n26095 & ~n23757;
  assign n36415 = ~n35995 & ~n32976;
  assign n27766 = ~n27757 | ~n27776;
  assign n23418 = ~n43098 & ~n41631;
  assign n23427 = ~n23468 | ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n23436 = ~n26838 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n23356 = ~n43098 & ~n23355;
  assign n23290 = ~n25652 & ~n43093;
  assign n41374 = ~n42025;
  assign n23997 = ~n23996 & ~n23995;
  assign n23992 = ~n26659 & ~n23991;
  assign n23993 = ~n28591 & ~n23990;
  assign n23987 = ~n27009 & ~n23984;
  assign n23303 = ~n43094 & ~n25605;
  assign n23056 = ~n43098 & ~n23136;
  assign n39775 = ~n40531 & ~n39786;
  assign n23065 = ~n23468 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n24861 = ~n24852 | ~P1_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n23455 = ~n43098 & ~n26298;
  assign n38207 = ~n37851 | ~n39114;
  assign n23959 = ~n22915 | ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n26848 = n43503 & n35715;
  assign n23958 = ~n43271 | ~P1_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n28117 = ~n28125 & ~n28124;
  assign n26858 = ~n25652;
  assign n23478 = ~n26838 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n23469 = ~n23468 | ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n25678 = ~n26789 & ~n25676;
  assign n23859 = ~n24526 & ~n23856;
  assign n24054 = ~n24527 & ~n24053;
  assign n24050 = ~n32121 & ~n24049;
  assign n23325 = ~n23468 | ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n24051 = ~n24526 & ~n24048;
  assign n24044 = ~n24539 & ~n24043;
  assign n24045 = ~n28585 & ~n24042;
  assign n23343 = ~n26838 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n24040 = ~n27006 & ~n24039;
  assign n23022 = ~n43098 & ~n26271;
  assign n24041 = ~n26095 & ~n24038;
  assign n23031 = ~n23468 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n37834 = ~n37610 | ~n39114;
  assign n23388 = ~n43098 & ~n25692;
  assign n24034 = ~n24033 & ~n24032;
  assign n23397 = ~n23468 | ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n24029 = ~n26659 & ~n24028;
  assign n24030 = ~n28591 & ~n24027;
  assign n23410 = ~n26838 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n24024 = ~n27009 & ~n24021;
  assign n22979 = ~n22978 | ~n22977;
  assign n22909 = ~n34042;
  assign n39097 = ~n39028 & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n22910 = ~n27230;
  assign n23017 = ~n22953 | ~n22952;
  assign n23015 = ~n23002 | ~n23001;
  assign n24100 = ~n23900 | ~n23899;
  assign n23014 = ~n23013 | ~n23012;
  assign n22901 = ~n22912;
  assign n27097 = ~n27301 & ~n34767;
  assign n37933 = ~n38220 | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n37542 = ~n39113 & ~n39114;
  assign n24227 = ~n29568 | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n26791 = ~n26862;
  assign n41145 = ~n40865;
  assign n22917 = n36286;
  assign n24250 = ~n39310 & ~n26587;
  assign n22980 = ~n22967 | ~n22966;
  assign n41516 = ~n28757 | ~P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n23329 = ~n43496 | ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n22915 = ~n28593;
  assign n23686 = ~n37852 & ~n39524;
  assign n23827 = ~n28587 & ~n26099;
  assign n23346 = ~n23481 | ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n37851 = ~n37030 & ~n38277;
  assign n23777 = ~n23772;
  assign n22986 = ~n22985 & ~P1_BE_N_REG_1__SCAN_IN;
  assign n23828 = ~n28593 & ~n26094;
  assign n24209 = ~n29574 | ~n29752;
  assign n23020 = ~n43496 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n27240 = ~n36311 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n39529 = ~n37362 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n23671 = ~n37951 & ~n39524;
  assign n39113 = ~n23653 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n26214 = ~n31488;
  assign n42023 = ~n41384 & ~n41382;
  assign n23759 = ~n28587 & ~n23758;
  assign n38220 = ~n37636 & ~n37635;
  assign n22977 = ~n22976 & ~P1_ADDRESS_REG_2__SCAN_IN;
  assign n27927 = ~n31816;
  assign n38481 = ~n24504 & ~n34677;
  assign n27066 = ~n36311 | ~P3_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n23811 = ~n28587 & ~n24355;
  assign n24437 = ~n24436 & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n23620 = ~n23619 & ~P2_STATE2_REG_1__SCAN_IN;
  assign n23123 = ~n23128 | ~n23129;
  assign n22902 = ~n34773;
  assign n23353 = ~n43496 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n22952 = ~n22951 & ~P2_BE_N_REG_0__SCAN_IN;
  assign n42626 = n42214 & P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n23453 = ~n43496 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n24852 = ~n24843 & ~n24842;
  assign n38884 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n37474;
  assign n23377 = ~n23481 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n36289 = ~n27071 & ~n27070;
  assign n23995 = ~n28587 & ~n24480;
  assign n27274 = ~n36311 | ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n23002 = ~n22994 & ~n22993;
  assign n23012 = ~n23011 & ~P2_ADDRESS_REG_2__SCAN_IN;
  assign n23996 = ~n28593 & ~n23994;
  assign n23001 = ~n23000 & ~n22999;
  assign n26807 = ~n23481;
  assign n23899 = ~n23898 | ~n23897;
  assign n22966 = ~n22965 & ~n22964;
  assign n27095 = ~n27049 | ~n27048;
  assign n23054 = ~n43496 | ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n23013 = ~n23008 & ~n23007;
  assign n43094 = ~n43496;
  assign n24033 = ~n28593 & ~n24031;
  assign n35624 = ~n35630 & ~n26050;
  assign n27206 = ~n36311 | ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n23046 = ~n23481 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n23386 = ~n43496 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n23403 = ~n23481 | ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n43033 = ~n31442 | ~n33710;
  assign n22978 = ~n22973 & ~n22972;
  assign n23900 = ~n23849 | ~n39937;
  assign n22967 = ~n22959 & ~n22958;
  assign n23482 = ~n23481 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n28608 = ~n24864;
  assign n27144 = ~n36311 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n23416 = ~n43496 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n36286 = ~n27070 & ~n27058;
  assign n24032 = ~n28587 & ~n24726;
  assign n23439 = ~n23481 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n27776 = ~n27790 | ~n27777;
  assign n23539 = ~n36366;
  assign n22964 = ~n22963 | ~n22962;
  assign n27777 = ~n35608 & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n23122 = ~n37635 | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n44100 = ~n31478;
  assign n34909 = n39508 & P2_STATEBS16_REG_SCAN_IN;
  assign n22972 = ~n22971 | ~n22970;
  assign n22965 = ~n22961 | ~n22960;
  assign n23849 = ~n31922 & ~n23897;
  assign n36048 = ~n36049;
  assign n26587 = ~n32336 | ~n33710;
  assign n22993 = ~n22992 | ~n22991;
  assign n27759 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~n41354;
  assign n22973 = ~n22969 | ~n22968;
  assign n23008 = ~n23004 | ~n23003;
  assign n23000 = ~n22996 | ~n22995;
  assign n27071 = ~n36047;
  assign n22994 = ~n22990 | ~n22989;
  assign n40168 = ~n36526 & ~n36352;
  assign n23850 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~n34677;
  assign n42214 = ~n42651 & ~n42658;
  assign n29574 = ~n29579 | ~n29055;
  assign n23271 = ~n36357 | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n23892 = ~n35163 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n27771 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~n29449;
  assign n29308 = P3_STATE_REG_1__SCAN_IN & n29149;
  assign n40221 = ~n27711;
  assign n22999 = ~n22998 | ~n22997;
  assign n41375 = ~n31667;
  assign n23937 = ~n24830 & ~P1_STATE2_REG_0__SCAN_IN;
  assign n32190 = ~P3_STATE2_REG_0__SCAN_IN & ~n31507;
  assign n22959 = ~n22955 | ~n22954;
  assign n23011 = ~n23010 | ~n23009;
  assign n39524 = ~n39508;
  assign n23103 = ~n23684 & ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n23679 = ~n39508 | ~n39114;
  assign n31938 = ~n31922 & ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n29580 = ~n29055 & ~P1_STATE_REG_0__SCAN_IN;
  assign n38316 = ~n37132 | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n23105 = ~n26878;
  assign n23619 = ~n37634 & ~P2_STATE2_REG_0__SCAN_IN;
  assign n22951 = ~n22950 | ~n22949;
  assign n22976 = ~n22975 | ~n22974;
  assign n22953 = ~n22948 & ~P2_BE_N_REG_1__SCAN_IN;
  assign n22987 = ~n22982 & ~P1_BE_N_REG_0__SCAN_IN;
  assign n22958 = ~n22957 | ~n22956;
  assign n23226 = ~n38277 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n39946 = ~n39315;
  assign n23007 = ~n23006 | ~n23005;
  assign n22985 = ~n22984 | ~n22983;
  assign n24505 = ~n34476 & ~n35163;
  assign n43146 = ~n42996 & ~n42906;
  assign n24843 = ~n24829 | ~P1_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n43612 = ~n43549 & ~n43187;
  assign n37805 = ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n42547 = ~P1_INSTADDRPOINTER_REG_27__SCAN_IN | ~P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n37629 = ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n22996 = ~P2_ADDRESS_REG_8__SCAN_IN & ~P2_ADDRESS_REG_7__SCAN_IN;
  assign n22998 = ~P2_ADDRESS_REG_12__SCAN_IN & ~P2_ADDRESS_REG_11__SCAN_IN;
  assign n42321 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n22997 = ~P2_ADDRESS_REG_14__SCAN_IN & ~P2_ADDRESS_REG_13__SCAN_IN;
  assign n22995 = ~P2_ADDRESS_REG_10__SCAN_IN & ~P2_ADDRESS_REG_9__SCAN_IN;
  assign n22948 = ~P2_M_IO_N_REG_SCAN_IN | ~P2_W_R_N_REG_SCAN_IN;
  assign n43097 = ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n33537 = ~P2_EBX_REG_6__SCAN_IN;
  assign n43082 = ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n23006 = ~P2_ADDRESS_REG_28__SCAN_IN & ~P2_ADDRESS_REG_27__SCAN_IN;
  assign n23005 = ~P2_ADDRESS_REG_1__SCAN_IN & ~P2_ADDRESS_REG_0__SCAN_IN;
  assign n41230 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n26779 = ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n22990 = ~P2_ADDRESS_REG_4__SCAN_IN & ~P2_ADDRESS_REG_3__SCAN_IN;
  assign n43093 = ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n23003 = ~P2_ADDRESS_REG_22__SCAN_IN & ~P2_ADDRESS_REG_21__SCAN_IN;
  assign n22989 = ~P2_ADDRESS_REG_6__SCAN_IN & ~P2_ADDRESS_REG_5__SCAN_IN;
  assign n35254 = ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n23010 = ~P2_ADDRESS_REG_24__SCAN_IN & ~P2_ADDRESS_REG_23__SCAN_IN;
  assign n22992 = ~P2_ADDRESS_REG_16__SCAN_IN & ~P2_ADDRESS_REG_15__SCAN_IN;
  assign n23009 = ~P2_ADDRESS_REG_26__SCAN_IN & ~P2_ADDRESS_REG_25__SCAN_IN;
  assign n22991 = ~P2_ADDRESS_REG_18__SCAN_IN & ~P2_ADDRESS_REG_17__SCAN_IN;
  assign n23004 = ~P2_ADDRESS_REG_20__SCAN_IN & ~P2_ADDRESS_REG_19__SCAN_IN;
  assign n42337 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n22968 = ~P1_ADDRESS_REG_22__SCAN_IN & ~P1_ADDRESS_REG_21__SCAN_IN;
  assign n42786 = ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n22971 = ~P1_ADDRESS_REG_28__SCAN_IN & ~P1_ADDRESS_REG_27__SCAN_IN;
  assign n23104 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n39511 = ~P2_STATE2_REG_2__SCAN_IN;
  assign n28129 = ~P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n36357 = ~P2_STATE2_REG_0__SCAN_IN;
  assign n42070 = ~P2_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n34677 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n38321 = ~P2_STATEBS16_REG_SCAN_IN;
  assign n24707 = ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n22970 = ~P1_ADDRESS_REG_1__SCAN_IN & ~P1_ADDRESS_REG_0__SCAN_IN;
  assign n32075 = ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n28132 = ~P2_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n37475 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n22975 = ~P1_ADDRESS_REG_24__SCAN_IN & ~P1_ADDRESS_REG_23__SCAN_IN;
  assign n23637 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n40527 = ~P3_STATE2_REG_2__SCAN_IN;
  assign n22974 = ~P1_ADDRESS_REG_26__SCAN_IN & ~P1_ADDRESS_REG_25__SCAN_IN;
  assign n39937 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n37634 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n35452 = ~P3_STATE2_REG_1__SCAN_IN;
  assign n22982 = ~P1_M_IO_N_REG_SCAN_IN | ~P1_W_R_N_REG_SCAN_IN;
  assign n32083 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23579 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n22984 = ~P1_D_C_N_REG_SCAN_IN & ~P1_ADS_N_REG_SCAN_IN;
  assign n22983 = ~P1_BE_N_REG_2__SCAN_IN & ~P1_BE_N_REG_3__SCAN_IN;
  assign n37635 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n31055 = ~P2_STATE2_REG_1__SCAN_IN;
  assign n23684 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n33579 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n39114 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n22950 = ~P2_D_C_N_REG_SCAN_IN & ~P2_ADS_N_REG_SCAN_IN;
  assign n41597 = ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n22949 = ~P2_BE_N_REG_2__SCAN_IN & ~P2_BE_N_REG_3__SCAN_IN;
  assign n39944 = ~P1_STATEBS16_REG_SCAN_IN;
  assign n41578 = ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n22955 = ~P1_ADDRESS_REG_4__SCAN_IN & ~P1_ADDRESS_REG_3__SCAN_IN;
  assign n22954 = ~P1_ADDRESS_REG_6__SCAN_IN & ~P1_ADDRESS_REG_5__SCAN_IN;
  assign n24830 = ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n32336 = ~P1_STATE2_REG_1__SCAN_IN & ~P1_STATE2_REG_3__SCAN_IN;
  assign n22957 = ~P1_ADDRESS_REG_16__SCAN_IN & ~P1_ADDRESS_REG_15__SCAN_IN;
  assign n22956 = ~P1_ADDRESS_REG_18__SCAN_IN & ~P1_ADDRESS_REG_17__SCAN_IN;
  assign n22961 = ~P1_ADDRESS_REG_8__SCAN_IN & ~P1_ADDRESS_REG_7__SCAN_IN;
  assign n22960 = ~P1_ADDRESS_REG_10__SCAN_IN & ~P1_ADDRESS_REG_9__SCAN_IN;
  assign n35163 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n23626 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n22963 = ~P1_ADDRESS_REG_12__SCAN_IN & ~P1_ADDRESS_REG_11__SCAN_IN;
  assign n41513 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n22962 = ~P1_ADDRESS_REG_14__SCAN_IN & ~P1_ADDRESS_REG_13__SCAN_IN;
  assign n22969 = ~P1_ADDRESS_REG_20__SCAN_IN & ~P1_ADDRESS_REG_19__SCAN_IN;
  assign n42104 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n29752 = ~P1_STATE_REG_1__SCAN_IN | ~P1_STATE_REG_2__SCAN_IN;
  assign n39440 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n26060 = ~P1_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n23994 = ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n23991 = ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n23990 = ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n23985 = ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n23984 = ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n23981 = ~P1_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n27880 = ~P2_EBX_REG_9__SCAN_IN;
  assign n27235 = ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n41023 = ~P1_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n33714 = ~P1_STATE2_REG_1__SCAN_IN;
  assign n26059 = ~P1_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n33710 = ~P1_STATE2_REG_0__SCAN_IN;
  assign n41128 = ~P1_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n40959 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN | ~P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n42707 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN | ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n40403 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n27048 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n41072 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n35608 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n23980 = ~P1_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n38277 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n35663 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n35728 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n29055 = ~P1_STATE_REG_1__SCAN_IN;
  assign n33933 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n43867 = ~n43864 | ~n43863;
  assign n43895 = ~n43890 | ~n43889;
  assign n43731 = ~n43717 | ~n43716;
  assign n43717 = ~n43708 | ~n43707;
  assign n43342 = n43030 ^ n43029;
  assign n28743 = ~n42832 & ~n43358;
  assign n28866 = ~n42933 & ~n43358;
  assign n43820 = ~n43812 & ~n43811;
  assign n42933 = n28857 ^ P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n42832 = ~n28734 & ~n43028;
  assign n42977 = ~n42976 | ~n42975;
  assign n43651 = ~n43644 | ~n43913;
  assign n43050 = ~n43042 & ~n43358;
  assign n43455 = ~n43453;
  assign n43142 = ~n43135 & ~n43358;
  assign n43705 = ~n43704 | ~n43703;
  assign n28857 = ~n28856 | ~n28855;
  assign n43783 = ~n43776 | ~n43913;
  assign n28492 = ~n42585 & ~n43358;
  assign n43866 = ~n43925 & ~n43893;
  assign n43453 = ~n43449 & ~n43448;
  assign n43529 = ~n43694 | ~n43523;
  assign n43641 = ~n43640 | ~n43639;
  assign n42585 = n42499 ^ n28483;
  assign n28519 = ~n28549 & ~n43358;
  assign n28504 = ~n42371 & ~n43358;
  assign n43640 = ~n43633 | ~n43693;
  assign n43925 = n43865 ^ P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n42487 = ~n42486 & ~n42485;
  assign n42821 = ~n42815 & ~n43358;
  assign n43216 = ~n43223 | ~n43913;
  assign n42974 = ~n42971 | ~n43462;
  assign n43643 = ~n43602 | ~n43746;
  assign n42549 = ~n42972 & ~n43462;
  assign n28510 = ~n28509 & ~n28508;
  assign n28848 = ~n28496 | ~n28852;
  assign n43022 = ~n43014 | ~n43876;
  assign n42486 = ~n42548 & ~n42483;
  assign n43522 = ~n43476 & ~n43475;
  assign n43476 = ~n43395 & ~n43394;
  assign n43806 = ~n43805 | ~n43804;
  assign n43387 = ~n43386 & ~n43385;
  assign n43323 = ~n43316 | ~n43913;
  assign n43201 = ~n43316 | ~n43876;
  assign n42534 = ~n42515 & ~n43755;
  assign n41952 = ~n41951 & ~n41950;
  assign n28895 = ~n28894 | ~n28893;
  assign n28508 = ~n28507 & ~n43462;
  assign n42959 = ~n42952 | ~n43913;
  assign n43598 = ~n43601 | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n41951 = ~n41949 & ~n22933;
  assign n42914 = ~n42952 | ~n43876;
  assign n42916 = ~n42951 & ~n43893;
  assign n43552 = ~n43597 | ~n43809;
  assign n42885 = ~n42800 & ~n43058;
  assign n43592 = ~n43597 | ~n43748;
  assign n42733 = ~n42854 & ~n43893;
  assign n42672 = ~n42840 & ~n43893;
  assign n43383 = ~n43382 | ~n43381;
  assign n27834 = ~n41742 & ~n43358;
  assign n42800 = n42799 & n42798;
  assign n42865 = ~n42855 | ~n43913;
  assign n43057 = ~n43056 & ~n43055;
  assign n42731 = ~n42855 | ~n43876;
  assign n42854 = ~n42710 | ~n42709;
  assign n42840 = ~n42661 | ~n42660;
  assign n43572 = ~n43571 & ~n43794;
  assign n43597 = ~n43170 | ~n43612;
  assign n28873 = ~n28872 | ~n28871;
  assign n43551 = ~n43550 & ~n43549;
  assign n42880 = ~n42869 & ~n43893;
  assign n43024 = ~n43013 & ~n43893;
  assign n42315 = ~n42450 & ~n43893;
  assign n42228 = ~n42422 & ~n43893;
  assign n42297 = ~n42436 & ~n43893;
  assign n43380 = ~n43377 & ~n43794;
  assign n28675 = ~n43377 & ~n44019;
  assign n42822 = ~n43377;
  assign n42536 = ~n42514 | ~n43748;
  assign n28727 = ~n42941 & ~n44019;
  assign n42359 = ~n42870 | ~n43913;
  assign n42295 = ~n42437 | ~n43876;
  assign n42433 = ~n42423 | ~n43913;
  assign n42128 = ~n42138 | ~n43748;
  assign n41186 = ~n41191 & ~n41187;
  assign n42608 = ~n42604 | ~n43748;
  assign n42878 = ~n42870 | ~n43876;
  assign n42226 = ~n42423 | ~n43876;
  assign n41669 = ~n41675 | ~n43693;
  assign n28870 = ~n42941 & ~n43794;
  assign n42447 = ~n42437 | ~n43913;
  assign n41679 = ~n41675 | ~n43523;
  assign n43550 = ~n42989 | ~n43146;
  assign n41846 = ~n41842 | ~n43523;
  assign n42897 = ~n42989 | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n42168 = ~n43031 & ~n43794;
  assign n42696 = ~n42687 | ~n32242;
  assign n42720 = ~n42716 & ~n42715;
  assign n42233 = ~n42276 | ~n43809;
  assign n42989 = ~n42708 & ~n42707;
  assign n42705 = ~n42708;
  assign n43039 = ~n43031 & ~n43729;
  assign n42379 = ~n42378 | ~n42628;
  assign n42563 = ~n42561 | ~n43748;
  assign n40806 = ~n40802 & ~n43341;
  assign n42572 = ~n42564 | ~n43876;
  assign n42625 = ~n42624 | ~n43748;
  assign n41711 = ~n41702 & ~n43755;
  assign n41269 = ~n41264 & ~n33538;
  assign n41696 = ~n41687 | ~n32242;
  assign n28839 = ~n28858 & ~n43794;
  assign n42276 = ~n42624 | ~n42232;
  assign n42126 = ~n42139 & ~n43755;
  assign n26940 = ~n41264 & ~n41754;
  assign n42378 = ~n42624 | ~n42626;
  assign n42750 = ~n42747;
  assign n27824 = ~n27822;
  assign n42051 = ~n42042 | ~n32242;
  assign n42670 = ~n42841 | ~n43876;
  assign n28060 = ~n42409 & ~n44019;
  assign n41619 = ~n41785 | ~n41616;
  assign n28075 = ~n42058 | ~n43748;
  assign n39585 = ~n39583 | ~n43525;
  assign n42415 = ~n42409 & ~n43794;
  assign n42851 = ~n42841 | ~n43913;
  assign n42624 = ~n42058 & ~n42104;
  assign n28464 = ~n28463 | ~n28462;
  assign n43527 = ~n43899 | ~n43525;
  assign n28534 = ~n28735 & ~n43794;
  assign n42058 = ~n41699 | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n42641 = ~n42632 & ~n43755;
  assign n26573 = ~n40692 & ~n43341;
  assign n41434 = ~n41425 | ~n32242;
  assign n41182 = ~n41171 | ~n43913;
  assign n42511 = ~n42505 & ~n43729;
  assign n42461 = ~n42451 | ~n43913;
  assign n41855 = ~n42505 & ~n43794;
  assign n39685 = ~n39713 | ~n43693;
  assign n41781 = ~n41772 | ~n32242;
  assign n42620 = ~n42611 & ~n43755;
  assign n42284 = ~n42281 | ~n42280;
  assign n39717 = ~n39713 | ~n43523;
  assign n40781 = ~n40942 & ~n43755;
  assign n43766 = ~n43756 & ~n43877;
  assign n42664 = ~n42203 | ~n42202;
  assign n28371 = ~n43524 | ~n41942;
  assign n27041 = ~n42505 & ~n44019;
  assign n41939 = ~n43756 & ~n41931;
  assign n25987 = ~n40784 & ~n43341;
  assign n41088 = ~n41170 & ~n43893;
  assign n28045 = ~n28044 | ~n28043;
  assign n43781 = ~n43777 & ~n43915;
  assign n40066 = ~n40067 | ~n43693;
  assign n43132 = ~n43777 | ~n43525;
  assign n41772 = ~n42173;
  assign n40497 = ~n40486 | ~n43707;
  assign n40071 = ~n40067 | ~n43523;
  assign n26557 = ~n26556 | ~n26555;
  assign n40100 = ~n40486 | ~n36906;
  assign n41048 = ~n41039 | ~n32242;
  assign n42181 = ~n42173 & ~n43794;
  assign n28225 = ~n43878 & ~n41931;
  assign n39562 = ~n39560 | ~n36906;
  assign n41488 = ~n27869 | ~n27868;
  assign n39645 = ~n39643 | ~n36906;
  assign n42095 = ~n42307 | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n38806 = n39560 & n43707;
  assign n39599 = ~n39643 | ~n43707;
  assign n41490 = ~n41079 | ~n41078;
  assign n41470 = ~n41461 | ~n32242;
  assign n41222 = ~n43611 & ~n41931;
  assign n41734 = ~n43682 | ~n41942;
  assign n27845 = ~n41953 & ~n43794;
  assign n42307 = ~n42093 | ~n42092;
  assign n26695 = ~n41953 & ~n44019;
  assign n27869 = ~n41077 | ~n41076;
  assign n41959 = ~n41953 & ~n43729;
  assign n38902 = ~n38897 & ~n33538;
  assign n41566 = ~n40053 & ~n40052;
  assign n39673 = ~n40053;
  assign n42062 = ~n27887 | ~n42090;
  assign n25798 = ~n38897 & ~n41754;
  assign n41461 = ~n41898;
  assign n27752 = ~n41399 & ~n42318;
  assign n41077 = ~n27864 | ~n27863;
  assign n41905 = ~n41898 & ~n43794;
  assign n41225 = ~n43645 & ~n41888;
  assign n40783 = ~n40941 | ~n43748;
  assign n41731 = ~n43672 & ~n41931;
  assign n43611 = ~n41211 | ~n41210;
  assign n38661 = ~n38659 | ~n36906;
  assign n27030 = ~n27029 | ~n27028;
  assign n39672 = ~n39671 & ~n39670;
  assign n40558 = ~n40549 | ~n32242;
  assign n39293 = ~n38970 & ~n39671;
  assign n38897 = ~n38969 | ~n25490;
  assign n43625 = ~n43645 & ~n43886;
  assign n43681 = ~n43672 & ~n43877;
  assign n43649 = ~n43645 & ~n43915;
  assign n39665 = ~n39664 | ~n39663;
  assign n42887 = ~n43645 | ~n43525;
  assign n41844 = ~n43317 | ~n43525;
  assign n41200 = ~n41194 & ~n43729;
  assign n43198 = ~n43317 & ~n43886;
  assign n26704 = ~n41194 & ~n43794;
  assign n40934 = ~n43196 & ~n41931;
  assign n40937 = ~n43317 & ~n41888;
  assign n26152 = ~n41194 & ~n44019;
  assign n43321 = ~n43317 & ~n43915;
  assign n41677 = ~n43582 | ~n43525;
  assign n39922 = ~n43582;
  assign n37564 = ~n37563 | ~n37562;
  assign n41613 = ~n41611 & ~n35967;
  assign n39587 = ~n39586;
  assign n26558 = ~n40152 & ~n43893;
  assign n41243 = ~n41254 | ~n41238;
  assign n41455 = ~n41454 | ~n41453;
  assign n27746 = ~n27745 | ~n27744;
  assign n43543 = ~n43582 & ~n43915;
  assign n42319 = ~n41152 | ~n41238;
  assign n39926 = ~n41657 & ~n41931;
  assign n26040 = ~n26033 & ~n44019;
  assign n39586 = ~n38798 | ~n22933;
  assign n28100 = ~n28099 & ~n28098;
  assign n39768 = ~n43224 & ~n41888;
  assign n27857 = ~n27852 | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n27856 = ~n27855 | ~n27854;
  assign n41030 = ~n41024 | ~n41453;
  assign n27745 = ~n28099 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n28762 = ~n28761 | ~n28760;
  assign n37561 = ~n37557 & ~n43811;
  assign n39921 = ~n39757 & ~n28323;
  assign n37503 = ~n37502 | ~n37501;
  assign n40070 = ~n40069 | ~n40068;
  assign n39907 = ~n41024 | ~n32242;
  assign n43586 = ~n43584 | ~n43583;
  assign n39757 = ~n40115 | ~n40114;
  assign n36908 = ~n36906 | ~n37498;
  assign n40855 = ~n40854 | ~n41147;
  assign n40716 = ~n40707 & ~n43794;
  assign n38638 = ~n39934 & ~n38636;
  assign n26090 = ~n26086 & ~n44019;
  assign n40856 = ~n40853 | ~n41149;
  assign n41151 = ~n41148 | ~n41147;
  assign n38394 = ~n38391 | ~n38390;
  assign n38266 = ~n38636 & ~n43794;
  assign n25092 = ~n38636 & ~n44019;
  assign n39689 = ~n32242 | ~n39688;
  assign n38960 = ~P2_INSTQUEUE_REG_2__3__SCAN_IN | ~n39020;
  assign n38983 = ~P2_INSTQUEUE_REG_2__4__SCAN_IN | ~n39020;
  assign n36126 = ~n36125 | ~n36124;
  assign n39023 = ~P2_INSTQUEUE_REG_2__2__SCAN_IN | ~n39020;
  assign n41148 = ~n41252 | ~n41146;
  assign n39010 = ~P2_INSTQUEUE_REG_2__6__SCAN_IN | ~n39020;
  assign n41150 = ~n41252 | ~n41149;
  assign n39002 = ~P2_INSTQUEUE_REG_2__5__SCAN_IN | ~n39020;
  assign n42725 = ~n42724 | ~n42858;
  assign n41253 = ~n41252 | ~n41251;
  assign n26389 = ~n38376 | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n41136 = ~n41130 | ~n41453;
  assign n38994 = ~P2_INSTQUEUE_REG_2__7__SCAN_IN | ~n39020;
  assign n40115 = ~n39703 & ~n28309;
  assign n40854 = ~n41252 | ~n41259;
  assign n36097 = ~n36096 | ~n36095;
  assign n37349 = ~n39934 & ~n44007;
  assign n37993 = ~n37992 | ~n37991;
  assign n39688 = ~n40493;
  assign n40494 = ~n40493 & ~n43729;
  assign n39273 = ~P2_INSTQUEUE_REG_10__4__SCAN_IN | ~n39284;
  assign n38810 = ~n38809 | ~n38808;
  assign n42294 = n42293 & n42526;
  assign n39235 = ~P2_INSTQUEUE_REG_10__2__SCAN_IN | ~n39284;
  assign n39263 = ~P2_INSTQUEUE_REG_10__7__SCAN_IN | ~n39284;
  assign n37218 = ~n44007 & ~n43794;
  assign n44012 = ~n44007 & ~n44019;
  assign n39288 = ~P2_INSTQUEUE_REG_10__3__SCAN_IN | ~n39284;
  assign n26079 = ~n40493 & ~n43794;
  assign n39020 = ~n38242 | ~n39531;
  assign n39246 = ~P2_INSTQUEUE_REG_10__0__SCAN_IN | ~n39284;
  assign n39202 = ~P2_INSTQUEUE_REG_10__6__SCAN_IN | ~n39284;
  assign n39703 = ~n37460 | ~n37459;
  assign n39255 = ~P2_INSTQUEUE_REG_10__1__SCAN_IN | ~n39284;
  assign n40064 = ~n40054 & ~n43695;
  assign n39176 = ~n40908 & ~n39191;
  assign n37878 = ~P2_INSTQUEUE_REG_8__1__SCAN_IN | ~n38217;
  assign n39142 = ~n41317 & ~n39191;
  assign n37894 = ~P2_INSTQUEUE_REG_8__6__SCAN_IN | ~n38217;
  assign n41076 = ~n27865 ^ P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n36122 = ~n43341 & ~n36121;
  assign n37886 = ~P2_INSTQUEUE_REG_8__0__SCAN_IN | ~n38217;
  assign n37460 = ~n37265 & ~n37264;
  assign n39150 = ~n39540 & ~n39191;
  assign n27861 = ~n40757 | ~n28062;
  assign n38577 = ~n40882 & ~n39603;
  assign n38898 = ~n42871;
  assign n38585 = ~n41317 & ~n39603;
  assign n39168 = ~n40896 & ~n39191;
  assign n39596 = ~n39595 | ~n39594;
  assign n27741 = ~n27740 | ~n40751;
  assign n42876 = ~n42871 & ~n43886;
  assign n36861 = ~n36860 | ~n36859;
  assign n38907 = ~n38906 | ~n41149;
  assign n39197 = ~n41289 & ~n39191;
  assign n37925 = ~P2_INSTQUEUE_REG_8__5__SCAN_IN | ~n38217;
  assign n38794 = ~n38793 | ~n38792;
  assign n38372 = ~n36857 | ~n26484;
  assign n38205 = ~P2_INSTQUEUE_REG_8__7__SCAN_IN | ~n38217;
  assign n39184 = ~n41301 & ~n39191;
  assign n38808 = ~n38807 | ~n43367;
  assign n38218 = ~P2_INSTQUEUE_REG_8__4__SCAN_IN | ~n38217;
  assign n38569 = ~n39515 & ~n39603;
  assign n38197 = ~P2_INSTQUEUE_REG_8__3__SCAN_IN | ~n38217;
  assign n37862 = ~P2_INSTQUEUE_REG_8__2__SCAN_IN | ~n38217;
  assign n39284 = ~n38301 | ~n39531;
  assign n39134 = ~n39191 & ~n39515;
  assign n37245 = ~n37242 & ~n43794;
  assign n27868 = ~n27867 | ~n27866;
  assign n38906 = ~n38905 | ~n38904;
  assign n26340 = ~n36860 | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n36859 = ~n26339 | ~n26338;
  assign n38217 = ~n37861 | ~n39531;
  assign n27865 = ~n27867 | ~n43835;
  assign n37630 = ~n37836 & ~n37629;
  assign n37265 = ~n37726 | ~n37725;
  assign n36857 = ~n26483 | ~n26482;
  assign n36487 = ~n36488;
  assign n36092 = ~n36090 | ~n36089;
  assign n41309 = ~n40891;
  assign n42640 = ~n42639 | ~n42638;
  assign n37848 = ~n39934 & ~n37846;
  assign n36860 = ~n26336 | ~n26337;
  assign n43443 = ~n43442 & ~n43441;
  assign n42875 = ~n42874 | ~n42873;
  assign n37726 = ~n36396 & ~n28282;
  assign n36396 = ~n37831 | ~n37830;
  assign n37206 = ~n37146 | ~n37145;
  assign n40891 = ~n39533 & ~n39532;
  assign n38938 = ~n38620 | ~n39531;
  assign n39364 = ~n39362 & ~n39361;
  assign n40258 = ~n40257 | ~n41257;
  assign n39096 = ~n39094 & ~n39093;
  assign n37597 = ~n36568 & ~n36567;
  assign n39332 = ~n39330 & ~n39329;
  assign n39109 = ~n39106 & ~n39105;
  assign n38856 = ~n38855 | ~n38854;
  assign n37604 = ~n36576 | ~n36575;
  assign n39965 = ~n39964 | ~n39963;
  assign n38864 = ~n38863 | ~n38862;
  assign n38872 = ~n38871 | ~n38870;
  assign n39340 = ~n39338 & ~n39337;
  assign n37621 = ~n37608 | ~n39508;
  assign n38848 = ~n38847 | ~n38846;
  assign n43837 = ~n43836 | ~n43835;
  assign n37214 = ~n37500 & ~n37499;
  assign n38840 = ~n38839 | ~n38838;
  assign n39348 = ~n39346 & ~n39345;
  assign n38880 = ~n38879 | ~n38878;
  assign n38152 = ~n41531 & ~n39796;
  assign n38892 = ~n38891 | ~n38890;
  assign n39874 = ~n39873 | ~n39872;
  assign n39072 = ~n39070 & ~n39069;
  assign n39080 = ~n39078 & ~n39077;
  assign n37416 = ~n37037 & ~n37036;
  assign n39532 = ~n39531 | ~n39530;
  assign n39866 = ~n39865 | ~n39864;
  assign n26332 = ~n36486 & ~n36485;
  assign n40046 = ~n40045 | ~n40044;
  assign n39998 = ~n39997 | ~n39996;
  assign n39088 = ~n39086 & ~n39085;
  assign n39834 = ~n39833 | ~n39832;
  assign n39324 = ~n39322 & ~n39321;
  assign n39048 = ~n39046 & ~n39045;
  assign n40009 = ~n40008 | ~n40007;
  assign n39385 = ~n39382 & ~n39381;
  assign n40020 = ~n40019 | ~n40018;
  assign n39987 = ~n39986 | ~n39985;
  assign n39826 = ~n39825 | ~n39824;
  assign n39886 = ~n39885 | ~n39884;
  assign n39858 = ~n39857 | ~n39856;
  assign n37547 = ~n36739 | ~n36738;
  assign n39976 = ~n39975 | ~n39974;
  assign n39850 = ~n39849 | ~n39848;
  assign n39356 = ~n39354 & ~n39353;
  assign n39064 = ~n39062 & ~n39061;
  assign n39372 = ~n39370 & ~n39369;
  assign n39056 = ~n39054 & ~n39053;
  assign n40031 = ~n40030 | ~n40029;
  assign n39842 = ~n39841 | ~n39840;
  assign n38102 = ~n38101 | ~n38100;
  assign n38524 = ~n38523 | ~n38522;
  assign n38432 = ~n38431 | ~n38430;
  assign n38532 = ~n38531 | ~n38530;
  assign n42983 = ~n42981 & ~n42980;
  assign n37539 = ~n36749 & ~n36748;
  assign n38540 = ~n38539 | ~n38538;
  assign n38130 = ~n38129 | ~n38128;
  assign n38416 = ~n38415 | ~n38414;
  assign n38508 = ~n38507 | ~n38506;
  assign n38118 = ~n38117 | ~n38116;
  assign n28223 = ~n43832 & ~n39482;
  assign n38456 = ~n38455 | ~n38454;
  assign n38548 = ~n38547 | ~n38546;
  assign n41316 = ~n39514 & ~n39513;
  assign n38078 = ~n38077 | ~n38076;
  assign n38516 = ~n38515 | ~n38514;
  assign n38086 = ~n38085 | ~n38084;
  assign n38560 = ~n38559 | ~n38558;
  assign n38094 = ~n38093 | ~n38092;
  assign n42492 = ~n43344 | ~n42491;
  assign n38500 = ~n38499 | ~n38498;
  assign n39345 = ~n39344 | ~n39343;
  assign n39069 = ~n39068 | ~n39067;
  assign n39361 = ~n39360 | ~n39359;
  assign n38448 = ~n38447 | ~n38446;
  assign n39077 = ~n39076 | ~n39075;
  assign n39321 = ~n39320 | ~n39319;
  assign n39085 = ~n39084 | ~n39083;
  assign n39329 = ~n39328 | ~n39327;
  assign n39045 = ~n39044 | ~n39043;
  assign n39337 = ~n39336 | ~n39335;
  assign n38440 = ~n38439 | ~n38438;
  assign n39381 = ~n39380 | ~n39379;
  assign n28872 = ~n43803 | ~n42491;
  assign n38476 = ~n38475 | ~n38474;
  assign n36373 = ~n36375 | ~n36374;
  assign n39353 = ~n39352 | ~n39351;
  assign n39061 = ~n39060 | ~n39059;
  assign n39105 = ~n39104 | ~n39103;
  assign n38424 = ~n38423 | ~n38422;
  assign n37934 = ~n37657 & ~n37656;
  assign n28725 = ~n42491 | ~n44021;
  assign n39369 = ~n39368 | ~n39367;
  assign n38070 = ~n38069 | ~n38068;
  assign n39093 = ~n39092 | ~n39091;
  assign n36801 = ~n36656 | ~n39531;
  assign n39053 = ~n39052 | ~n39051;
  assign n38110 = ~n38109 | ~n38108;
  assign n37356 = ~n36553 | ~n36552;
  assign n37372 = ~n39524 & ~n37365;
  assign n38464 = ~n38463 | ~n38462;
  assign n28894 = ~n43803 | ~n42551;
  assign n41876 = ~n41872 | ~n41871;
  assign n38625 = ~n39508 | ~n38616;
  assign n27858 = ~n26430 & ~n26429;
  assign n39286 = ~n38280;
  assign n42981 = ~n40077 & ~n40073;
  assign n42552 = ~n43344 | ~n42551;
  assign n28827 = ~n42551 | ~n44021;
  assign n37038 = ~n39508 | ~n37033;
  assign n37767 = ~n40239 | ~n40857;
  assign n37143 = ~n39508 | ~n37135;
  assign n40256 = ~n40239 | ~n40980;
  assign n43828 = ~n43753 | ~n43835;
  assign n43832 = ~n41872 ^ n28209;
  assign n36553 = ~n36206 & ~n36205;
  assign n43195 = ~n43659 | ~n43835;
  assign n28673 = ~n43376 | ~n44021;
  assign n38280 = ~n37045 | ~n37947;
  assign n41872 = ~n41933 & ~n41932;
  assign n37364 = ~n38773 & ~n39543;
  assign n36745 = ~n39508 | ~n36736;
  assign n38556 = ~n39818 | ~n38497;
  assign n42006 = ~n43344 | ~n43376;
  assign n44013 = ~n24869 | ~n34815;
  assign n38319 = ~n37147 & ~n37947;
  assign n38612 = ~n38615 | ~n37947;
  assign n43382 = ~n43803 | ~n43376;
  assign n37651 = ~n39508 | ~n37642;
  assign n38615 = ~n37946 & ~n37945;
  assign n39509 = n39508 & n39507;
  assign n37025 = ~n39445 | ~n40857;
  assign n41554 = ~n42338 | ~n41553;
  assign n39446 = ~n39445 | ~n40980;
  assign n26427 = ~n26411 | ~n26410;
  assign n36253 = ~n36248 | ~n25113;
  assign n44098 = ~n34521 | ~n34520;
  assign n28722 = ~n28721 & ~n28720;
  assign n38127 = ~n38067 | ~n38066;
  assign n36653 = ~n36652 & ~n38321;
  assign n39607 = n37650 & n37947;
  assign n26426 = ~n26425 | ~n26424;
  assign n39411 = ~n39410 | ~n40980;
  assign n26582 = ~n26581 | ~P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n37570 = ~n38147 & ~n38143;
  assign n37627 = ~n37626 | ~n39531;
  assign n24722 = ~n24720 | ~n24719;
  assign n41875 = ~n41874 | ~n41873;
  assign n26411 = ~n26404 & ~n26403;
  assign n28841 = ~n43803 | ~n42934;
  assign n37946 = ~n23700 | ~n37638;
  assign n43193 = ~n43192 | ~n43835;
  assign n42645 = ~n42934 | ~n44021;
  assign n42936 = ~n43344 | ~n42934;
  assign n37650 = ~n23700 & ~n37639;
  assign n37367 = ~n38334 & ~n37361;
  assign n42908 = ~n43209 | ~n43207;
  assign n43183 = ~n43209;
  assign n38473 = ~n38413 | ~n38412;
  assign n39507 = ~n23700 | ~n37363;
  assign n43176 = ~n43530 | ~n43549;
  assign n43184 = ~n43530;
  assign n26410 = ~n26409 & ~n26408;
  assign n28473 = ~n43343 | ~n44021;
  assign n34599 = ~n34094 | ~n34093;
  assign n26425 = ~n26417 & ~n26416;
  assign n43192 = n40926 ^ n40925;
  assign n26424 = ~n26423 & ~n26422;
  assign n43174 = ~n43207;
  assign n40977 = ~n40976 | ~n41257;
  assign n39410 = ~n36886 | ~n37569;
  assign n26352 = ~n26350 | ~n26349;
  assign n26404 = ~n26402 | ~n26401;
  assign n43347 = ~n43344 | ~n43343;
  assign n43027 = ~n28853;
  assign n35096 = ~n35185 | ~n35037;
  assign n34513 = ~n35627 | ~n44102;
  assign n41395 = ~n41394 | ~n41683;
  assign n40347 = ~n40345 & ~n42336;
  assign n34363 = ~n34131 | ~n34130;
  assign n41394 = ~n41392 | ~n41391;
  assign n38298 = ~n38297 | ~n39524;
  assign n35330 = ~n35332;
  assign n26323 = ~n26322 | ~n26321;
  assign n39119 = ~n39118 & ~n39511;
  assign n25933 = ~n26569 | ~n25932;
  assign n25968 = ~n43462 | ~n25967;
  assign n43171 = n39928 ^ n39927;
  assign n37644 = ~n37641 & ~n39508;
  assign n28536 = ~n43803 | ~n42833;
  assign n24670 = ~n24669;
  assign n24620 = ~n35332 & ~n35366;
  assign n25971 = ~n43462 | ~n38642;
  assign n39127 = ~n39126 | ~n39524;
  assign n35244 = ~n35185 | ~n35184;
  assign n34584 = ~n37486 | ~n33733;
  assign n26564 = ~n43462 | ~n25981;
  assign n42835 = ~n43344 | ~n42833;
  assign n26350 = ~n26344 & ~n26343;
  assign n34752 = ~n35185 | ~n34425;
  assign n28728 = ~n43462 | ~n42367;
  assign n26358 = ~n26356 | ~n26355;
  assign n26368 = ~n26367 | ~n26366;
  assign n40148 = ~n42336 & ~n40147;
  assign n27825 = ~n43462 | ~n40798;
  assign n25977 = ~n43462 | ~n40091;
  assign n42417 = ~n43803 | ~n42408;
  assign n38385 = ~n43462 & ~n38643;
  assign n41684 = ~n41681 | ~n41683;
  assign n42373 = ~n43344 | ~n42408;
  assign n24858 = ~n24851 & ~n24873;
  assign n38619 = ~n38614 & ~n39508;
  assign n42003 = ~n22933 & ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n42901 = ~n42997 | ~n42996;
  assign n33793 = ~n24840 & ~n24839;
  assign n43448 = ~n22933 & ~P1_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n28729 = ~n22933 | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n40851 = ~n40850 | ~n41259;
  assign n34425 = ~n34424 & ~n34423;
  assign n24851 = ~n24716 | ~n25897;
  assign n28476 = ~n22933 | ~P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n27722 = ~n27721 | ~n41149;
  assign n26251 = ~n26250 | ~n26249;
  assign n26355 = ~n37870 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n24737 = ~n24859 & ~n24745;
  assign n41381 = ~n41380 | ~n41670;
  assign n25979 = ~n22933 | ~P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n41386 = ~n41385 | ~n41670;
  assign n42500 = ~n22933 | ~n42579;
  assign n38383 = ~n22933 | ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n24860 = ~n24859 & ~n24873;
  assign n40813 = ~n40812 | ~n41390;
  assign n38239 = ~n38238 | ~n39524;
  assign n25972 = ~n22933 & ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n26407 = ~n38329 | ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n25970 = ~n22933 | ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n35014 = ~n34269 | ~n34268;
  assign n41769 = ~n42172 | ~n44021;
  assign n22933 = n25897 & n24746;
  assign n38238 = ~n38237 | ~n39522;
  assign n42183 = ~n43803 | ~n42172;
  assign n26233 = ~n26364 & ~n26232;
  assign n26245 = ~n26240 | ~n26239;
  assign n27718 = ~n27720 | ~n27717;
  assign n41907 = ~n43803 | ~n42586;
  assign n37376 = ~n26370;
  assign n40234 = ~n42336 & ~n40232;
  assign n40528 = ~n40527 & ~n40526;
  assign n25931 = ~n25897 | ~n25896;
  assign n41441 = ~n42586 | ~n44021;
  assign n37639 = ~n37638 | ~n37637;
  assign n28553 = ~n43344 | ~n42172;
  assign n40479 = ~n40478 & ~n40527;
  assign n37363 = ~n37638 & ~n37945;
  assign n28056 = n28055 & n28054;
  assign n28092 = ~n41114 | ~n41542;
  assign n41008 = ~n41007 | ~n41006;
  assign n41010 = ~n41003 | ~n41002;
  assign n42904 = ~n40121 ^ n40120;
  assign n42588 = ~n43344 | ~n42586;
  assign n33918 = ~n35262 | ~n35261;
  assign n27721 = ~n27720 | ~P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n40401 = ~n40400 & ~n40527;
  assign n41063 = ~P3_EBX_REG_26__SCAN_IN & ~n41390;
  assign n40812 = ~n40811 | ~n40810;
  assign n37130 = ~n37638 & ~n37637;
  assign n41670 = ~n41379 | ~n41378;
  assign n41515 = ~n41514 | ~n41513;
  assign n40547 = ~n40546 | ~n40810;
  assign n41115 = ~n41397 & ~n41114;
  assign n36648 = ~n26361;
  assign n40517 = ~n42336 & ~n40516;
  assign n40850 = ~n41514 | ~P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n35354 = ~n35185 | ~n34730;
  assign n41003 = ~n41001 | ~n41229;
  assign n39745 = ~n39744 | ~n40545;
  assign n39447 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN | ~n39444;
  assign n41514 = ~n40847 & ~n41233;
  assign n40746 = ~n41541 | ~n40743;
  assign n26310 = ~n38628 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n42682 = ~n43344 | ~n42680;
  assign n26312 = ~n37039 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n42899 = n39710 ^ n39709;
  assign n41543 = n41542 & n41541;
  assign n24710 = ~n24715 | ~n24712;
  assign n24828 = ~n24615 | ~n24623;
  assign n26240 = ~n37039 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n27719 = ~n37710 | ~n27715;
  assign n41857 = ~n43803 | ~n42680;
  assign n24841 = ~n24715 ^ n24712;
  assign n35623 = ~n33731 | ~n33730;
  assign n35262 = ~n27894 & ~n27893;
  assign n39505 = ~n39504 | ~n39741;
  assign n27847 = ~n43803 | ~n41969;
  assign n40462 = ~n42336 & ~n40460;
  assign n27894 = ~n36258 | ~n36257;
  assign n41439 = ~n41435;
  assign n40847 = ~n40748 | ~n40747;
  assign n40476 = ~n40475 | ~n40474;
  assign n42882 = ~n42868 | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n42711 = ~n42466 & ~n42353;
  assign n32895 = ~n32894 | ~n32893;
  assign n32800 = ~n32347 | ~n32263;
  assign n24496 = ~n24495;
  assign n40747 = ~n40998 & ~n39437;
  assign n36258 = ~n35250 & ~n35249;
  assign n42351 = ~n42352 | ~n43835;
  assign n27349 = ~n42321 & ~n38924;
  assign n42024 = ~n41373 | ~n41372;
  assign n24609 = ~n24614 | ~n24610;
  assign n41438 = ~n41437 & ~n41436;
  assign n38153 = ~n39437 & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n32347 = ~n32264;
  assign n40245 = ~n41235 & ~n40244;
  assign n32264 = ~n32345 | ~n32344;
  assign n39771 = ~n39450 | ~n40341;
  assign n41745 = ~n43344 | ~n41743;
  assign n27844 = ~n27843 | ~n27842;
  assign n40405 = ~n40381 & ~n42336;
  assign n26691 = n26690 & n26689;
  assign n39437 = ~n39775 | ~n38142;
  assign n39789 = ~n39788 | ~n39787;
  assign n39393 = ~n39391 & ~n40341;
  assign n26706 = ~n43803 | ~n41276;
  assign n26703 = ~n26702 | ~n43033;
  assign n32891 = ~n23697 ^ n23695;
  assign n41456 = ~n43803 | ~n41743;
  assign n35250 = ~n26521 | ~n26520;
  assign n23698 = ~n23697 | ~n23696;
  assign n42414 = ~n42413 | ~n42412;
  assign n37772 = ~n40244 & ~n41397;
  assign n40745 = ~n41545 | ~n40744;
  assign n37509 = ~n37226 & ~n43566;
  assign n26521 = ~n26516 | ~n26515;
  assign n26520 = ~n26519 | ~n26518;
  assign n40985 = ~n40984 | ~n40983;
  assign n42700 = ~n42111 | ~n42110;
  assign n36143 = ~n35467 & ~n41453;
  assign n37919 = ~n37921;
  assign n32545 = ~n24494 | ~n24493;
  assign n41276 = ~n26148 & ~n26715;
  assign n41113 = ~n41545 & ~n41516;
  assign n40341 = ~n39390 | ~n39389;
  assign n41547 = ~n41546 | ~n41545;
  assign n40411 = ~n39395 | ~n40470;
  assign n41545 = ~n27749 | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n27707 = ~n36192 | ~n27704;
  assign n42199 = ~n42246;
  assign n26516 = ~n26517 | ~n26514;
  assign n41034 = ~n43803 | ~n41022;
  assign n32629 = n31796 & n31795;
  assign n42247 = ~n42245 | ~n42244;
  assign n39636 = ~n39635 & ~n42336;
  assign n42243 = n40630 ^ n40629;
  assign n43583 = ~n43877;
  assign n23694 = ~n32143 | ~n32144;
  assign n34575 = ~n34124 & ~n39944;
  assign n40706 = ~n25945 & ~n26142;
  assign n42237 = ~n42236 & ~n42235;
  assign n35173 = ~n34124 | ~n34551;
  assign n40278 = ~n40277 & ~n42336;
  assign n36169 = ~n36168 | ~n36167;
  assign n43794 = ~n41894 | ~n26062;
  assign n28370 = ~n28369 & ~n28368;
  assign n40630 = ~n40587 & ~n40586;
  assign n28213 = ~n37288 | ~n28212;
  assign n28210 = ~P2_EBX_REG_31__SCAN_IN | ~n37288;
  assign n38923 = ~n40242 | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n24781 = ~n23690;
  assign n34279 = n42922 & n43331;
  assign n41979 = ~n42922 | ~n34287;
  assign n43893 = ~n26550 | ~n26431;
  assign n25670 = ~n36829 | ~n36828;
  assign n40960 = ~n40376 & ~n40375;
  assign n41308 = ~n39271;
  assign n40895 = ~n39285;
  assign n37774 = ~n40242 & ~n41408;
  assign n40185 = ~n40182 | ~n40181;
  assign n35546 = ~n35545 | ~n35544;
  assign n40204 = ~n40200 | ~n40199;
  assign n42110 = ~n26215 | ~n28156;
  assign n41206 = ~n41919;
  assign n39948 = ~n39959 | ~n39942;
  assign n38696 = ~n36694 | ~n36693;
  assign n43735 = ~n43734 & ~P1_EAX_REG_31__SCAN_IN;
  assign n39811 = ~n39821 | ~n39942;
  assign n38715 = ~n36560 | ~n36559;
  assign n43738 = n43734 & n39902;
  assign n43737 = n43734 & n39897;
  assign n43306 = n43734 & n39893;
  assign n40376 = ~n40371 & ~n41235;
  assign n38706 = ~n36621 | ~n36620;
  assign n36193 = ~n27709 | ~n41149;
  assign n43441 = ~n43344;
  assign n36692 = ~n36802 | ~BUF2_REG_30__SCAN_IN;
  assign n40911 = ~n36561 & ~n36794;
  assign n24132 = ~n24205;
  assign n43689 = ~n25102 & ~n36557;
  assign n23689 = ~n35790 | ~n31816;
  assign n36694 = ~n36802 | ~BUF2_REG_22__SCAN_IN;
  assign n36693 = ~n36803 | ~BUF1_REG_22__SCAN_IN;
  assign n36591 = ~n36803 | ~BUF1_REG_31__SCAN_IN;
  assign n36587 = ~n36802 | ~BUF2_REG_23__SCAN_IN;
  assign n36560 = ~n36802 | ~BUF2_REG_18__SCAN_IN;
  assign n36592 = ~n36802 | ~BUF2_REG_31__SCAN_IN;
  assign n36691 = ~n36803 | ~BUF1_REG_30__SCAN_IN;
  assign n32107 = ~n32237;
  assign n36633 = ~BUF2_REG_24__SCAN_IN | ~n36802;
  assign n34687 = ~n35185;
  assign n36632 = ~BUF1_REG_24__SCAN_IN | ~n36803;
  assign n39516 = ~n37289 & ~n36794;
  assign n36559 = ~n36803 | ~BUF1_REG_18__SCAN_IN;
  assign n36642 = ~BUF2_REG_16__SCAN_IN | ~n36802;
  assign n25625 = ~n36831 | ~n36830;
  assign n36682 = ~n36803 | ~BUF1_REG_21__SCAN_IN;
  assign n36624 = ~n36803 | ~BUF1_REG_25__SCAN_IN;
  assign n35381 = ~n41754 | ~n43695;
  assign n36683 = ~n36802 | ~BUF2_REG_21__SCAN_IN;
  assign n36643 = ~BUF1_REG_16__SCAN_IN | ~n36803;
  assign n36586 = ~n36803 | ~BUF1_REG_23__SCAN_IN;
  assign n40668 = ~n44002 | ~n40350;
  assign n36799 = ~n36803 | ~BUF1_REG_27__SCAN_IN;
  assign n36800 = ~n36802 | ~BUF2_REG_27__SCAN_IN;
  assign n40838 = ~n40837 | ~n40836;
  assign n36805 = ~n36802 | ~BUF2_REG_19__SCAN_IN;
  assign n36621 = ~n36802 | ~BUF2_REG_17__SCAN_IN;
  assign n36784 = ~n36803 | ~BUF1_REG_20__SCAN_IN;
  assign n37488 = ~n37476 & ~n39942;
  assign n36785 = ~n36802 | ~BUF2_REG_20__SCAN_IN;
  assign n36804 = ~n36803 | ~BUF1_REG_19__SCAN_IN;
  assign n36620 = ~n36803 | ~BUF1_REG_17__SCAN_IN;
  assign n43547 = ~n43911 & ~n43546;
  assign n41340 = ~n41353;
  assign n41355 = ~n41354 | ~n41353;
  assign n36677 = ~n36802 | ~BUF2_REG_29__SCAN_IN;
  assign n36676 = ~n36803 | ~BUF1_REG_29__SCAN_IN;
  assign n40676 = ~n40607 & ~n40606;
  assign n36783 = ~n36802 | ~BUF2_REG_28__SCAN_IN;
  assign n43734 = ~n32237 | ~n32236;
  assign n39821 = ~n37476;
  assign n36782 = ~n36803 | ~BUF1_REG_28__SCAN_IN;
  assign n43297 = ~n44019;
  assign n36578 = ~n36803 | ~BUF1_REG_26__SCAN_IN;
  assign n39818 = ~n37486 & ~n39956;
  assign n42089 = ~n42066 & ~n42353;
  assign n26069 = ~n26068 | ~n35473;
  assign n26056 = ~P1_EBX_REG_31__SCAN_IN | ~n35473;
  assign n36002 = ~n41759 | ~n32218;
  assign n40017 = ~n37486 & ~n34074;
  assign n40028 = ~n37486 & ~n34151;
  assign n40043 = ~n37486 & ~n34606;
  assign n39984 = ~n37486 & ~n34136;
  assign n39995 = ~n37486 & ~n34166;
  assign n40006 = ~n37486 & ~n34228;
  assign n39973 = ~n37486 & ~n34189;
  assign n39962 = ~n37486 & ~n34243;
  assign n36162 = ~n41401 | ~n35940;
  assign n35766 = n23538 & n23537;
  assign n32237 = ~n31722 | ~n31721;
  assign n43713 = ~n40693 | ~n26591;
  assign n24205 = ~n24129 | ~n44102;
  assign n40503 = ~n40372 | ~n36447;
  assign n23617 = ~n26235 & ~n23676;
  assign n39953 = ~n38058 | ~n38057;
  assign n34165 = ~n34241 & ~n34164;
  assign n35473 = ~n26047 | ~n31273;
  assign n34242 = ~n34241 & ~n22947;
  assign n42081 = ~n40282 | ~n43835;
  assign n25587 = ~n25584 | ~n25583;
  assign n34188 = ~n34241 & ~n34187;
  assign n25584 = ~n34903 | ~n34902;
  assign n41495 = ~n39461 & ~n42353;
  assign n41301 = ~n40056 | ~n39531;
  assign n34914 = ~n39531 & ~n32074;
  assign n43811 = ~n43913;
  assign n43924 = ~n27923 | ~n43061;
  assign n26497 = ~n26496 & ~n42353;
  assign n40908 = ~n38018 | ~n39531;
  assign n40896 = ~n36792 | ~n39531;
  assign n27348 = ~n27343 & ~n27344;
  assign n40167 = ~n38595 | ~n38594;
  assign n24486 = ~n24485;
  assign n24813 = ~n24812 & ~n43294;
  assign n34241 = ~n34071 | ~n34070;
  assign n43295 = ~n43558 | ~n43294;
  assign n31439 = n44028 & n31382;
  assign n41289 = ~n36590 | ~n39531;
  assign n39540 = ~n37434 | ~n39531;
  assign n40882 = ~n39675 | ~n39531;
  assign n32236 = ~n32235 | ~n44102;
  assign n39515 = ~n37112 | ~n39531;
  assign n26203 = ~n26185 & ~n26184;
  assign n41317 = ~n38972 | ~n39531;
  assign n24128 = ~n24107 | ~n24106;
  assign n32235 = ~n32234 | ~n32233;
  assign n26185 = ~n26183 & ~n26182;
  assign n28773 = ~n28716 & ~n28715;
  assign n34119 = ~n34551;
  assign n34355 = ~P3_EAX_REG_10__SCAN_IN | ~n34966;
  assign n37830 = ~n28275 | ~n28274;
  assign n28817 = ~n43138 | ~n43294;
  assign n34903 = n25583 ^ n25578;
  assign n37355 = ~n28268 | ~n28267;
  assign n41491 = ~n38945 | ~n43835;
  assign n36158 = ~P3_REIP_REG_28__SCAN_IN | ~n35640;
  assign n24765 = ~P2_PHYADDRPOINTER_REG_30__SCAN_IN | ~n28147;
  assign n37725 = ~n28288 | ~n28287;
  assign n40114 = ~n28315 | ~n28314;
  assign n36552 = ~n28261 | ~n28260;
  assign n26061 = ~n43293 | ~P1_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n36063 = ~n36061;
  assign n23667 = ~n23642 | ~n23641;
  assign n39702 = ~n28308 | ~n28307;
  assign n31905 = ~n31904 | ~n31903;
  assign n37459 = ~n28301 | ~n28300;
  assign n36395 = ~n28281 | ~n28280;
  assign n24127 = ~n24126 & ~n31894;
  assign n35695 = n34967 & n34966;
  assign n35534 = ~n41401 | ~n35532;
  assign n39404 = ~n42322 & ~n36509;
  assign n36901 = ~n35821 | ~n25076;
  assign n26183 = ~n28150 & ~n37289;
  assign n23644 = n26515 ^ n26518;
  assign n24445 = ~n24442;
  assign n36061 = ~n32377 | ~n32376;
  assign n36429 = ~n27688 | ~n27687;
  assign n36039 = ~n36038 & ~n36041;
  assign n23516 = ~n31779 | ~n31768;
  assign n24096 = ~n31927 | ~n24095;
  assign n24126 = ~n31927 & ~n24108;
  assign n28274 = ~n39578 | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n28234 = ~n39578 | ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n28233 = ~n28361 & ~n28229;
  assign n28273 = ~n28361 & ~n29506;
  assign n28246 = ~n28361 & ~n29221;
  assign n27632 = ~n41539 | ~n40968;
  assign n35541 = ~n34628 | ~n34659;
  assign n28247 = ~n39578 | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n26182 = ~n31524 & ~n23127;
  assign n28254 = ~n39578 | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n28253 = ~n28361 & ~n28249;
  assign n28294 = ~n39578 | ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n27898 = ~n28361 & ~n29199;
  assign n27899 = ~n39578 | ~P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n26528 = ~n39578 | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n28145 = ~P2_PHYADDRPOINTER_REG_28__SCAN_IN | ~n28107;
  assign n28240 = ~n28361 & ~n28236;
  assign n26535 = ~n39578 | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n28241 = ~n39578 | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n26534 = ~n28361 & ~n26530;
  assign n31912 = ~n31909 & ~n31908;
  assign n41540 = ~n40968;
  assign n27919 = ~n28361 & ~n27915;
  assign n27920 = ~n39578 | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n26495 = ~n27879;
  assign n36042 = ~n36041 | ~n40968;
  assign n26541 = ~n28361 & ~n26537;
  assign n28260 = ~n39578 | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n26542 = ~n39578 | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n28259 = ~n28361 & ~n29471;
  assign n28280 = ~n39578 | ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n28655 = ~n43378 | ~n43294;
  assign n28287 = ~n39578 | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n27905 = ~n28361 & ~n27901;
  assign n27911 = ~n28361 & ~n29204;
  assign n28267 = ~n39578 | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n26526 = ~n28361 & ~n26522;
  assign n39958 = n39942 & n39315;
  assign n25574 = ~n32890 & ~n32889;
  assign n26515 = ~n23629 & ~n23628;
  assign n24442 = ~n24434 & ~n24433;
  assign n42339 = ~n42338 & ~n42337;
  assign n24808 = ~n34552 | ~n25932;
  assign n27341 = ~n36022 & ~n40196;
  assign n27687 = ~n27686 | ~n27685;
  assign n41016 = ~n42338 & ~n41002;
  assign n40843 = ~n42338 & ~n42321;
  assign n36282 = ~n36239;
  assign n35823 = ~n34818 | ~n34817;
  assign n40529 = ~n42338;
  assign n34641 = ~n41401 | ~n34673;
  assign n26494 = ~n26493 & ~n26492;
  assign n33772 = ~n33923;
  assign n24433 = ~n24432 & ~n24431;
  assign n40968 = ~n32361 | ~n27631;
  assign n31524 = ~n23288 | ~n23287;
  assign n31909 = ~n23949 | ~n23948;
  assign n23635 = ~n23591;
  assign n32147 = ~n23722 & ~n23415;
  assign n25566 = ~n25565 | ~n25564;
  assign n34843 = ~n32206 | ~n32807;
  assign n31765 = ~n26199 & ~n26198;
  assign n32608 = ~n36242 | ~n43957;
  assign n28460 = ~n43035 | ~n43294;
  assign n42338 = ~n42336 | ~n40865;
  assign n36021 = ~n27340 & ~n27339;
  assign n28153 = ~n28152 | ~n31525;
  assign n32566 = ~n32485 | ~n36242;
  assign n31286 = ~n31202 | ~n23127;
  assign n41371 = ~n41331;
  assign n32606 = ~n33090 & ~n32488;
  assign n32807 = ~n33090;
  assign n34611 = ~n32866 & ~n32849;
  assign n35609 = ~n41537 & ~n35608;
  assign n25572 = ~n25562 | ~n25563;
  assign n41331 = ~n32373 | ~n32372;
  assign n25565 = ~n25562;
  assign n26484 = ~n40570 | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n36359 = n36358 & n36357;
  assign n27682 = ~n36020 | ~n36019;
  assign n23674 = ~n23612 & ~n23611;
  assign n32678 = ~n32672 | ~n32671;
  assign n26207 = ~n23717 & ~n23716;
  assign n26488 = ~n26478 | ~n26477;
  assign n28346 = ~n23571 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n28511 = ~n27974 & ~n27973;
  assign n28037 = ~n43294 | ~n42410;
  assign n23632 = ~n23630 & ~n35715;
  assign n28142 = ~P2_PHYADDRPOINTER_REG_24__SCAN_IN | ~n28109;
  assign n25562 = ~n25555 | ~n25554;
  assign n27620 = ~n27617 | ~n27793;
  assign n23935 = ~n23928 & ~n23927;
  assign n23264 = ~n23263 | ~n23564;
  assign n32201 = ~n41374 & ~n32368;
  assign n32370 = ~n32369 | ~n32368;
  assign n25555 = ~n32168 | ~n32167;
  assign n31771 = ~n26508 | ~n32509;
  assign n27817 = ~n27816 | ~n27815;
  assign n31954 = ~n31953 & ~n32526;
  assign n26197 = ~n26196 | ~n26445;
  assign n23927 = ~n23926 & ~n23925;
  assign n41408 = ~n40744;
  assign n23222 = ~n23219 | ~n23218;
  assign n24430 = ~n24428 & ~n33710;
  assign n24226 = ~n24215 & ~n24214;
  assign n27815 = ~n27814 & ~n27813;
  assign n32368 = ~n32200 | ~n32199;
  assign n27027 = ~n42507 | ~n43294;
  assign n32369 = ~n32367 | ~n32366;
  assign n28140 = ~P2_PHYADDRPOINTER_REG_22__SCAN_IN | ~n28110;
  assign n27335 = ~n27331 & ~n27330;
  assign n23611 = ~n23610 | ~n23609;
  assign n23560 = ~n23593 | ~n23558;
  assign n32366 = ~n31825 & ~n31824;
  assign n31768 = ~n26545 & ~n23545;
  assign n23551 = ~n23550 & ~n23549;
  assign n23552 = ~n23701 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n32197 = ~n33487 | ~n32196;
  assign n24215 = ~n24213 | ~n24212;
  assign n27873 = ~n27871 | ~n23085;
  assign n32846 = ~n32845 | ~n32844;
  assign n32167 = ~n32214 | ~n32213;
  assign n23639 = ~n23638 | ~n23637;
  assign n28149 = ~n31766 & ~n32149;
  assign n24246 = ~n24133 | ~n22947;
  assign n25064 = ~n25063 | ~n25062;
  assign n26431 = ~n31764;
  assign n32213 = ~n25552 | ~n25551;
  assign n25564 = ~n25563;
  assign n26545 = ~n23492 | ~n23491;
  assign n31659 = ~n31826 | ~n41324;
  assign n27675 = ~n36974 | ~n36973;
  assign n41402 = ~P3_PHYADDRPOINTER_REG_29__SCAN_IN | ~n35654;
  assign n26678 = ~n41955 | ~n43294;
  assign n28138 = ~P2_PHYADDRPOINTER_REG_20__SCAN_IN | ~n28111;
  assign n37123 = ~n25776 | ~n25775;
  assign n32373 = ~n27802 & ~n27801;
  assign n23546 = ~n23544 & ~n23543;
  assign n26436 = ~n26434 | ~n41873;
  assign n25715 = ~n41473 | ~P2_REIP_REG_7__SCAN_IN;
  assign n26636 = ~n41444 | ~n43294;
  assign n26091 = ~n26032 & ~n26031;
  assign n41324 = ~n33486 & ~n31532;
  assign n25629 = ~n41473 | ~P2_REIP_REG_5__SCAN_IN;
  assign n27812 = ~n29940 | ~n27811;
  assign n28111 = ~n42354 & ~n28137;
  assign n36272 = ~n24912 | ~n24911;
  assign n25591 = ~n41473 | ~P2_REIP_REG_4__SCAN_IN;
  assign n31810 = ~n31809 & ~n32371;
  assign n25674 = ~n41473 | ~P2_REIP_REG_6__SCAN_IN;
  assign n41250 = ~n41147 & ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n37213 = ~n24987 | ~n24986;
  assign n25570 = ~n41473 | ~P2_REIP_REG_2__SCAN_IN;
  assign n23657 = ~n23656 | ~n23655;
  assign n25537 = ~n25539;
  assign n32214 = ~n25546 | ~n25545;
  assign n24751 = ~n31477 | ~n24750;
  assign n37568 = ~n41147 | ~n40421;
  assign n25551 = ~n41473 | ~P2_REIP_REG_0__SCAN_IN;
  assign n35654 = ~n41092 & ~n35529;
  assign n43055 = ~n42797 | ~n42796;
  assign n24427 = ~n24426 | ~n24425;
  assign n23228 = ~n23227 | ~n23226;
  assign n25538 = ~n25536 & ~n25535;
  assign n23692 = ~n23691;
  assign n23681 = ~n23680 | ~n23679;
  assign n27700 = ~n41147 | ~n27699;
  assign n26434 = ~n23217 & ~n23216;
  assign n25721 = ~n25550 & ~n27901;
  assign n23499 = ~n23548;
  assign n27729 = ~n41149 | ~n27728;
  assign n27704 = ~n41149 | ~n27703;
  assign n25735 = ~n25550 & ~n27915;
  assign n25789 = ~n25550 & ~n29493;
  assign n25756 = ~n25550 & ~n29221;
  assign n26439 = ~n26437 | ~n41873;
  assign n23567 = ~n31058 & ~n36357;
  assign n27670 = ~n36665 | ~n36664;
  assign n26136 = ~n41196 | ~n43294;
  assign n25763 = ~n25550 & ~n28249;
  assign n32371 = ~n31808 & ~n31807;
  assign n23733 = ~n31058;
  assign n23132 = ~n23131 | ~n24775;
  assign n25743 = ~n25550 & ~n28229;
  assign n27715 = ~n41149 & ~P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n23133 = ~n26437 & ~n31498;
  assign n28137 = ~P2_PHYADDRPOINTER_REG_18__SCAN_IN | ~n28112;
  assign n38143 = ~n41149 | ~P3_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n25780 = ~n25550 & ~n29506;
  assign n26677 = ~n26676 | ~n26675;
  assign n24223 = ~n24231 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n25749 = ~n25550 & ~n28236;
  assign n26924 = ~n25550 & ~n29511;
  assign n23680 = ~n23678 | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n27695 = ~n41149 | ~n27694;
  assign n35529 = ~n40732 | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n23662 = ~n42796 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n28665 = ~n28664 | ~n28663;
  assign n25770 = ~n25550 & ~n29471;
  assign n23556 = ~n23555 | ~n23554;
  assign n23691 = ~n42796 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n25582 = ~n25550 & ~n38814;
  assign n27742 = ~n41149 & ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n23695 = ~n42796 | ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n23227 = ~n23225 | ~n23224;
  assign n42748 = ~n41829 | ~n42796;
  assign n27608 = ~n27602 | ~n27626;
  assign n25729 = ~n25550 & ~n29204;
  assign n31371 = ~n27797 | ~n27796;
  assign n25561 = ~n25556 & ~n26282;
  assign n24192 = ~n40080 | ~P1_EBX_REG_7__SCAN_IN;
  assign n31447 = ~n32082 | ~n31793;
  assign n24195 = ~n40080 | ~P1_EBX_REG_8__SCAN_IN;
  assign n24189 = ~n40080 | ~P1_EBX_REG_6__SCAN_IN;
  assign n25078 = ~n40080 | ~P1_EBX_REG_9__SCAN_IN;
  assign n25081 = ~n40080 | ~P1_EBX_REG_10__SCAN_IN;
  assign n27800 = ~n32361;
  assign n25084 = ~n40080 | ~P1_EBX_REG_11__SCAN_IN;
  assign n24186 = ~n40080 | ~P1_EBX_REG_5__SCAN_IN;
  assign n25087 = ~n40080 | ~P1_EBX_REG_12__SCAN_IN;
  assign n25843 = ~n40080 | ~P1_EBX_REG_13__SCAN_IN;
  assign n31807 = ~n29940 | ~n27597;
  assign n25938 = ~n40080 | ~P1_EBX_REG_14__SCAN_IN;
  assign n25941 = ~n40080 | ~P1_EBX_REG_15__SCAN_IN;
  assign n23548 = ~n23498 & ~n32217;
  assign n41235 = ~n41542;
  assign n24183 = ~n40080 | ~P1_EBX_REG_4__SCAN_IN;
  assign n24180 = ~n40080 | ~P1_EBX_REG_3__SCAN_IN;
  assign n25545 = ~n25557 & ~n41474;
  assign n31823 = ~n32361 & ~n33487;
  assign n24105 = ~n24104 | ~n24103;
  assign n27343 = ~n27342 | ~n39615;
  assign n27607 = ~n27606 | ~n29940;
  assign n23452 = ~n23448 | ~n23447;
  assign n26437 = ~n23126 | ~n23125;
  assign n27602 = ~n27601 | ~n29940;
  assign n23170 = ~n23558;
  assign n41149 = ~n27689 & ~n35858;
  assign n24780 = ~n24779 & ~n24778;
  assign n23678 = ~n23685;
  assign n23587 = ~n25532 | ~n23584;
  assign n23217 = n23223 ^ n23185;
  assign n25726 = ~n26914 & ~n41697;
  assign n25739 = ~n26916 & ~n25738;
  assign n25725 = ~n26916 & ~n25724;
  assign n24220 = ~n24241 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n25727 = ~n25758 | ~n34645;
  assign n25723 = ~n25717 | ~n25758;
  assign n25741 = ~n25758 | ~n35425;
  assign n23894 = ~n23945 | ~n23933;
  assign n23578 = ~n23577 | ~n23085;
  assign n23586 = ~n25094 | ~n23585;
  assign n25748 = ~n25747 | ~n25746;
  assign n25751 = ~n25745 | ~n25758;
  assign n25714 = ~n26914 & ~n28062;
  assign n25711 = ~n25758 | ~n43835;
  assign n25577 = ~n25758 | ~n25575;
  assign n26191 = ~n26505 & ~n26428;
  assign n27665 = ~n35446 | ~n35445;
  assign n41093 = ~n40738 | ~P3_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n25894 = ~n40708 | ~n43294;
  assign n23908 = ~n24130 & ~n22947;
  assign n24222 = ~n24134 & ~n24119;
  assign n25737 = ~n25731 | ~n25758;
  assign n24483 = ~n24482 & ~n24481;
  assign n27323 = ~n27322;
  assign n23938 = n23936 & n23945;
  assign n26193 = ~n26505 | ~n26157;
  assign n23905 = ~n23945;
  assign n24219 = ~n24655 | ~n34187;
  assign n25548 = ~n25547 | ~n39522;
  assign n25672 = ~n26916 & ~n25671;
  assign n25673 = ~n26914 & ~n28061;
  assign n25549 = ~n26914 & ~n33579;
  assign n25669 = ~n25758 | ~n26428;
  assign n23185 = ~n26505 | ~n23224;
  assign n24656 = ~n24655 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n24425 = ~n32232 | ~n39895;
  assign n27876 = ~n41873 | ~n42353;
  assign n40980 = ~n40202 & ~n35858;
  assign n26447 = ~n41873 & ~n26446;
  assign n27336 = ~n27334 | ~n27333;
  assign n23261 = ~n26505 | ~n23270;
  assign n23125 = ~n26505 | ~n26167;
  assign n25586 = ~n25758 | ~n25585;
  assign n26490 = ~n41873 & ~n33537;
  assign n25589 = ~n26916 & ~n25588;
  assign n25568 = ~n26916 & ~n25567;
  assign n25569 = ~n26914 & ~n34858;
  assign n27680 = n27683 ^ n32515;
  assign n28206 = ~n40120;
  assign n25734 = ~n25733 | ~n25732;
  assign n25590 = ~n26914 & ~n39656;
  assign n25754 = ~n25758 | ~n35963;
  assign n41932 = ~n41873 & ~n28208;
  assign n25627 = ~n26916 & ~n25626;
  assign n25628 = ~n26914 & ~n39651;
  assign n25624 = ~n25758 | ~n26384;
  assign n25493 = ~n32217 | ~n39522;
  assign n43727 = ~n43726 | ~n43725;
  assign n27601 = ~n27802 & ~n27600;
  assign n26450 = ~n41873 | ~n26449;
  assign n36973 = n27673 ^ P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n25762 = ~n25761 | ~n25760;
  assign n23223 = ~n26505 | ~n23267;
  assign n25765 = ~n25759 | ~n25758;
  assign n25086 = ~n40081 | ~P1_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n25083 = ~n40081 | ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n25842 = ~n40081 | ~P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n23504 = ~n23503 | ~n26184;
  assign n23126 = ~n23085 | ~n26282;
  assign n23918 = ~n24872 | ~n23916;
  assign n25077 = ~n40081 | ~P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n23904 = ~n24654 | ~n23906;
  assign n25080 = ~n40081 | ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n24194 = ~n40081 | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n24746 = ~n25895 & ~n24745;
  assign n27318 = ~n27316 | ~n35974;
  assign n24191 = ~n40081 | ~P1_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n24730 = ~n24872 & ~n24726;
  assign n26029 = ~n25995 | ~n25994;
  assign n32857 = ~n31825 | ~n31511;
  assign n24188 = ~n40081 | ~P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n35445 = ~n27661 | ~n27660;
  assign n23168 = ~n23085 | ~n34879;
  assign n24185 = ~n40081 | ~P1_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n25579 = ~n28191 | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n25580 = ~n41474 | ~P2_EAX_REG_3__SCAN_IN;
  assign n24130 = ~n24200;
  assign n27333 = ~n32501 | ~n27332;
  assign n28051 = ~n40081 | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n28048 = ~n40081 | ~P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n26909 = ~n41790 & ~n23127;
  assign n27035 = ~n40081 | ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n27032 = ~n40081 | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n26686 = ~n40081 | ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n31451 = ~n24208 & ~n24207;
  assign n25533 = ~n28191 | ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n25534 = ~n41474 | ~P2_EAX_REG_1__SCAN_IN;
  assign n27673 = ~n27672 ^ n32208;
  assign n26683 = ~n40081 | ~P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n25719 = ~n41474 | ~P2_EAX_REG_8__SCAN_IN;
  assign n25718 = ~n28191 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n27605 = ~n27603 | ~n33501;
  assign n27328 = ~n27327;
  assign n26143 = ~n40081 | ~P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n42745 = ~n23127 & ~n42753;
  assign n26034 = ~n40081 | ~P1_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n25940 = ~n40081 | ~P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n25937 = ~n40081 | ~P1_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n24199 = ~n31921 | ~n24406;
  assign n24329 = ~n24387 | ~n24749;
  assign n33357 = ~n23728 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n24179 = ~n40081 | ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n24176 = ~n40081 | ~P1_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n24411 = ~n24396 | ~n24395;
  assign n24182 = ~n40081 | ~P1_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n27795 = ~n27596 | ~n27599;
  assign n24170 = ~n28825 & ~P1_EBX_REG_0__SCAN_IN;
  assign n24732 = ~n24664 | ~n24663;
  assign n26505 = ~n23085;
  assign n25109 = ~n36688 & ~n25108;
  assign n31716 = ~n31715 | ~n44100;
  assign n25833 = ~n43721 | ~P1_EAX_REG_13__SCAN_IN;
  assign n24908 = ~n43721 | ~P1_EAX_REG_8__SCAN_IN;
  assign n25585 = ~n26341;
  assign n31056 = ~n37289 & ~n32149;
  assign n25059 = ~n43721 | ~P1_EAX_REG_12__SCAN_IN;
  assign n24983 = ~n43721 | ~P1_EAX_REG_10__SCAN_IN;
  assign n27249 = ~n27248 | ~n27656;
  assign n24946 = ~n43721 | ~P1_EAX_REG_9__SCAN_IN;
  assign n24729 = ~n25895 | ~n24728;
  assign n24118 = ~n24802 | ~n34097;
  assign n24405 = ~n34097 | ~n31382;
  assign n23851 = ~n31721 & ~n23916;
  assign n31921 = ~n32239 & ~n24149;
  assign n24607 = ~n24706 & ~n24658;
  assign n25093 = ~n36561;
  assign n24232 = ~n24394 & ~n31721;
  assign n23917 = ~n24706 | ~n24098;
  assign n23910 = ~n35466;
  assign n23085 = ~n43061 & ~n37289;
  assign n38909 = ~n37754 | ~P3_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n23909 = ~n34097 & ~n31721;
  assign n27747 = ~n27592 & ~n27591;
  assign n31448 = ~n24102 & ~n24101;
  assign n24745 = ~n39891 | ~n31721;
  assign n23896 = ~n24706 & ~n34187;
  assign n26223 = ~n34885 & ~n33579;
  assign n27792 = ~n29940 | ~n27610;
  assign n24856 = ~n43721 | ~P1_EAX_REG_6__SCAN_IN;
  assign n24846 = ~n43721 | ~P1_EAX_REG_5__SCAN_IN;
  assign n24836 = ~n24831 & ~n24830;
  assign n24834 = ~n43721 | ~P1_EAX_REG_4__SCAN_IN;
  assign n25995 = ~n43721 | ~P1_EAX_REG_16__SCAN_IN;
  assign n27614 = ~n27613 & ~n31801;
  assign n25494 = ~n43061 | ~n39522;
  assign n25575 = ~n26327;
  assign n26328 = ~n43061 | ~n26327;
  assign n23501 = ~n23321 | ~n23320;
  assign n26177 = ~n23512;
  assign n36561 = ~n23446 & ~n23445;
  assign n25062 = ~n38389 | ~n43294;
  assign n27613 = ~n32672 & ~n27803;
  assign n27611 = ~n27803;
  assign n35976 = ~n27282 ^ P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n27610 = ~n33501 | ~n33486;
  assign n35425 = ~n25236 | ~n25235;
  assign n26282 = ~n23121 & ~n23120;
  assign n27627 = ~n27796 & ~n29940;
  assign n24208 = ~n24406 | ~n31382;
  assign n24728 = ~n24727 | ~n24734;
  assign n24866 = ~n28810 & ~n24862;
  assign n27671 = ~n27657 | ~n32808;
  assign n24659 = ~n24569 | ~n24568;
  assign n24169 = ~n24235 & ~n31705;
  assign n26428 = ~n25668 | ~n25667;
  assign n24109 = ~n24802 | ~n39891;
  assign n27248 = ~n32808;
  assign n31803 = ~n31802 | ~n31801;
  assign n25710 = ~n25691 | ~n25690;
  assign n23052 = ~n23051 | ~n23050;
  assign n24099 = ~n24098 | ~n24097;
  assign n34645 = ~n25176 | ~n25175;
  assign n27320 = ~n27656 | ~P3_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n27660 = ~n32284 | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n26440 = ~n25528 | ~n25527;
  assign n25021 = ~n39592 & ~n43725;
  assign n28810 = ~n39892 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n33486 = ~n33487;
  assign n27788 = ~n27773 | ~n27772;
  assign n27805 = ~n27781 & ~n27780;
  assign n27595 = ~n30706 & ~n31801;
  assign n31805 = ~n32475 | ~n29940;
  assign n36546 = ~n25359 | ~n25358;
  assign n27591 = ~n29940 | ~n31801;
  assign n23083 = ~n23082 | ~n23081;
  assign n35963 = ~n25297 | ~n25296;
  assign n27656 = ~n27143 & ~n27142;
  assign n25837 = ~n25061 | ~P1_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n24985 = ~n38804 | ~n43294;
  assign n24733 = ~n24705 & ~n24704;
  assign n23486 = ~n23485 & ~n23484;
  assign n23414 = ~n23406 & ~n23405;
  assign n23446 = ~n23432 | ~n23431;
  assign n24391 = ~n22947 | ~n24488;
  assign n34164 = ~n23979 & ~n23978;
  assign n40038 = ~n34102 | ~n34101;
  assign n39981 = ~n34140 | ~n34139;
  assign n39989 = ~n34142 | ~n34141;
  assign n40011 = ~n34232 | ~n34231;
  assign n39967 = ~n34251 | ~n34250;
  assign n23277 = ~n23276 | ~n23275;
  assign n39939 = ~n34247 | ~n34246;
  assign n39970 = ~n34195 | ~n34194;
  assign n40000 = ~n34172 | ~n34171;
  assign n40014 = ~n34081 | ~n34080;
  assign n40022 = ~n34083 | ~n34082;
  assign n40025 = ~n34157 | ~n34156;
  assign n39992 = ~n34170 | ~n34169;
  assign n40033 = ~n34155 | ~n34154;
  assign n40003 = ~n34234 | ~n34233;
  assign n40049 = ~n34104 | ~n34103;
  assign n39978 = ~n34193 | ~n34192;
  assign n23485 = ~n23483 | ~n23482;
  assign n23442 = ~n23440 | ~n23439;
  assign n27380 = ~n27364 | ~n27363;
  assign n27379 = ~n27378 | ~n27377;
  assign n27440 = ~n27424 | ~n27423;
  assign n23370 = ~n23362 & ~n23361;
  assign n27079 = ~n27057 | ~n27056;
  assign n24948 = ~n37516 & ~n43725;
  assign n23080 = ~n23078 | ~n23077;
  assign n27559 = ~n27558 | ~n27557;
  assign n23402 = ~n23394 & ~n23393;
  assign n23049 = ~n23047 | ~n23046;
  assign n24489 = ~n24295 | ~n24294;
  assign n23338 = ~n23337 | ~n23336;
  assign n24488 = ~n24386 | ~n24385;
  assign n27410 = ~n27394 | ~n27393;
  assign n27314 = ~n27313 | ~n27312;
  assign n23936 = ~n23941 & ~n23942;
  assign n23944 = ~n23942 | ~n23941;
  assign n27529 = ~n27528 | ~n27527;
  assign n25061 = ~n25020 & ~n25019;
  assign n23406 = ~n23404 | ~n23403;
  assign n23027 = ~n23026 | ~n23025;
  assign n23336 = n23335 & n23334;
  assign n23351 = ~n23345 & ~n23344;
  assign n23078 = ~n26828 | ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n23361 = ~n23360 | ~n23359;
  assign n23238 = ~n26780 & ~n42787;
  assign n23061 = ~n23060 | ~n23059;
  assign n23301 = ~n23295 | ~n23294;
  assign n23310 = ~n23306 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23413 = ~n23412 & ~n23411;
  assign n23487 = ~n23480 & ~n23479;
  assign n31189 = ~U214;
  assign n27226 = ~n27225 & ~n27224;
  assign n27227 = ~n27219 & ~n27218;
  assign n24910 = ~n37243 | ~n43294;
  assign n25020 = ~n24981 | ~P1_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n25619 = ~n25615 | ~n25614;
  assign n25612 = ~n25611 | ~n25610;
  assign n27409 = ~n27408 | ~n27407;
  assign n23963 = ~n23955 & ~n23954;
  assign n23977 = ~n23969 & ~n23968;
  assign n24089 = ~n24081 & ~n24080;
  assign n27770 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n27760;
  assign n27446 = ~n27442 | ~n27441;
  assign n27452 = ~n27448 | ~n27447;
  assign n23768 = ~n23756 | ~n23755;
  assign n27244 = ~n27243 & ~n27242;
  assign n23655 = ~n37853 | ~n39508;
  assign n24602 = ~n24598 | ~n24597;
  assign n24687 = ~n24683 | ~n24682;
  assign n24686 = ~n24685 | ~n24684;
  assign n23962 = ~n23961 & ~n23960;
  assign n23376 = ~n23372 | ~n23371;
  assign n24058 = ~n24057 | ~n24056;
  assign n24037 = ~n24026 | ~n24025;
  assign n23438 = ~n23434 | ~n23433;
  assign n23059 = ~n22926 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n23369 = ~n23368 & ~n23367;
  assign n23025 = ~n22926 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n23359 = ~n22926 | ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n23028 = ~n23024 & ~n35715;
  assign n23832 = ~n23824 | ~n23823;
  assign n23968 = ~n23967 | ~n23966;
  assign n23401 = ~n23400 & ~n23399;
  assign n23391 = ~n22926 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n23480 = ~n23476 | ~n23475;
  assign n23976 = ~n23975 & ~n23974;
  assign n23873 = ~n23861 | ~n23860;
  assign n23872 = ~n23871 | ~n23870;
  assign n23076 = ~n23072 | ~n23071;
  assign n24067 = ~n24063 | ~n24062;
  assign n24080 = ~n24079 | ~n24078;
  assign n23345 = ~n23341 | ~n23340;
  assign n23043 = ~n23038 | ~n23037;
  assign n23316 = ~n23315 & ~n23314;
  assign n23062 = ~n23058 & ~n35715;
  assign n24383 = ~n24382 | ~n24381;
  assign n23334 = ~n22926 | ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n23459 = ~n22926 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n23421 = ~n22926 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n23955 = ~n23951 | ~n23950;
  assign n23954 = ~n23953 | ~n23952;
  assign n23317 = ~n23312 & ~n23311;
  assign n23412 = ~n23408 | ~n23407;
  assign n23823 = ~n23822 & ~n23821;
  assign n27185 = ~n22903 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n23831 = ~n23830 | ~n23829;
  assign n27538 = ~n22903 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n27166 = ~n22903 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n23969 = ~n23965 | ~n23964;
  assign n23884 = ~n23883 | ~n23882;
  assign n23951 = ~n43241 | ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n24063 = ~n43241 | ~P1_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n23033 = ~n23032 | ~n23031;
  assign n27368 = ~n22919 | ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n23885 = ~n23881 | ~n23880;
  assign n23411 = ~n23410 | ~n23409;
  assign n23344 = ~n23343 | ~n23342;
  assign n23042 = ~n23041 | ~n23040;
  assign n24059 = ~n24047 | ~n24046;
  assign n23974 = ~n23973 | ~n23972;
  assign n27104 = ~n22903 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n27546 = ~n22919 | ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n27051 = ~n22903 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n23767 = ~n23766 | ~n23765;
  assign n23870 = ~n23869 & ~n23868;
  assign n27269 = ~n22903 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n23975 = ~n23971 | ~n23970;
  assign n23861 = ~n23855 & ~n23854;
  assign n23824 = ~n23820 & ~n23819;
  assign n27115 = ~n22903 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n24036 = ~n24035 | ~n24034;
  assign n27221 = ~n22903 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n27492 = ~n22919 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n24596 = ~n24592 | ~n24591;
  assign n24595 = ~n24594 | ~n24593;
  assign n24601 = ~n24600 | ~n24599;
  assign n27478 = ~n22903 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n27465 = ~n27464 | ~n27463;
  assign n39896 = ~P1_ADDRESS_REG_29__SCAN_IN | ~n22981;
  assign n23375 = ~n23374 | ~n23373;
  assign n27387 = ~n22903 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n24587 = ~n24586 | ~n24585;
  assign n27420 = ~n22919 | ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n23067 = ~n23066 | ~n23065;
  assign n27418 = ~n22903 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n23075 = ~n23074 | ~n23073;
  assign n23068 = ~n23064 | ~n23063;
  assign n27760 = ~n27759 | ~n27758;
  assign n24361 = ~n24360 | ~n24359;
  assign n27451 = ~n27450 | ~n27449;
  assign n23312 = ~n26818 & ~n43085;
  assign n23437 = ~n23436 | ~n23435;
  assign n24440 = ~n24439 | ~n24438;
  assign n27508 = ~n22903 | ~P3_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n23837 = ~n23836 | ~n23835;
  assign n27518 = ~n22919 | ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n23210 = ~n25687 & ~n41805;
  assign n23838 = ~n23834 | ~n23833;
  assign n27358 = ~n22903 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n27562 = ~n22903 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n27572 = ~n27568 | ~n27567;
  assign n27564 = ~n22919 | ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n23435 = ~n26858 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n27434 = ~n35392 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n27477 = ~n36317 | ~P3_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n24251 = ~n24250 & ~n24249;
  assign n27433 = ~n22920 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n23366 = ~n23467 | ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n27073 = ~n22902 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n25687 = ~n23458;
  assign n27480 = ~n36310 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n27426 = ~n22917 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n23903 = ~n24100 & ~n33710;
  assign n23363 = ~n23464 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n27472 = ~n36294 | ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n27488 = ~n22917 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n27487 = ~n35392 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n23371 = ~n26832 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n27491 = ~n22923 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n26820 = ~n26832;
  assign n23298 = ~n26848 | ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n24229 = ~n24228 | ~n24227;
  assign n23117 = ~n25641 & ~n23114;
  assign n27251 = ~n36299 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n27258 = ~n36286 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n27260 = ~n35392 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n23477 = ~n26858 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n27137 = ~n35392 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n23184 = ~n23182 | ~n23181;
  assign n38059 = ~n38062 & ~n43722;
  assign n22925 = ~n26853;
  assign n27411 = ~n22923 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n23073 = ~n26858 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n23071 = ~n26832 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n24453 = ~n43260 | ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n27081 = ~n22902 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n31825 = ~n32867;
  assign n27273 = ~n22902 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n32880 = ~n36415 | ~n35842;
  assign n23340 = ~n26832 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n27523 = ~n35392 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n36363 = ~n28159 & ~n28158;
  assign n27353 = ~n35392 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n27359 = ~n22923 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n23860 = ~n23859 & ~n23858;
  assign n23871 = ~n23865 & ~n23864;
  assign n27548 = ~n22917 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n27547 = ~n35392 | ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n27552 = ~n36294 | ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n27553 = ~n22923 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n24084 = ~n43261 | ~P1_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n27503 = ~n22923 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n23970 = ~n43260 | ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n23971 = ~n43270 | ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n27583 = ~n22902 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n27561 = ~n36307 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n27584 = ~n36294 | ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n27582 = ~n36310 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n23409 = ~n26858 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n27577 = ~n22923 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n23964 = ~n43246 | ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n23957 = ~n43275 | ~P1_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n23037 = ~n26832 | ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n27389 = ~n35392 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n27145 = ~n22902 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n23040 = ~n26858 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n24083 = ~n43270 | ~P1_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n27570 = ~n22917 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n23972 = ~n43261 | ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n27569 = ~n35392 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n27397 = ~n22923 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n23830 = ~n23826 & ~n23825;
  assign n24082 = ~n43260 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n27510 = ~n22917 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n27199 = ~n22902 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n43729 = ~n29569 | ~n39315;
  assign n27232 = ~n34773 & ~n27228;
  assign n27231 = ~n27230 & ~n27229;
  assign n32867 = ~n27782 | ~n29436;
  assign n23296 = ~n26807 & ~n26768;
  assign n23374 = ~n26838 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n23365 = ~n23468 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n35804 = ~P2_STATE2_REG_1__SCAN_IN & ~n28155;
  assign n23041 = ~n26838 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n34515 = ~n24209 & ~P1_STATE_REG_0__SCAN_IN;
  assign n41310 = ~n39529 & ~n39114;
  assign n41560 = ~n40865 & ~n40723;
  assign n24838 = ~n35518 & ~n43725;
  assign n22905 = ~n26848;
  assign n23182 = ~n23123 | ~n23122;
  assign n23074 = ~n26838 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n27188 = ~n27288 & ~n27187;
  assign n27183 = ~n27230 & ~n27182;
  assign n27256 = ~n27288 & ~n27255;
  assign n23891 = ~n23900 | ~n23850;
  assign n27118 = ~n27288 & ~n27117;
  assign n23829 = ~n23828 & ~n23827;
  assign n22907 = ~n24517;
  assign n23877 = ~n43271 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n27101 = ~n27288 & ~n27100;
  assign n29305 = n29245 & n29244;
  assign n27096 = ~n27095 & ~n27094;
  assign n28494 = ~n41999;
  assign n27748 = ~n40127 | ~n36190;
  assign n31495 = n36357 & n35811;
  assign n22908 = ~n27009;
  assign n24506 = ~n24505;
  assign n43499 = ~n23019 & ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n23275 = ~n23270;
  assign n29439 = ~n29308;
  assign n22927 = ~n23720 | ~n35718;
  assign n23077 = ~n23481 | ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n24833 = ~n43294 & ~n24832;
  assign n22912 = ~n35408;
  assign n27061 = ~n27069;
  assign n27539 = ~n36311 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n36316 = ~n27068 | ~n36052;
  assign n24510 = ~n24509 | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n29553 = ~n29175;
  assign n24825 = ~n35889 & ~n43725;
  assign n24438 = ~n24509 | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n39310 = ~n24248 | ~n34476;
  assign n24228 = ~n26587 | ~n39937;
  assign n23631 = ~n31488 & ~n38277;
  assign n44099 = ~n32136 & ~n33710;
  assign n27431 = ~n36311 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n29721 = ~n29580;
  assign n27479 = ~n36311 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n23608 = ~n31488 & ~n39114;
  assign n26862 = n23105 & n23103;
  assign n23570 = ~n31488 & ~n37635;
  assign n23943 = ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n33734;
  assign n23942 = ~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN | ~n24830;
  assign n35630 = ~n43722 | ~n33714;
  assign n23932 = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n37475;
  assign n25114 = ~n37805 & ~n35254;
  assign n27757 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~n41341;
  assign n24864 = ~n43722 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n26877 = ~n23039 | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n43496 = ~n32506 & ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n23183 = ~n37634 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23720 = ~n23045;
  assign n27058 = ~n33933 | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n36311 = ~n36049 & ~n29442;
  assign n40127 = ~n40959 & ~n40981;
  assign n35811 = ~n31055 | ~n39511;
  assign n36366 = ~P2_STATE2_REG_2__SCAN_IN | ~n31055;
  assign n31488 = ~n36357 | ~n31055;
  assign n26174 = ~P2_FLUSH_REG_SCAN_IN & ~n31055;
  assign n24436 = ~n34476;
  assign n42011 = ~P3_STATE2_REG_3__SCAN_IN | ~n32362;
  assign n24504 = ~n37475 | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n24248 = ~n34677 | ~n39937;
  assign n35802 = ~n36364;
  assign n37023 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN | ~P3_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n27182 = ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n27181 = ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n36364 = ~READY21_REG_SCAN_IN | ~READY12_REG_SCAN_IN;
  assign n24842 = ~P1_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n23039 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n24829 = P1_PHYADDRPOINTER_REG_1__SCAN_IN & P1_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n34550 = ~P1_STATE2_REG_2__SCAN_IN | ~P1_STATE2_REG_1__SCAN_IN;
  assign n31507 = ~P3_STATE2_REG_2__SCAN_IN | ~P3_STATE2_REG_1__SCAN_IN;
  assign n41671 = ~P3_STATE2_REG_0__SCAN_IN;
  assign n33842 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN | ~P3_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n40196 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n31667 = ~READY22_REG_SCAN_IN | ~READY2;
  assign n40998 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n27117 = ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n26099 = ~P1_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n29726 = ~P3_STATE2_REG_2__SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN;
  assign n28755 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN | ~P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n34476 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n29997 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n41341 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n29171 = ~P2_ADDRESS_REG_29__SCAN_IN;
  assign n27153 = ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n31953 = ~P3_EBX_REG_5__SCAN_IN | ~P3_EBX_REG_6__SCAN_IN;
  assign n33734 = ~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n36307 = ~n27070 & ~n27061;
  assign n23665 = ~n23634 | ~n23633;
  assign n23634 = ~n23617 & ~n23616;
  assign n42746 = n42747 ^ n42748;
  assign n42747 = ~n41785 | ~n41784;
  assign n34726 = n24575 ^ n24610;
  assign n43864 = ~n43914 | ~n43876;
  assign n43905 = ~n43898 | ~n43913;
  assign n43898 = ~n43875 | ~n43874;
  assign n43795 = ~n43728 ^ n43727;
  assign n43728 = ~n43720 | ~n43719;
  assign n32238 = ~n24061 | ~n24060;
  assign n27070 = ~n35663 | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n36295 = ~n27071 & ~n33502;
  assign n23724 = ~n23490;
  assign n36306 = ~n27061 & ~n33502;
  assign n34576 = n24499 ^ n24497;
  assign n22920 = ~n35408;
  assign n22921 = ~n22912;
  assign n22922 = ~n22920;
  assign n40306 = ~n23668 ^ n23667;
  assign n36299 = ~n33502 & ~n29442;
  assign n26235 = n23613 ^ n23614;
  assign n22924 = ~n22927 & ~n35715;
  assign n23019 = ~n26153 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23571 = ~n26546 & ~n26505;
  assign n24743 = ~n24742;
  assign n24406 = ~n34164 & ~n31891;
  assign n24508 = ~n26587;
  assign n24115 = ~n31921 & ~n34164;
  assign n24426 = ~n24424;
  assign n23583 = ~n23569 | ~n35707;
  assign n23566 = ~n23731 & ~n23565;
  assign n23603 = ~n23552 | ~n23551;
  assign n42197 = ~n42305 | ~n42303;
  assign n27860 = ~n26391 | ~n26390;
  assign n23709 = ~n23708 | ~n23707;
  assign n23708 = ~n23705 | ~n36561;
  assign n27689 = n32515 | n27683;
  assign n42002 = ~n42501 | ~n41995;
  assign n25936 = ~n25841 | ~n25840;
  assign n42285 = n36385 ^ n36384;
  assign n42066 = ~n39481 ^ n39480;
  assign n40395 = ~n40394 | ~n40393;
  assign n27668 = ~n27667;
  assign n41332 = ~n41331 & ~n41330;
  assign n43379 = n43559 & n43378;
  assign n25076 = n24196 ^ n40073;
  assign n37000 = ~n25962 ^ n24755;
  assign n35821 = ~n35823 & ~n35822;
  assign n43016 = n39701 ^ n39700;
  assign n39671 = ~n38969 & ~n38968;
  assign n42872 = n36373 ^ n26913;
  assign n38016 = ~n25487;
  assign n37839 = ~n36577 & ~n37947;
  assign n34906 = ~n37363;
  assign n36625 = ~n36802 | ~BUF2_REG_25__SCAN_IN;
  assign n36579 = ~n36802 | ~BUF2_REG_26__SCAN_IN;
  assign n24631 = ~n28775 | ~P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n24630 = ~n43264 | ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n24633 = ~n43245 | ~P1_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n24624 = ~n43271 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n24625 = ~n22915 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n24626 = ~n43275 | ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n24640 = ~n22908 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n24641 = ~n43274 | ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n24639 = ~n22907 | ~P1_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n24679 = ~n28775 | ~P1_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n24678 = ~n22915 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n24677 = ~n43246 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n24599 = ~n43271 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n24600 = ~n43260 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n24598 = ~n43265 | ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n24591 = ~n22908 | ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n24592 = ~n43270 | ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n24594 = ~n43275 | ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n24585 = ~n43246 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n24586 = ~n43251 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n24583 = ~n43245 | ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n23172 = ~n24775 | ~n23171;
  assign n25615 = ~n26831 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n25614 = ~n26827 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n25616 = ~n26841 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n25611 = ~n26852 | ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n25595 = ~n26828 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n23191 = ~n26831 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n23190 = ~n26852 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n23204 = ~n26858 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n23092 = ~n26831 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n23091 = ~n26852 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n23096 = ~n26837 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n23097 = ~n26827 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n23108 = ~n26726 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n23110 = ~n26858 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n23897 = P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n27003 = ~P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n27010 = ~P1_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n24717 = ~n24851;
  assign n24576 = ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n23853 = ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n23857 = ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n25285 = ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n25635 = ~n23481 | ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n25636 = ~n26849 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n23245 = ~n22906 | ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n23232 = ~n26858 | ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n23235 = ~n26726 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n27228 = ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n27537 = ~n36317 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n27533 = ~n36320 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n27462 = ~n22917 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n27464 = ~n22914 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n27457 = ~n22923 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n27458 = ~n22913 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n27456 = ~n36294 | ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n27443 = ~n22920 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n24726 = ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n24027 = ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n24735 = ~n24734 ^ n24747;
  assign n35325 = ~n35324;
  assign n24133 = ~n24216;
  assign n24333 = ~n24298 & ~n24297;
  assign n24296 = ~n24489;
  assign n24485 = ~n24333 & ~n24334;
  assign n31891 = ~n24016 | ~n24015;
  assign n24015 = n24014 & n24013;
  assign n33720 = ~n33717 | ~n33721;
  assign n33719 = ~n33718 | ~n34495;
  assign n33717 = ~n34495;
  assign n23591 = ~n28346;
  assign n43099 = ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n25559 = ~n25557;
  assign n28284 = ~n39573 | ~P2_EBX_REG_19__SCAN_IN;
  assign n42204 = n40676 ^ n40675;
  assign n42094 = n40652 ^ n40651;
  assign n42084 = ~n42083 | ~n42082;
  assign n38945 = n27882 ^ n27881;
  assign n26499 = ~n26498 & ~n26497;
  assign n26496 = ~n39727;
  assign n23534 = ~n25099;
  assign n23321 = ~n23301 & ~n23300;
  assign n23490 = ~n23384 & ~n23383;
  assign n23383 = ~n23382 | ~n23381;
  assign n26167 = n23182 ^ n23124;
  assign n23124 = ~n23181;
  assign n35771 = ~n35768 | ~n35767;
  assign n35772 = ~n35717 | ~n35716;
  assign n27388 = ~n22902 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n27384 = ~n22919 | ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n27383 = ~n22917 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n27381 = ~n22920 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n27765 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n27521 = ~n36320 | ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n27516 = ~n36294 | ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n27501 = ~n36311 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n27502 = ~n22902 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n27413 = ~n36320 | ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n27414 = ~n36310 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n27594 = ~n27604;
  assign n27374 = ~n36320 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n27373 = ~n36311 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n40823 = ~n39774 | ~n39773;
  assign n39773 = ~n40471 | ~n40968;
  assign n41349 = ~n41348 | ~n41347;
  assign n41348 = ~n41343 | ~n41342;
  assign n24171 = n24168 ^ n28825;
  assign n26634 = ~n26600 | ~n26599;
  assign n26600 = ~n43721 | ~P1_EAX_REG_18__SCAN_IN;
  assign n24874 = ~n25928;
  assign n25023 = ~n28608 | ~P1_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n37500 = ~n36273 | ~n36272;
  assign n24848 = n36110 & n43294;
  assign n34344 = ~n33794 & ~n33793;
  assign n40079 = ~n42981;
  assign n42483 = ~n43462 | ~P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n41435 = ~n41437 | ~n41436;
  assign n26146 = n26145 ^ n28825;
  assign n26715 = ~n26147 & ~n26146;
  assign n26142 = ~n25944 & ~n25943;
  assign n25984 = ~n25936 & ~n25935;
  assign n25841 = ~n37532 & ~n37531;
  assign n37219 = n25082 ^ n40073;
  assign n36905 = ~n43462 ^ P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n23888 = ~n23873 & ~n23872;
  assign n24388 = n24734 ^ n24488;
  assign n24443 = ~n24441 & ~n24440;
  assign n24503 = ~n24435;
  assign n24117 = ~n24130 & ~n31382;
  assign n31903 = ~n31902 | ~n31901;
  assign n23979 = ~n23963 | ~n23962;
  assign n33716 = ~n34485 | ~n33714;
  assign n34505 = ~n34504 | ~n34503;
  assign n23510 = n23220 ^ P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n23220 = ~n23266;
  assign n26195 = ~n26194 | ~n26193;
  assign n28277 = ~n39573 | ~P2_EBX_REG_18__SCAN_IN;
  assign n42256 = n39211 ^ n39210;
  assign n40282 = n28199 ^ n28198;
  assign n39461 = ~n27889 ^ n27888;
  assign n37329 = n27879 ^ n27878;
  assign n28271 = ~n39573 | ~P2_EBX_REG_17__SCAN_IN;
  assign n25222 = ~n25214 | ~n25213;
  assign n25234 = ~n25230 | ~n25229;
  assign n25159 = ~n25158 | ~n25157;
  assign n25160 = ~n25156 | ~n25155;
  assign n25162 = ~n25154 & ~n25153;
  assign n25174 = ~n25170 | ~n25169;
  assign n25169 = ~n25168 & ~n25167;
  assign n42749 = ~n42748;
  assign n43829 = ~n43828;
  assign n43613 = ~n43163 | ~n43162;
  assign n28309 = ~n39702;
  assign n37466 = ~n37269;
  assign n28282 = ~n36395;
  assign n42202 = ~n42236;
  assign n23729 = ~n23500 & ~n23499;
  assign n23500 = ~n23547;
  assign n23714 = ~n23713 | ~n44000;
  assign n26209 = ~n26207 | ~n26506;
  assign n37796 = ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n42782 = ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n39525 = ~n39523 | ~n39522;
  assign n39528 = ~n39527;
  assign n27255 = ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n40861 = ~n41146;
  assign n27347 = ~n27344 ^ n27343;
  assign n27677 = n32501 ^ n27655;
  assign n27317 = ~n32284 | ~n36352;
  assign n39788 = ~n41542 | ~n39785;
  assign n40412 = ~n41542 | ~n40411;
  assign n40210 = ~n39448;
  assign n39401 = ~n39400 | ~n40226;
  assign n27685 = ~n27684;
  assign n40269 = ~n40174 | ~n40173;
  assign n38594 = ~n40422 | ~n40170;
  assign n43374 = ~n43797 | ~P1_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n28820 = ~n28774 | ~n28773;
  assign n28044 = ~n28512 | ~n28511;
  assign n28512 = ~n27029 & ~n27028;
  assign n26680 = ~n26712 | ~n26711;
  assign n28485 = ~n26680 & ~n26679;
  assign n26138 = ~n26092 | ~n26091;
  assign n25850 = ~n25065 | ~n25064;
  assign n36900 = n25079 ^ n28825;
  assign n37220 = ~n36901 & ~n36900;
  assign n34814 = ~n34344 | ~n34343;
  assign n41898 = ~n28485 ^ n28484;
  assign n25992 = n25934 & n25933;
  assign n37536 = ~n37214 | ~n37213;
  assign n31908 = ~n31907;
  assign n43571 = n43720 ^ n43718;
  assign n28854 = ~n28852;
  assign n28505 = ~n42500 & ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n26581 = ~n26580;
  assign n25975 = ~n38383;
  assign n38798 = ~n38799;
  assign n37551 = n37500 ^ n37499;
  assign n43359 = n42977 ^ P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n43135 = n43449 ^ n42975;
  assign n42551 = n42979 ^ n40072;
  assign n28723 = ~n42979;
  assign n42815 = n42548 ^ n42005;
  assign n42833 = n28523 ^ n28522;
  assign n42680 = n41435 ^ n28047;
  assign n41127 = n25984 ^ n25983;
  assign n37498 = ~n36905 ^ n36904;
  assign n35237 = ~n35169 | ~n35168;
  assign n38406 = ~n39818 | ~n38405;
  assign n28196 = ~n22900 & ~n37289;
  assign n40932 = ~n43192 | ~n41934;
  assign n37729 = ~n37728 | ~n37727;
  assign n37727 = ~n38898 | ~n41942;
  assign n37728 = ~n42872 | ~n40602;
  assign n23663 = ~n23662;
  assign n23605 = ~n23597 & ~n23596;
  assign n41657 = ~n43584;
  assign n41565 = ~n41564;
  assign n36377 = ~n36373;
  assign n42219 = n35376 ^ n35316;
  assign n35380 = ~n35376;
  assign n42564 = ~n42069 ^ n42068;
  assign n43667 = ~n43664 & ~n43663;
  assign n43224 = n39757 ^ n39756;
  assign n42857 = ~n37460 ^ n37459;
  assign n42516 = ~n37265 ^ n37264;
  assign n42515 = n42472 ^ P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n42437 = n42286 ^ n42346;
  assign n42288 = ~n42287 | ~n43583;
  assign n42526 = ~n42727 | ~n42292;
  assign n42612 = ~n37445 ^ n37444;
  assign n42611 = n42279 ^ n42259;
  assign n42259 = ~n42280 | ~n42278;
  assign n42632 = ~n42388 ^ n42387;
  assign n42111 = ~n43158 | ~n43150;
  assign n42139 = ~n42103 ^ n42102;
  assign n36613 = n36852 ^ n36851;
  assign n36846 = ~n26216 | ~n42110;
  assign n27100 = ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n39445 = ~n38147 ^ n37022;
  assign n28091 = ~n41113 | ~n41546;
  assign n40241 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~n40240;
  assign n40239 = ~n37766 ^ n37765;
  assign n40253 = ~n41006 | ~n40252;
  assign n40331 = ~n40226 | ~n40225;
  assign n40229 = n36211 ^ P3_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n40963 = ~n40982 | ~n40961;
  assign n40972 = ~n40971 | ~n40970;
  assign n41537 = ~n27620 & ~n27619;
  assign n40374 = ~n40372 | ~n41546;
  assign n39631 = ~n39630 | ~n39629;
  assign n43575 = ~n43791 | ~P1_REIP_REG_30__SCAN_IN;
  assign n28879 = ~n43371 | ~P1_REIP_REG_28__SCAN_IN;
  assign n28533 = ~n28532 | ~n28531;
  assign n42180 = ~n42179 | ~n42178;
  assign n37520 = ~n37515 | ~n43033;
  assign n36115 = ~n36114 | ~n36113;
  assign n35887 = ~n35886 | ~n35885;
  assign n36149 = ~n36148 | ~n36147;
  assign n35512 = ~n43566;
  assign n42941 = ~n28774 ^ n28773;
  assign n28660 = ~n28774;
  assign n28465 = ~n28835;
  assign n26693 = ~n41969 | ~n44021;
  assign n26713 = ~n41454;
  assign n26717 = ~n41743 | ~n44021;
  assign n26150 = ~n41276 | ~n44021;
  assign n26033 = ~n41024;
  assign n26038 = ~n41022 | ~n44021;
  assign n41454 = n26712 ^ n26711;
  assign n41024 = n26092 ^ n26091;
  assign n40707 = ~n25993 ^ n25992;
  assign n39593 = n37536 ^ n37535;
  assign n43029 = ~n43462 ^ n43351;
  assign n42679 = n42504 ^ P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n41968 = n41952 ^ P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n40784 = n26565 ^ n25982;
  assign n26585 = ~n31361;
  assign n38659 = n38387 ^ n38386;
  assign n40795 = ~n40797 | ~n26562;
  assign n40793 = ~n40092 | ~n26563;
  assign n26572 = ~n26571 | ~n26570;
  assign n40099 = ~n43344 | ~n40098;
  assign n24757 = ~n24756 | ~n37006;
  assign n24756 = ~n36906 | ~n37000;
  assign n35836 = ~n35835 | ~n35834;
  assign n39765 = ~n43175 | ~n41934;
  assign n39754 = ~n39753 | ~n39752;
  assign n39704 = ~n43015;
  assign n42439 = n36396 ^ n36395;
  assign n36393 = ~n36392 | ~n36391;
  assign n38956 = ~n38955 | ~n38954;
  assign n39715 = ~n42857 | ~n43525;
  assign n39295 = ~n42516 | ~n43525;
  assign n42637 = ~n37356 ^ n37355;
  assign n42424 = n36553 ^ n36552;
  assign n38980 = n42517 & n41756;
  assign n38970 = n38969 & n38968;
  assign n25796 = ~n42872 | ~n41756;
  assign n38015 = ~n38014 | ~n38013;
  assign n40152 = n27852 ^ n28061;
  assign n42514 = ~n42708 ^ P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n42138 = n42656 ^ n42100;
  assign n39667 = n38376 ^ P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n37626 = ~n37625 | ~n37834;
  assign n37602 = ~n37601 | ~n37600;
  assign n37527 = ~n37526 | ~n37525;
  assign n37914 = ~n37913 | ~n37912;
  assign n37906 = ~n37905 | ~n37904;
  assign n37545 = ~n37544 | ~n37543;
  assign n37430 = ~n37429 | ~n37428;
  assign n37412 = ~n37411 | ~n37410;
  assign n37421 = ~n37420 | ~n37419;
  assign n37404 = ~n37403 | ~n37402;
  assign n38936 = ~n38935 | ~n38934;
  assign n38623 = ~n38622 | ~n38621;
  assign n40914 = ~n40913 | ~n40912;
  assign n40902 = ~n40901 | ~n40900;
  assign n40889 = ~n40888 | ~n40887;
  assign n41299 = ~n41298 | ~n41297;
  assign n41298 = ~P2_INSTQUEUE_REG_15__6__SCAN_IN | ~n41309;
  assign n41319 = ~n39548;
  assign n41287 = ~n41286 | ~n41285;
  assign n41286 = ~P2_INSTQUEUE_REG_15__7__SCAN_IN | ~n41309;
  assign n35941 = ~n41519 ^ n36162;
  assign n40810 = ~n41058;
  assign n36401 = ~n36403;
  assign n41398 = P3_INSTADDRPOINTER_REG_31__SCAN_IN ^ n27350;
  assign n41414 = ~n41401 | ~n41400;
  assign n37776 = ~n37772 | ~n37771;
  assign n38167 = ~n40744 | ~n39790;
  assign n38168 = ~n40743 | ~n39785;
  assign n38029 = ~n38142 | ~n40431;
  assign n37593 = ~n40743 | ~n40411;
  assign n40958 = ~n37109 | ~n37108;
  assign n40983 = ~n40982 | ~n40981;
  assign n40994 = ~n40993 | ~n42338;
  assign n40993 = ~n40992 | ~P3_STATE2_REG_2__SCAN_IN;
  assign n40992 = ~n40991 | ~n40990;
  assign n38589 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n38609 = ~n38608 | ~n38607;
  assign n41372 = ~n41371 | ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n26398 = ~n37039;
  assign n26393 = ~n38628;
  assign n26397 = ~n37654;
  assign n26392 = ~n36569;
  assign n25605 = ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n26346 = ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n28586 = ~P1_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n26100 = ~P1_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n24646 = ~n43242 | ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n24647 = ~n43246 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n24644 = ~n43260 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n24645 = ~n43251 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n24632 = ~n43261 | ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n24627 = ~n43270 | ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n24638 = ~n43265 | ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n24685 = ~n43245 | ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n24684 = ~n43270 | ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n24682 = ~n43251 | ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n24683 = ~n22907 | ~P1_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n24701 = ~n24697 | ~n24696;
  assign n24700 = ~n24699 | ~n24698;
  assign n24694 = ~n24693 | ~n24692;
  assign n24695 = ~n24691 | ~n24690;
  assign n24676 = ~n43242 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n24355 = ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n24364 = ~P1_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n24368 = ~P1_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n24378 = ~P1_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n24367 = ~P1_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n24356 = ~P1_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n26094 = ~P1_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n24267 = ~P1_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n24255 = ~P1_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n23131 = ~n23278 | ~n26167;
  assign n23174 = ~n33357 | ~n24775;
  assign n43085 = ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n26260 = ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n26405 = ~n38237;
  assign n26345 = ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n23289 = ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n23313 = ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n23355 = ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n23890 = n32083 ^ P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n23933 = ~n23929 ^ n23930;
  assign n23930 = P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ n37475;
  assign n26096 = ~P1_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n28616 = ~n28601 | ~n28600;
  assign n23761 = ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n23757 = ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n23762 = ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n43251 = ~n24526;
  assign n43245 = ~n27004;
  assign n43265 = ~n27011;
  assign n24578 = ~n43241 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n24577 = ~n22907 | ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n24580 = ~n43264 | ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n24579 = ~n43242 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n24597 = ~n43261 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n24593 = ~n22915 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n24584 = ~n43274 | ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n24613 = ~n24612 & ~n24611;
  assign n24345 = ~P1_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n24363 = ~P1_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n23862 = ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n23867 = ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n23866 = ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n23863 = ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n28592 = ~P1_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n24210 = ~n24209;
  assign n24373 = ~P1_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n24341 = ~P1_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n24377 = ~P1_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n24352 = ~P1_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n24342 = ~P1_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n24346 = ~P1_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n24374 = ~P1_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n24264 = ~P1_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n24275 = ~P1_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n43260 = ~n27006;
  assign n43261 = ~n24539;
  assign n43274 = ~n28585;
  assign n43264 = ~n26659;
  assign n43241 = ~n24515;
  assign n43242 = ~n24527;
  assign n40587 = ~n40676 | ~n40675;
  assign n28202 = ~P2_EBX_REG_15__SCAN_IN;
  assign n26301 = ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n25676 = ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n43086 = ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n41805 = ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n26790 = ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n26768 = ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n41588 = ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n26396 = ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n25657 = ~n26862 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n25658 = ~n26859 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n25660 = ~n25656 & ~n43407;
  assign n25617 = ~n22906 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n25613 = ~n25609 | ~n25608;
  assign n25599 = ~n25598 | ~n25597;
  assign n42787 = ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n26232 = ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n25517 = ~n23481 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n25518 = ~n26849 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n25506 = ~n26862 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n25507 = ~n26859 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n25508 = ~n25645 & ~n26260;
  assign n43172 = ~n43536;
  assign n28201 = ~P2_EBX_REG_13__SCAN_IN;
  assign n25697 = ~n22926 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n23198 = ~n23197 | ~n23196;
  assign n23199 = ~n23195 | ~n23194;
  assign n23193 = ~n23189 | ~n23188;
  assign n23208 = ~n23207 | ~n23206;
  assign n23089 = ~n26848 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n23098 = ~n22906 | ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n23112 = ~n23111 | ~n23110;
  assign n41631 = ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n26298 = ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n23128 = n37635 ^ P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n23181 = n37634 ^ P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n27761 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n29449;
  assign n27600 = ~n27599;
  assign n27603 = ~n27616 | ~n27611;
  assign n27339 = ~n32515 ^ n27333;
  assign n27551 = ~n36310 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n27554 = ~n36298 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n27563 = ~n36298 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n27568 = ~n36317 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n27473 = ~n22920 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n27493 = ~n36320 | ~P3_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n27494 = ~n22902 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n23898 = ~n39937 | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n24098 = n23891 ^ n23890;
  assign n43239 = ~n28807 | ~n28806;
  assign n24053 = ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n24049 = ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n24048 = ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n24052 = ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n24043 = ~P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n24038 = ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n24042 = ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n24021 = ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n24022 = ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n24017 = ~P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n27971 = ~n27937 | ~n27936;
  assign n26978 = ~n26944 | ~n26943;
  assign n26944 = ~n43721 | ~P1_EAX_REG_20__SCAN_IN;
  assign n23752 = ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n23749 = ~P1_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n25926 = ~n25925 | ~n25924;
  assign n25927 = ~n25911 | ~n25910;
  assign n25896 = ~n25895;
  assign n24978 = ~n24977 | ~n24976;
  assign n24982 = ~n28608 | ~P1_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n24941 = ~n24940 | ~n24939;
  assign n24945 = ~n28608 | ~P1_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n24903 = ~n24902 | ~n24901;
  assign n24904 = ~n24888 | ~n24887;
  assign n24907 = ~n28608 | ~P1_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n24859 = ~n25897 ^ n24731;
  assign n24845 = ~n28608 | ~P1_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n24823 = ~n24817 | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n43456 = ~n43462 ^ P1_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n24718 = n24732 ^ n24733;
  assign n24418 = ~n24416;
  assign n24137 = ~n24406;
  assign n23852 = ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n23856 = ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n24387 = ~n24477;
  assign n24734 = ~n24749;
  assign n24238 = ~n24234;
  assign n24242 = ~n24241;
  assign n24233 = ~n24231;
  assign n24480 = ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n34682 = ~n34717;
  assign n33709 = ~n35630 | ~n34550;
  assign n23266 = n23267 ^ P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23493 = ~n23724 | ~n23501;
  assign n23224 = n35715 ^ P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n28203 = ~P2_EBX_REG_17__SCAN_IN;
  assign n42209 = n40587 ^ n40586;
  assign n28200 = ~P2_EBX_REG_11__SCAN_IN;
  assign n26444 = ~n26459;
  assign n23136 = ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n26460 = n26459 ^ n26462;
  assign n28211 = ~n41879;
  assign n43426 = ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n25241 = ~n25240 | ~n25239;
  assign n25257 = ~n25256 | ~n25255;
  assign n25258 = ~n25254 | ~n25253;
  assign n26257 = ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n25167 = ~n25166 | ~n25165;
  assign n41602 = ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n41598 = ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n43092 = ~n43499;
  assign n41592 = ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n26819 = ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n25768 = ~n25758 | ~n36546;
  assign n25761 = ~n41474 | ~P2_EAX_REG_14__SCAN_IN;
  assign n25202 = ~n25198 | ~n25197;
  assign n25181 = ~n25180 | ~n25179;
  assign n25182 = ~n25178 | ~n25177;
  assign n25187 = ~n25186 | ~n25185;
  assign n25188 = ~n25184 | ~n25183;
  assign n25196 = ~n25194 | ~n25193;
  assign n25120 = ~n25119 | ~n25118;
  assign n25121 = ~n25117 | ~n25116;
  assign n25140 = ~n25136 | ~n25135;
  assign n25139 = ~n25138 | ~n25137;
  assign n25664 = ~n26831 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n25663 = ~n26827 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n25632 = ~n26780 & ~n25631;
  assign n23247 = ~n26832 | ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n23234 = ~n26838 | ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n25492 = ~n37635 | ~P2_STATE2_REG_3__SCAN_IN;
  assign n25524 = ~n22926 | ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n25523 = ~n26848 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n26271 = ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n23155 = ~n26849 | ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n43659 = ~n43606;
  assign n28291 = ~n23598 | ~P2_EBX_REG_20__SCAN_IN;
  assign n42099 = n40607 ^ n40606;
  assign n27885 = ~n27884 | ~n40762;
  assign n23723 = ~n23587 & ~n23586;
  assign n25685 = ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n25686 = ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n25703 = ~n26848 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n25681 = ~n26838 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n26391 = ~n26342 & ~n26341;
  assign n26390 = ~n26386 & ~n26385;
  assign n26476 = ~n36490 | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n23547 = ~n26200 & ~n25093;
  assign n26286 = ~n26285;
  assign n23169 = ~n26505 | ~n26154;
  assign n23458 = ~n22927 & ~n35715;
  assign n25692 = ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n23468 = ~n43100 & ~n35715;
  assign n26157 = n23130 ^ n23129;
  assign n23130 = ~n23128;
  assign n26159 = ~n23510;
  assign n27768 = ~n27767;
  assign n27417 = ~n36317 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n27049 = ~n36041;
  assign n34767 = ~P3_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n33298 = ~n22913;
  assign n27158 = ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n27151 = ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n27154 = ~n22919;
  assign n27157 = ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n27146 = ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n34766 = ~n36307;
  assign n27710 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN | ~P3_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n27345 = ~n39615 ^ n27342;
  assign n27366 = ~n36294 | ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n27365 = ~n36298 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n27367 = ~n22920 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n27357 = ~n36317 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n27360 = ~n22917 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n28747 = ~n28755 | ~n40968;
  assign n42323 = ~n40422 | ~n27642;
  assign n27229 = ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n27684 = ~n27689 ^ n35858;
  assign n27327 = ~n27250 ^ n32208;
  assign n27667 = n27666 ^ n32808;
  assign n27672 = ~n27671;
  assign n27798 = ~n27794 | ~n27793;
  assign n32198 = ~n33487 ^ n29940;
  assign n27545 = ~n22920 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n27540 = ~n22902 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n27531 = ~n36307 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n27447 = ~n36317 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n27449 = ~n36307 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n27466 = ~n27462 | ~n27461;
  assign n27463 = ~n35392 | ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n27459 = ~n27458 | ~n27457;
  assign n27444 = ~n36298 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n27578 = ~n36320 | ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n27485 = ~n36307 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n27486 = ~n36298 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n41330 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n26676 = ~n26671 | ~n28604;
  assign n26134 = ~n26129 | ~n28604;
  assign n25943 = n25942 ^ n28825;
  assign n24853 = ~n28608 | ~P1_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n24854 = ~n35681 | ~n43294;
  assign n24791 = ~n24790 | ~n24789;
  assign n24031 = ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n24028 = ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n26977 = ~n26976 | ~n43725;
  assign n28478 = ~n41949;
  assign n25836 = ~P1_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n25019 = ~P1_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n24798 = ~n24797 | ~n24796;
  assign n24797 = ~n43721 | ~P1_EAX_REG_1__SCAN_IN;
  assign n40072 = n42978 ^ n28825;
  assign n28720 = n28719 ^ n40073;
  assign n28719 = ~n28718 | ~n28717;
  assign n28669 = n28668 ^ n28825;
  assign n28668 = ~n28667 | ~n28666;
  assign n28832 = n28665 ^ n40073;
  assign n28663 = ~n40081 | ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n28522 = n28468 ^ n40073;
  assign n28466 = ~n40081 | ~P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n28054 = n28053 ^ n28825;
  assign n28052 = ~n40080 | ~P1_EBX_REG_23__SCAN_IN;
  assign n28523 = ~n28055 & ~n28054;
  assign n28550 = n28050 ^ n40073;
  assign n28049 = ~n40080 | ~P1_EBX_REG_22__SCAN_IN;
  assign n28047 = n27037 ^ n28825;
  assign n27036 = ~n40080 | ~P1_EBX_REG_21__SCAN_IN;
  assign n41436 = n27034 ^ n40073;
  assign n27033 = ~n40080 | ~P1_EBX_REG_20__SCAN_IN;
  assign n26689 = n26688 ^ n28825;
  assign n26687 = ~n40080 | ~P1_EBX_REG_19__SCAN_IN;
  assign n41437 = ~n26690 & ~n26689;
  assign n26714 = n26685 ^ n40073;
  assign n26141 = n26036 ^ n40073;
  assign n25983 = n25939 ^ n40073;
  assign n25935 = n25844 ^ n28825;
  assign n25840 = n25088 ^ n40073;
  assign n37532 = ~n37220 | ~n37219;
  assign n37531 = n25085 ^ n28825;
  assign n24753 = ~n24754;
  assign n24725 = ~n24724;
  assign n24740 = ~n24739;
  assign n34817 = n24190 ^ n40073;
  assign n24173 = ~n24171;
  assign n32549 = n24178 ^ n40073;
  assign n34058 = ~n34056 | ~n34055;
  assign n24494 = ~n34576 | ~n26568;
  assign n24157 = ~n42924 | ~n32552;
  assign n26568 = ~n24745;
  assign n31916 = ~n24162;
  assign n24103 = ~n31910;
  assign n24108 = ~n31921 | ~n31721;
  assign n32131 = ~n32080;
  assign n32116 = ~n31920 | ~n31919;
  assign n24125 = ~n26044 | ~n24121;
  assign n24121 = ~n24120 | ~n24222;
  assign n34691 = ~n39315 | ~n34685;
  assign n34685 = ~n34684 | ~n22916;
  assign n38403 = ~n38410;
  assign n38492 = n38484 & n38483;
  assign n38484 = ~n38482 | ~n39301;
  assign n38490 = ~n38557;
  assign n39316 = ~n39302;
  assign n38063 = ~n39316 | ~n39301;
  assign n34684 = n34679 & n34575;
  assign n34508 = ~n34494 | ~n34493;
  assign n23507 = ~n26157;
  assign n43668 = n41727 ^ n41726;
  assign n43607 = n41874 ^ n41212;
  assign n39764 = ~n40121 & ~n28206;
  assign n37274 = ~n37736 & ~n37735;
  assign n36385 = ~n39211 & ~n39210;
  assign n25746 = ~n28191 | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n25747 = ~n41474 | ~P2_EAX_REG_12__SCAN_IN;
  assign n40355 = n26488 ^ n26487;
  assign n26446 = ~P2_EBX_REG_4__SCAN_IN;
  assign n38821 = n26457 ^ n26456;
  assign n39569 = ~n28367 | ~n28366;
  assign n43512 = ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n43503 = ~n43100;
  assign n28264 = ~n39573 | ~P2_EBX_REG_16__SCAN_IN;
  assign n28257 = ~n39573 | ~P2_EBX_REG_15__SCAN_IN;
  assign n25327 = ~n25326 | ~n25325;
  assign n25328 = ~n25311 | ~n25310;
  assign n25281 = ~n25280 | ~n25279;
  assign n25295 = ~n25291 | ~n25290;
  assign n23592 = ~P2_REIP_REG_0__SCAN_IN;
  assign n23630 = ~n23603 & ~n23561;
  assign n28186 = ~n41724;
  assign n40921 = ~n28176 | ~n28175;
  assign n41564 = n41789 ^ n41569;
  assign n26923 = ~n26922 | ~n26921;
  assign n25788 = ~n25787 | ~n25786;
  assign n25784 = ~n41473 | ~P2_REIP_REG_18__SCAN_IN;
  assign n25487 = ~n38014 & ~n38013;
  assign n25732 = ~n28191 | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n25733 = ~n41474 | ~P2_EAX_REG_10__SCAN_IN;
  assign n26384 = ~n26449;
  assign n25558 = ~P2_STATE2_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n25491 = ~n25544;
  assign n28139 = ~P2_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n28136 = ~P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n28134 = ~P2_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n35971 = ~n35602 & ~n35601;
  assign n28127 = ~P2_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n28124 = ~P2_PHYADDRPOINTER_REG_4__SCAN_IN | ~n28118;
  assign n28125 = ~P2_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n23163 = ~n26848 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n23149 = ~n23148 | ~n23147;
  assign n23150 = ~n23146 | ~n23145;
  assign n23144 = ~n23140 | ~n23139;
  assign n23143 = ~n23142 | ~n23141;
  assign n43753 = n41933 ^ n41932;
  assign n28353 = ~n41732;
  assign n41940 = ~n28360 | ~n28359;
  assign n28336 = ~n39578 | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n28329 = ~n39578 | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n28330 = ~n28328 & ~n28327;
  assign n43584 = n39910 ^ n39909;
  assign n28321 = ~n39578 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n28314 = ~n39578 | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n28307 = ~n39578 | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n28305 = ~n28304 | ~n28303;
  assign n28300 = ~n39578 | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n28298 = ~n28297 | ~n28296;
  assign n28292 = ~n28291 | ~n28290;
  assign n26919 = ~n41473 | ~P2_REIP_REG_20__SCAN_IN;
  assign n42713 = ~n42717;
  assign n28285 = ~n28284 | ~n28283;
  assign n42716 = ~n42349 | ~n42348;
  assign n42347 = ~n42284 | ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n42348 = ~n42283 | ~n42282;
  assign n42283 = ~n42284;
  assign n25779 = ~n25778 | ~n25777;
  assign n42279 = ~n42255 | ~n42254;
  assign n42253 = ~n42252;
  assign n42257 = ~n42258;
  assign n25775 = ~n41473 | ~P2_REIP_REG_16__SCAN_IN;
  assign n42387 = n42252 ^ P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n42245 = ~n42662 | ~n42658;
  assign n26503 = ~n38374 | ~n26486;
  assign n26500 = ~n26499;
  assign n42382 = ~n42242;
  assign n36840 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n25544 = ~n23490 | ~n23501;
  assign n36489 = ~n36488 | ~n36840;
  assign n36486 = n26330 ^ P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n23645 = ~n26513 | ~n23644;
  assign n32944 = P2_INSTADDRPOINTER_REG_2__SCAN_IN ^ n26226;
  assign n32945 = n26285 ^ n26282;
  assign n25547 = ~n22904 | ~P2_EAX_REG_0__SCAN_IN;
  assign n41474 = ~n23415 & ~P2_STATE2_REG_3__SCAN_IN;
  assign n34879 = ~n34885;
  assign n23537 = ~n28150 | ~n23536;
  assign n23538 = n23534 & n23533;
  assign n43091 = ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n37620 = ~n38323 | ~n37951;
  assign n38237 = ~n26248 & ~n37302;
  assign n38329 = ~n26365;
  assign n37139 = ~n26371;
  assign n36746 = ~n26375;
  assign n37870 = ~n26354;
  assign n24777 = ~n24775;
  assign n38626 = ~n38278 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n37951 = P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ n23669;
  assign n36635 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n37362 = ~n36635;
  assign n26172 = ~n26171 | ~n26170;
  assign n26171 = ~n26169 | ~n31055;
  assign n23568 = ~n31493;
  assign n35777 = ~n35773 | ~n35772;
  assign n27396 = ~n36294 | ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n27398 = ~n36298 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n27390 = ~n36307 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n27382 = ~n36317 | ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n27402 = ~n36310 | ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n27790 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n27804 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ^ n29997;
  assign n27774 = ~n27766 ^ n27765;
  assign n31665 = ~n31670;
  assign n35641 = ~n35527 | ~n41682;
  assign n33741 = ~n33738 | ~n33739;
  assign n36164 = ~n41401 | ~n35930;
  assign n35408 = n27070 | n29442;
  assign n35420 = ~P3_EBX_REG_16__SCAN_IN;
  assign n33620 = ~P3_EBX_REG_8__SCAN_IN;
  assign n27507 = ~n36317 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n27509 = ~n22920 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n27524 = ~n36307 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n27515 = ~n36298 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n27504 = ~n36310 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n27428 = ~n22902 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n27425 = ~n36307 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n27412 = ~n36298 | ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n36310 = ~n27230;
  assign n36298 = ~n34042;
  assign n27187 = ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n27797 = ~n27795;
  assign n38905 = ~n38903;
  assign n32883 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN | ~P3_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n39450 = ~n37023;
  assign n40726 = ~n41403;
  assign n27321 = ~n27320;
  assign n27663 = ~n27662;
  assign n36664 = ~n27667 ^ P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n27319 = ~n32826 | ~n36526;
  assign n35446 = ~n27662 ^ P3_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n27352 = ~n22902 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n27351 = ~n36307 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n27372 = ~n36310 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n41407 = P3_INSTADDRPOINTER_REG_31__SCAN_IN ^ n27750;
  assign n28745 = ~n42337 | ~n40508;
  assign n40997 = ~n40826 | ~n40825;
  assign n37765 = ~n41149 ^ P3_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n39449 = ~n40221 | ~n39450;
  assign n39774 = ~n40422 | ~n39451;
  assign n40215 = ~n39388;
  assign n40213 = ~n39387;
  assign n40211 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN | ~n40210;
  assign n35861 = ~n27692 & ~n27691;
  assign n27690 = ~n36429;
  assign n36075 = n41149 ^ P3_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n35988 = ~n27686 ^ n27684;
  assign n36020 = n27680 ^ P3_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n40194 = ~n40178 | ~n40177;
  assign n27809 = ~n27808 | ~n33486;
  assign n27784 = ~n29940;
  assign n29841 = ~n42011 | ~n29447;
  assign n33502 = ~n35663 | ~n35608;
  assign n36294 = ~n27288;
  assign n41337 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n41351 = ~n41350 | ~n41349;
  assign n42160 = ~P1_REIP_REG_25__SCAN_IN | ~n42161;
  assign n28661 = n28471 ^ n28825;
  assign n28469 = ~n40081 | ~P1_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n42412 = ~n43559 | ~n42411;
  assign n42404 = ~P1_REIP_REG_23__SCAN_IN | ~n42403;
  assign n42184 = ~P1_REIP_REG_21__SCAN_IN | ~n28526;
  assign n41848 = ~P1_REIP_REG_19__SCAN_IN | ~n27840;
  assign n27843 = ~n41955 | ~n43559;
  assign n27841 = ~n27840 | ~n41894;
  assign n26702 = ~n41196 | ~n43559;
  assign n27836 = ~P1_REIP_REG_16__SCAN_IN | ~n41020;
  assign n40703 = ~P1_REIP_REG_14__SCAN_IN | ~n41125;
  assign n37241 = ~P1_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n34823 = ~P1_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n36990 = ~n35512 | ~n36982;
  assign n26065 = ~n31895 | ~n39944;
  assign n39942 = ~n35165 ^ n31936;
  assign n28656 = ~n28653 | ~n28652;
  assign n28461 = ~n28458 | ~n28457;
  assign n27026 = ~n27025 | ~n27024;
  assign n25849 = ~n25839 & ~n25838;
  assign n33791 = n24184 ^ n40073;
  assign n31794 = n24171 ^ n24172;
  assign n31697 = ~n24172;
  assign n25071 = ~n25070 | ~n25069;
  assign n28858 = ~n28835 ^ n28834;
  assign n28735 = ~n28525 ^ n28524;
  assign n42173 = ~n28512 ^ n28511;
  assign n26633 = ~n26632 | ~n43725;
  assign n26028 = ~n26027 | ~n43725;
  assign n37242 = ~n37001;
  assign n31360 = ~n31359 | ~n34515;
  assign n31359 = ~n32080 | ~n34517;
  assign n43712 = P1_PHYADDRPOINTER_REG_31__SCAN_IN ^ n26061;
  assign n43558 = P1_PHYADDRPOINTER_REG_30__SCAN_IN ^ n43293;
  assign n43138 = ~P1_PHYADDRPOINTER_REG_29__SCAN_IN ^ n28816;
  assign n43046 = ~P1_PHYADDRPOINTER_REG_28__SCAN_IN ^ n28714;
  assign n43378 = P1_PHYADDRPOINTER_REG_27__SCAN_IN ^ n28654;
  assign n28860 = ~P1_PHYADDRPOINTER_REG_26__SCAN_IN ^ n28612;
  assign n43035 = P1_PHYADDRPOINTER_REG_25__SCAN_IN ^ n28459;
  assign n28737 = ~P1_PHYADDRPOINTER_REG_24__SCAN_IN ^ n28413;
  assign n28731 = ~n22933 | ~P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n42410 = ~P1_PHYADDRPOINTER_REG_23__SCAN_IN ^ n28036;
  assign n42174 = ~P1_PHYADDRPOINTER_REG_22__SCAN_IN ^ n27972;
  assign n42507 = P1_PHYADDRPOINTER_REG_21__SCAN_IN ^ n26982;
  assign n42498 = ~n43462 | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n41899 = P1_PHYADDRPOINTER_REG_20__SCAN_IN ^ n26979;
  assign n41955 = P1_PHYADDRPOINTER_REG_19__SCAN_IN ^ n26637;
  assign n41444 = ~P1_PHYADDRPOINTER_REG_18__SCAN_IN ^ n26598;
  assign n41196 = P1_PHYADDRPOINTER_REG_17__SCAN_IN ^ n26093;
  assign n41025 = P1_PHYADDRPOINTER_REG_16__SCAN_IN ^ n26058;
  assign n40708 = P1_PHYADDRPOINTER_REG_15__SCAN_IN ^ n26030;
  assign n26578 = ~n26580 ^ P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n41131 = P1_PHYADDRPOINTER_REG_14__SCAN_IN ^ n25889;
  assign n40490 = P1_PHYADDRPOINTER_REG_13__SCAN_IN ^ n25885;
  assign n38389 = P1_PHYADDRPOINTER_REG_12__SCAN_IN ^ n25837;
  assign n39592 = P1_PHYADDRPOINTER_REG_11__SCAN_IN ^ n25061;
  assign n38804 = P1_PHYADDRPOINTER_REG_10__SCAN_IN ^ n25020;
  assign n36269 = n35820 ^ n35819;
  assign n24812 = ~n24811;
  assign n43442 = n40085 ^ n40084;
  assign n43569 = ~n42983 ^ n42982;
  assign n43042 = n42487 ^ P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n42817 = ~n43469 | ~P1_REIP_REG_27__SCAN_IN;
  assign n42935 = ~n43469 | ~P1_REIP_REG_26__SCAN_IN;
  assign n42934 = n28833 ^ n28832;
  assign n43329 = ~n42966 | ~n42925;
  assign n42834 = ~n43469 | ~P1_REIP_REG_24__SCAN_IN;
  assign n42172 = n28551 ^ n28550;
  assign n41743 = n26715 ^ n26714;
  assign n43330 = ~n28546 | ~n28545;
  assign n26148 = n26147 & n26146;
  assign n41022 = n26142 ^ n26141;
  assign n40798 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n40797 = ~n40088;
  assign n26571 = ~n43344 | ~n40706;
  assign n40098 = n25936 ^ n25935;
  assign n38662 = n25841 ^ n25840;
  assign n38643 = ~P1_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n35822 = n24193 ^ n28825;
  assign n36264 = n35832 ^ n35831;
  assign n35682 = ~n35111 | ~n35110;
  assign n34339 = n24187 ^ n28825;
  assign n34818 = ~n34340 & ~n34339;
  assign n35334 = ~n35333 | ~n35332;
  assign n33309 = n24181 ^ n28825;
  assign n33792 = ~n33310 & ~n33309;
  assign n36893 = ~n38650;
  assign n32532 = ~n24205 | ~n43033;
  assign n24339 = ~n24338;
  assign n39301 = ~n39942;
  assign n34725 = ~n34576 | ~n34575;
  assign n33718 = ~n32135 & ~n32134;
  assign n34258 = ~n24513 & ~n24512;
  assign n35180 = ~n35167 | ~n35166;
  assign n34748 = ~n34413 | ~n34412;
  assign n34421 = ~n34411 | ~n34410;
  assign n35351 = ~n34722 | ~n34721;
  assign n34090 = ~n34089 | ~n34088;
  assign n34088 = ~n34684 | ~n34270;
  assign n35089 = ~n35025 | ~n35024;
  assign n35033 = ~n35023 | ~n35022;
  assign n33726 = n33716 & n33715;
  assign n44106 = ~n35629 | ~n44098;
  assign n29579 = ~P1_STATE_REG_2__SCAN_IN;
  assign n23509 = ~n23508 | ~n23507;
  assign n26199 = ~n26489;
  assign n27871 = ~n27870;
  assign n43524 = ~n39571 ^ n39569;
  assign n41936 = ~n41935 | ~P2_EBX_REG_29__SCAN_IN;
  assign n41728 = ~n41935 | ~P2_EBX_REG_28__SCAN_IN;
  assign n43175 = n39764 ^ n39763;
  assign n42721 = n37469 ^ n37468;
  assign n42467 = n37274 ^ n37273;
  assign n28278 = ~n28277 | ~n28276;
  assign n40570 = n26478 ^ n26477;
  assign n41783 = ~n41617 ^ n41787;
  assign n41265 = ~n42953;
  assign n37831 = ~n37356 & ~n28269;
  assign n28269 = ~n37355;
  assign n28272 = ~n28271 | ~n28270;
  assign n35964 = ~n35599 & ~n35598;
  assign n36203 = ~n35964 | ~n35963;
  assign n35598 = ~n25745;
  assign n28227 = ~n28226;
  assign n25233 = ~n25232 | ~n25231;
  assign n35426 = ~n34917 & ~n34918;
  assign n34918 = ~n25731;
  assign n25176 = n25162 & n25161;
  assign n25173 = ~n25172 | ~n25171;
  assign n35253 = ~n25115 | ~n25114;
  assign n36248 = ~n25112 | ~n25111;
  assign n43056 = ~n43054;
  assign n43389 = n43393 ^ n43391;
  assign n43672 = n41725 ^ n41724;
  assign n41211 = ~n41725;
  assign n42799 = n43054 ^ n43055;
  assign n42909 = ~n28162 ^ n28163;
  assign n40053 = ~n39671 | ~n39670;
  assign n38014 = ~n37442 | ~n37441;
  assign n37121 = ~n37120 | ~n37119;
  assign n41703 = ~n32802 | ~n32801;
  assign n32217 = ~n25544 | ~n23415;
  assign n43777 = ~n43682;
  assign n28141 = ~P2_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n42354 = ~P2_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n42215 = ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n42658 = ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n42140 = ~n35971 ^ n35970;
  assign n42561 = ~n42624;
  assign n41702 = n41499 ^ n41498;
  assign n26519 = ~n26517;
  assign n33563 = ~n33585 ^ n26440;
  assign n43842 = n43837 ^ P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n43891 = ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n43743 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n43814 = n41941 ^ n41940;
  assign n43682 = ~n41733 ^ n41732;
  assign n43661 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n43645 = ~n41224 ^ n41223;
  assign n43315 = n43597 ^ P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n43316 = ~n43605 ^ n43603;
  assign n43317 = n40936 ^ n40935;
  assign n43155 = ~n43148 | ~n43160;
  assign n43154 = ~n43158 | ~n43153;
  assign n43582 = ~n39921 ^ n39920;
  assign n43581 = n43538 ^ n43537;
  assign n43537 = n43536 ^ P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n39761 = ~n39758;
  assign n43549 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n43223 = n43532 ^ n43211;
  assign n43211 = ~n43530 ^ P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n42953 = ~n40115 ^ n40114;
  assign n42952 = n43206 ^ n42908;
  assign n42906 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n42992 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n43015 = n39703 ^ n39702;
  assign n43018 = ~n43016 | ~n43583;
  assign n43014 = n42999 ^ n42998;
  assign n42998 = ~n42997 ^ n42996;
  assign n42855 = n42993 ^ n42722;
  assign n42722 = ~n42990 ^ n42992;
  assign n42871 = ~n37726 ^ n37725;
  assign n42874 = ~n42872 | ~n43583;
  assign n42870 = ~n42716 ^ n42464;
  assign n42598 = ~n42597 | ~n42596;
  assign n42628 = ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n42224 = ~n42221 | ~n42220;
  assign n42423 = n42213 ^ n42212;
  assign n42212 = ~n42211 | ~n42248;
  assign n42668 = ~n42666 | ~n42843;
  assign n42841 = n42664 ^ n42663;
  assign n42451 = n42307 ^ n42306;
  assign n28076 = n42062 ^ n27890;
  assign n41171 = n41490 ^ n41080;
  assign n27854 = ~n27853;
  assign n42600 = ~n43165;
  assign n39656 = ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n25576 = ~P2_STATE2_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n26546 = ~n23729;
  assign n36612 = ~n36486 ^ n36485;
  assign n35790 = n23683 ^ n26235;
  assign n43164 = ~n42110;
  assign n26211 = ~n26210 | ~n23415;
  assign n26210 = ~n26209 | ~n26208;
  assign n36500 = ~n24769 | ~n24768;
  assign n37945 = n32145 ^ n32144;
  assign n32893 = ~n32892;
  assign n32894 = ~n32891;
  assign n32509 = ~n26507;
  assign n37625 = ~n37624 | ~n39522;
  assign n37624 = ~n37623 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n37641 = ~n37640 | ~n37933;
  assign n37640 = ~n37654 | ~n39522;
  assign n38331 = ~n38330 | ~n39524;
  assign n38330 = ~n38329 | ~n39522;
  assign n39125 = ~n26374;
  assign n37858 = ~n37857 | ~n39524;
  assign n37857 = ~n37870 | ~n39522;
  assign n38212 = ~n37854;
  assign n37947 = ~n24781 & ~n24780;
  assign n38294 = ~n37076;
  assign n38297 = ~n38296 | ~n39522;
  assign n38614 = ~n38613 | ~n38929;
  assign n37953 = ~n37952 | ~n39524;
  assign n37952 = ~n37965 | ~n39522;
  assign n36634 = ~n36652;
  assign n37360 = ~n37359 | ~n39524;
  assign n37359 = ~n37376 | ~n39522;
  assign n37373 = ~n37609 | ~n37362;
  assign n39526 = ~n39525 | ~n39524;
  assign n41284 = ~n39601;
  assign n32966 = ~n29726 | ~n35452;
  assign n36161 = ~n35944 | ~n35943;
  assign n41518 = ~P3_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n34656 = ~n34655 | ~n41389;
  assign n32858 = ~n32866 | ~n32857;
  assign n32859 = ~n33500;
  assign n33124 = ~n33067 | ~n33066;
  assign n33622 = ~n33621 | ~n33620;
  assign n33514 = ~n33516 | ~n33496;
  assign n41389 = ~P3_EBX_REG_26__SCAN_IN;
  assign n32253 = ~P3_EBX_REG_0__SCAN_IN | ~P3_EBX_REG_1__SCAN_IN;
  assign n32472 = ~n30706;
  assign n34011 = ~P3_EAX_REG_21__SCAN_IN | ~n34013;
  assign n35307 = ~P3_EAX_REG_14__SCAN_IN | ~n35695;
  assign n32826 = ~n27656;
  assign n32284 = ~n27281 & ~n27280;
  assign n27315 = ~n27298 | ~n27297;
  assign n41399 = ~n27746 ^ P3_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n41091 = ~n28762 ^ P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n40859 = ~n41147 | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n41156 = ~n41158 ^ n35529;
  assign n40732 = ~n41093;
  assign n41100 = ~P3_STATE2_REG_0__SCAN_IN & ~n40527;
  assign n41233 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n40817 = ~n42321 ^ n38924;
  assign n40410 = ~n39394 | ~n40470;
  assign n40335 = n37710 ^ n37709;
  assign n36869 = ~n40743 | ~n39388;
  assign n32881 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN | ~P3_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n36195 = ~n36194 | ~n36193;
  assign n36439 = ~P3_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n36433 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN | ~P3_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n36444 = ~n36427 | ~n41147;
  assign n36446 = ~n36429 | ~n36428;
  assign n40371 = ~n27348 & ~n36078;
  assign n36927 = ~n27336 ^ n27335;
  assign n36913 = n27677 ^ n27676;
  assign n36659 = ~n36661 & ~n33945;
  assign n27282 = ~n32284;
  assign n27653 = ~n27652 | ~n28088;
  assign n27654 = ~n27635 | ~n27634;
  assign n41535 = ~n40125;
  assign n41556 = n40752 ^ P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n40836 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~n40835;
  assign n41011 = n39422 ^ n39421;
  assign n39796 = ~n38151 ^ P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n40532 = ~n38174 ^ n40531;
  assign n40466 = ~n37574 ^ P3_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n40425 = ~n40475 | ~n40416;
  assign n40408 = ~n38030 ^ n40431;
  assign n39444 = ~n39443 | ~n39442;
  assign n39412 = ~n39409 | ~n39408;
  assign n39409 = ~n39403 | ~n39442;
  assign n41240 = ~n41546;
  assign n40398 = ~n40397 | ~n40964;
  assign n40981 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n40200 = ~n40192 | ~n40196;
  assign n27593 = ~n27747;
  assign n40182 = ~n40179 | ~n40194;
  assign n40179 = ~n40191 | ~n40270;
  assign n38605 = ~n38604 | ~n38603;
  assign n27810 = ~n27803 | ~n31787;
  assign n27786 = ~n27783 | ~n32475;
  assign n43990 = ~n29726 | ~P3_STATEBS16_REG_SCAN_IN;
  assign n41354 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n36055 = ~n40422 | ~n36054;
  assign n36052 = ~n29442;
  assign n42016 = ~n41375 | ~n40527;
  assign n42013 = ~n41670;
  assign n31442 = n39315 & n33714;
  assign n43800 = ~n43799 | ~n43798;
  assign n43384 = ~n43375 | ~n43374;
  assign n42166 = ~n42159 | ~n42158;
  assign n43343 = n28662 ^ n28661;
  assign n41854 = ~n41853 | ~n41852;
  assign n41904 = ~n41903 | ~n41902;
  assign n26708 = ~n26701 | ~n26700;
  assign n40718 = ~n43803 | ~n40706;
  assign n40715 = ~n40714 | ~n40713;
  assign n41140 = ~n43803 | ~n41127;
  assign n26078 = ~n26077 | ~n26076;
  assign n26081 = ~n43803 | ~n40098;
  assign n38792 = ~n39593 | ~n41453;
  assign n37519 = ~n37518 | ~n37517;
  assign n37507 = ~n37239 | ~n37238;
  assign n43570 = ~n43803;
  assign n35515 = ~n35514 | ~n35513;
  assign n43796 = ~n26070 & ~n26069;
  assign n28046 = ~n28525;
  assign n40493 = ~n25850 ^ n25849;
  assign n38636 = ~n38388;
  assign n44007 = ~n38807;
  assign n37550 = ~n36903 | ~n36902;
  assign n34815 = ~n34814 | ~n34813;
  assign n42028 = ~n43031;
  assign n41425 = ~n42505;
  assign n41039 = ~n41953;
  assign n40549 = ~n41194;
  assign n41130 = n26085 ^ n26084;
  assign n32233 = ~n32232 | ~n32231;
  assign n44092 = ~n44028 & ~n44093;
  assign n31748 = ~n32107 | ~n42736;
  assign n31757 = ~n32107 | ~n43121;
  assign n42371 = ~n28848 ^ n28497;
  assign n28497 = ~n43462 ^ P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n28549 = ~n28510 ^ P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n28483 = ~n43462 ^ P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n41742 = n28477 ^ n27827;
  assign n40802 = n27822 ^ n26584;
  assign n40692 = ~n26579 ^ n26578;
  assign n40486 = ~n40097 ^ n40096;
  assign n39643 = n39590 ^ n39589;
  assign n39594 = ~n39593 | ~n43367;
  assign n37516 = P1_PHYADDRPOINTER_REG_9__SCAN_IN ^ n24981;
  assign n37501 = ~n37551 | ~n43367;
  assign n37502 = ~n37498 | ~n43707;
  assign n37243 = P1_PHYADDRPOINTER_REG_8__SCAN_IN ^ n24944;
  assign n37003 = ~n43707 | ~n37000;
  assign n37002 = ~n37001 | ~n43367;
  assign n36993 = ~n36269;
  assign n35681 = P1_PHYADDRPOINTER_REG_6__SCAN_IN ^ n24861;
  assign n36110 = n24844 ^ n24852;
  assign n35518 = P1_PHYADDRPOINTER_REG_4__SCAN_IN ^ n24843;
  assign n42829 = ~n42676 | ~n42369;
  assign n41749 = ~n41965 | ~P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n41279 = ~n41278 | ~n41277;
  assign n41278 = ~n43344 | ~n41276;
  assign n40805 = ~n40804 | ~n40803;
  assign n40804 = ~n43344 | ~n41022;
  assign n25986 = ~n25985 | ~n40786;
  assign n25985 = ~n43344 | ~n41127;
  assign n39563 = ~n43344 | ~n44008;
  assign n24203 = ~n24202 | ~n31449;
  assign n32340 = ~n31915 | ~n31914;
  assign n39964 = ~P1_INSTQUEUE_REG_0__0__SCAN_IN | ~n40041;
  assign n39975 = ~P1_INSTQUEUE_REG_0__1__SCAN_IN | ~n40041;
  assign n40008 = ~P1_INSTQUEUE_REG_0__2__SCAN_IN | ~n40041;
  assign n39997 = ~P1_INSTQUEUE_REG_0__3__SCAN_IN | ~n40041;
  assign n39986 = ~P1_INSTQUEUE_REG_0__4__SCAN_IN | ~n40041;
  assign n40045 = ~P1_INSTQUEUE_REG_0__5__SCAN_IN | ~n40041;
  assign n40030 = ~P1_INSTQUEUE_REG_0__6__SCAN_IN | ~n40041;
  assign n40019 = ~P1_INSTQUEUE_REG_0__7__SCAN_IN | ~n40041;
  assign n39076 = ~P1_INSTQUEUE_REG_2__0__SCAN_IN | ~n39101;
  assign n39068 = ~P1_INSTQUEUE_REG_2__1__SCAN_IN | ~n39101;
  assign n39084 = ~P1_INSTQUEUE_REG_2__2__SCAN_IN | ~n39101;
  assign n39044 = ~P1_INSTQUEUE_REG_2__3__SCAN_IN | ~n39101;
  assign n39052 = ~P1_INSTQUEUE_REG_2__4__SCAN_IN | ~n39101;
  assign n39060 = ~P1_INSTQUEUE_REG_2__5__SCAN_IN | ~n39101;
  assign n39104 = ~P1_INSTQUEUE_REG_2__6__SCAN_IN | ~n39101;
  assign n39092 = ~P1_INSTQUEUE_REG_2__7__SCAN_IN | ~n39101;
  assign n38446 = ~n39962 | ~n38473;
  assign n38447 = ~P1_INSTQUEUE_REG_4__0__SCAN_IN | ~n38472;
  assign n38438 = ~n39973 | ~n38473;
  assign n38439 = ~P1_INSTQUEUE_REG_4__1__SCAN_IN | ~n38472;
  assign n38474 = ~n40006 | ~n38473;
  assign n38475 = ~P1_INSTQUEUE_REG_4__2__SCAN_IN | ~n38472;
  assign n38462 = ~n39995 | ~n38473;
  assign n38463 = ~P1_INSTQUEUE_REG_4__3__SCAN_IN | ~n38472;
  assign n38422 = ~n39984 | ~n38473;
  assign n38423 = ~P1_INSTQUEUE_REG_4__4__SCAN_IN | ~n38472;
  assign n38430 = ~n40043 | ~n38473;
  assign n38431 = ~P1_INSTQUEUE_REG_4__5__SCAN_IN | ~n38472;
  assign n38414 = ~n40028 | ~n38473;
  assign n38415 = ~P1_INSTQUEUE_REG_4__6__SCAN_IN | ~n38472;
  assign n38454 = ~n40017 | ~n38473;
  assign n38455 = ~P1_INSTQUEUE_REG_4__7__SCAN_IN | ~n38472;
  assign n38531 = ~P1_INSTQUEUE_REG_6__0__SCAN_IN | ~n38556;
  assign n38523 = ~P1_INSTQUEUE_REG_6__1__SCAN_IN | ~n38556;
  assign n38539 = ~P1_INSTQUEUE_REG_6__2__SCAN_IN | ~n38556;
  assign n38507 = ~P1_INSTQUEUE_REG_6__3__SCAN_IN | ~n38556;
  assign n38547 = ~P1_INSTQUEUE_REG_6__4__SCAN_IN | ~n38556;
  assign n38515 = ~P1_INSTQUEUE_REG_6__5__SCAN_IN | ~n38556;
  assign n38559 = ~P1_INSTQUEUE_REG_6__6__SCAN_IN | ~n38556;
  assign n38499 = ~P1_INSTQUEUE_REG_6__7__SCAN_IN | ~n38556;
  assign n34730 = ~n34729 | ~n34728;
  assign n39328 = ~P1_INSTQUEUE_REG_8__0__SCAN_IN | ~n39377;
  assign n39360 = ~P1_INSTQUEUE_REG_8__1__SCAN_IN | ~n39377;
  assign n39344 = ~P1_INSTQUEUE_REG_8__2__SCAN_IN | ~n39377;
  assign n39336 = ~P1_INSTQUEUE_REG_8__3__SCAN_IN | ~n39377;
  assign n39352 = ~P1_INSTQUEUE_REG_8__4__SCAN_IN | ~n39377;
  assign n39368 = ~P1_INSTQUEUE_REG_8__5__SCAN_IN | ~n39377;
  assign n39380 = ~P1_INSTQUEUE_REG_8__6__SCAN_IN | ~n39377;
  assign n39320 = ~P1_INSTQUEUE_REG_8__7__SCAN_IN | ~n39377;
  assign n38108 = ~n39962 | ~n38127;
  assign n38109 = ~P1_INSTQUEUE_REG_10__0__SCAN_IN | ~n38126;
  assign n38068 = ~n39973 | ~n38127;
  assign n38069 = ~P1_INSTQUEUE_REG_10__1__SCAN_IN | ~n38126;
  assign n38100 = ~n40006 | ~n38127;
  assign n38101 = ~P1_INSTQUEUE_REG_10__2__SCAN_IN | ~n38126;
  assign n38116 = ~n39995 | ~n38127;
  assign n38117 = ~P1_INSTQUEUE_REG_10__3__SCAN_IN | ~n38126;
  assign n38084 = ~n39984 | ~n38127;
  assign n38085 = ~P1_INSTQUEUE_REG_10__4__SCAN_IN | ~n38126;
  assign n38092 = ~n40043 | ~n38127;
  assign n38093 = ~P1_INSTQUEUE_REG_10__5__SCAN_IN | ~n38126;
  assign n38076 = ~n40028 | ~n38127;
  assign n38077 = ~P1_INSTQUEUE_REG_10__6__SCAN_IN | ~n38126;
  assign n38128 = ~n40017 | ~n38127;
  assign n38129 = ~P1_INSTQUEUE_REG_10__7__SCAN_IN | ~n38126;
  assign n39873 = ~P1_INSTQUEUE_REG_12__0__SCAN_IN | ~n39882;
  assign n39865 = ~P1_INSTQUEUE_REG_12__1__SCAN_IN | ~n39882;
  assign n39833 = ~P1_INSTQUEUE_REG_12__2__SCAN_IN | ~n39882;
  assign n39885 = ~P1_INSTQUEUE_REG_12__3__SCAN_IN | ~n39882;
  assign n39825 = ~P1_INSTQUEUE_REG_12__4__SCAN_IN | ~n39882;
  assign n39849 = ~P1_INSTQUEUE_REG_12__5__SCAN_IN | ~n39882;
  assign n39857 = ~P1_INSTQUEUE_REG_12__6__SCAN_IN | ~n39882;
  assign n39841 = ~P1_INSTQUEUE_REG_12__7__SCAN_IN | ~n39882;
  assign n38855 = ~P1_INSTQUEUE_REG_14__1__SCAN_IN | ~n38888;
  assign n38863 = ~P1_INSTQUEUE_REG_14__2__SCAN_IN | ~n38888;
  assign n38847 = ~P1_INSTQUEUE_REG_14__3__SCAN_IN | ~n38888;
  assign n38839 = ~P1_INSTQUEUE_REG_14__4__SCAN_IN | ~n38888;
  assign n38891 = ~P1_INSTQUEUE_REG_14__5__SCAN_IN | ~n38888;
  assign n38879 = ~P1_INSTQUEUE_REG_14__6__SCAN_IN | ~n38888;
  assign n38871 = ~P1_INSTQUEUE_REG_14__7__SCAN_IN | ~n38888;
  assign n29568 = ~n24509;
  assign n44000 = ~n23712 | ~n31522;
  assign n28151 = ~n31771;
  assign n29550 = ~P2_REIP_REG_1__SCAN_IN;
  assign n41916 = ~n41913 | ~n43808;
  assign n28148 = ~n41916 | ~n41718;
  assign n28222 = ~n28221 | ~n28220;
  assign n41737 = ~n41723 | ~n41722;
  assign n40933 = ~n40932 | ~n40931;
  assign n37470 = ~n42721 | ~n41934;
  assign n37461 = ~n42857;
  assign n37275 = ~n42467 | ~n41934;
  assign n37267 = ~n37266 | ~n41942;
  assign n42352 = n37736 ^ n37735;
  assign n37731 = ~P2_EBX_REG_19__SCAN_IN | ~n41935;
  assign n37730 = ~n37724 | ~n37723;
  assign n40687 = ~n40686 | ~n40685;
  assign n42452 = n35602 ^ n35601;
  assign n40663 = ~n40662 | ~n40661;
  assign n39491 = ~n39487 | ~n40668;
  assign n39470 = ~n39466 | ~n40668;
  assign n37338 = ~n37334 | ~n40668;
  assign n40367 = ~n40361 | ~n40360;
  assign n38833 = ~n38827 | ~n38826;
  assign n40579 = n37289 & n37288;
  assign n40324 = ~n40318 | ~n40317;
  assign n28368 = ~n37288;
  assign n43633 = n43476 ^ n43475;
  assign n41755 = n41785 ^ n41783;
  assign n26911 = ~n26908;
  assign n40069 = ~n43015 | ~n43525;
  assign n42616 = n37831 ^ n37830;
  assign n42842 = ~n36206 ^ n36205;
  assign n42565 = n35432 ^ n35431;
  assign n35599 = ~n35426 | ~n35425;
  assign n34917 = ~n34646 | ~n34645;
  assign n40580 = ~n36249 ^ n36248;
  assign n40325 = ~n37638;
  assign n43130 = n43390 ^ n43389;
  assign n41842 = n42746 ^ n42745;
  assign n41675 = n41656 ^ n41786;
  assign n40067 = n40053 ^ n40052;
  assign n40298 = ~n32798 ^ n28079;
  assign n25097 = ~n25095 | ~n25094;
  assign n36958 = ~n36957 | ~n36956;
  assign n36957 = ~n36954 | ~n36953;
  assign n36011 = ~n36010 | ~n36009;
  assign n31353 = ~n31344 & ~n31202;
  assign n43912 = P2_PHYADDRPOINTER_REG_31__SCAN_IN ^ n24765;
  assign n43808 = ~n28146 ^ n28145;
  assign n43013 = ~n42989 ^ P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n42709 = ~n42989;
  assign n42431 = ~n42428 | ~n42427;
  assign n42059 = ~n42058;
  assign n42076 = ~n42564 | ~n43913;
  assign n41170 = ~n41077 ^ n41076;
  assign n38379 = ~n38378 | ~n38377;
  assign n38377 = ~n39667 | ~n43809;
  assign n37556 = n36861 ^ P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n36493 = ~n36492 | ~n36491;
  assign n36492 = ~n36613 | ~n43913;
  assign n43812 = ~n43827 ^ n43754;
  assign n43754 = ~n43828 ^ P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n43776 = ~n43750 ^ n43671;
  assign n43775 = n43746 ^ P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n43644 = n43610 ^ n43661;
  assign n43578 = ~n43549 & ~n43156;
  assign n43156 = ~n43187 | ~n43617;
  assign n43222 = n43550 ^ n43549;
  assign n42894 = ~n42704 | ~n42703;
  assign n42520 = ~n42519 | ~n42518;
  assign n42519 = ~n42517 | ~n43583;
  assign n42868 = ~n42527 | ~n42526;
  assign n42282 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n42289 = ~n42288 | ~n42440;
  assign n42560 = ~n41698 | ~n28071;
  assign n41697 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n40941 = n40759 ^ n40758;
  assign n40758 = ~n40757 ^ P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n28061 = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n40769 = ~n40767 | ~n28061;
  assign n39651 = ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n36862 = ~n43893 & ~n37556;
  assign n36616 = ~n36615 | ~n36614;
  assign n36615 = ~n36613 | ~n43876;
  assign n34913 = ~n34914;
  assign n36532 = ~n31055 | ~n39522;
  assign n37782 = ~n37839 | ~n38706;
  assign n37739 = ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n37799 = ~n37839 | ~n38669;
  assign n37840 = ~n37839 | ~n38678;
  assign n37817 = ~n37839 | ~n38687;
  assign n37790 = ~n37839 | ~n38696;
  assign n37809 = ~n37839 | ~n37808;
  assign n36940 = ~n36939 | ~n36938;
  assign n36680 = ~n36679 | ~n36678;
  assign n37596 = ~n37610 | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n37648 = ~n37647 | ~n37646;
  assign n37939 = ~n37938 | ~n37937;
  assign n38567 = ~n38566 | ~n38565;
  assign n38565 = ~P2_INSTQUEUE_REG_4__0__SCAN_IN | ~n39612;
  assign n38357 = ~n38356 | ~n38355;
  assign n38356 = ~P2_INSTQUEUE_REG_4__1__SCAN_IN | ~n39612;
  assign n38341 = ~n38340 | ~n38339;
  assign n38340 = ~P2_INSTQUEUE_REG_4__2__SCAN_IN | ~n39612;
  assign n38349 = ~n38348 | ~n38347;
  assign n38348 = ~P2_INSTQUEUE_REG_4__3__SCAN_IN | ~n39612;
  assign n38581 = ~P2_INSTQUEUE_REG_4__4__SCAN_IN | ~n39612;
  assign n38575 = ~n38574 | ~n38573;
  assign n38573 = ~P2_INSTQUEUE_REG_4__5__SCAN_IN | ~n39612;
  assign n38365 = ~n38364 | ~n38363;
  assign n38364 = ~P2_INSTQUEUE_REG_4__6__SCAN_IN | ~n39612;
  assign n37150 = ~n37149 | ~n37148;
  assign n37209 = ~n37208 | ~n37207;
  assign n37198 = ~n37197 | ~n37196;
  assign n37174 = ~n37173 | ~n37172;
  assign n37158 = ~n37157 | ~n37156;
  assign n37182 = ~n37181 | ~n37180;
  assign n37166 = ~n37165 | ~n37164;
  assign n37190 = ~n37189 | ~n37188;
  assign n39147 = ~n39193 | ~n39542;
  assign n39173 = ~n39193 | ~n39233;
  assign n39165 = ~n39193 | ~n39285;
  assign n39139 = ~n39193 | ~n39271;
  assign n39157 = ~n39193 | ~n39156;
  assign n39181 = ~n39193 | ~n39201;
  assign n39194 = ~n39193 | ~n39606;
  assign n37048 = ~n37047 | ~n37046;
  assign n37081 = ~n37080 | ~n37079;
  assign n37064 = ~n37063 | ~n37062;
  assign n37072 = ~n37071 | ~n37070;
  assign n37056 = ~n37055 | ~n37054;
  assign n39203 = ~n39286 | ~n39201;
  assign n38709 = ~n38708 | ~n38707;
  assign n38718 = ~n38717 | ~n38716;
  assign n38672 = ~n38671 | ~n38670;
  assign n38681 = ~n38680 | ~n38679;
  assign n38690 = ~n38689 | ~n38688;
  assign n38929 = ~n38627;
  assign n38699 = ~n38698 | ~n38697;
  assign n37976 = ~P2_INSTQUEUE_REG_12__0__SCAN_IN | ~n38313;
  assign n37957 = ~P2_INSTQUEUE_REG_12__1__SCAN_IN | ~n38313;
  assign n38008 = ~P2_INSTQUEUE_REG_12__2__SCAN_IN | ~n38313;
  assign n37992 = ~P2_INSTQUEUE_REG_12__3__SCAN_IN | ~n38313;
  assign n38000 = ~P2_INSTQUEUE_REG_12__5__SCAN_IN | ~n38313;
  assign n38304 = ~n37944 | ~n39114;
  assign n37984 = ~P2_INSTQUEUE_REG_12__7__SCAN_IN | ~n38313;
  assign n36729 = ~n36728 | ~n36727;
  assign n36808 = ~n36807 | ~n36806;
  assign n36788 = ~n36787 | ~n36786;
  assign n36705 = ~n36704 | ~n36703;
  assign n36697 = ~n36696 | ~n36695;
  assign n36796 = ~n37944 | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n36713 = ~n36712 | ~n36711;
  assign n37368 = ~P2_INSTQUEUE_REG_14__0__SCAN_IN | ~n38778;
  assign n37392 = ~P2_INSTQUEUE_REG_14__1__SCAN_IN | ~n38778;
  assign n37384 = ~P2_INSTQUEUE_REG_14__5__SCAN_IN | ~n38778;
  assign n38769 = ~n37375;
  assign n41314 = ~n41313 | ~n41312;
  assign n38814 = ~P2_REIP_REG_3__SCAN_IN;
  assign n29204 = ~P2_REIP_REG_9__SCAN_IN;
  assign n29221 = ~P2_REIP_REG_13__SCAN_IN;
  assign n41365 = ~n31675 | ~n31674;
  assign n36168 = ~n36160 | ~n36159;
  assign n35644 = ~n35525 | ~n35949;
  assign n34545 = ~n33951;
  assign n33756 = ~n35525 | ~n33514;
  assign n35525 = ~n35951;
  assign n41864 = ~P3_EBX_REG_29__SCAN_IN | ~n43930;
  assign n41681 = ~P3_EBX_REG_28__SCAN_IN | ~n43930;
  assign n41863 = ~n41865;
  assign n34400 = ~P3_EBX_REG_14__SCAN_IN;
  assign n43933 = ~n43930 | ~n33162;
  assign n42135 = ~n32526 & ~n32672;
  assign n41059 = ~n42052;
  assign n36281 = ~n36243 | ~n36283;
  assign n33062 = ~n32986 | ~n32985;
  assign n32501 = n27112 | n27111;
  assign n33095 = ~n27659;
  assign n32193 = ~n43982;
  assign n43984 = ~n32190 & ~n32156;
  assign n41532 = n28100 ^ P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n41118 = ~n41514;
  assign n41111 = ~n41110 | ~n41109;
  assign n40848 = ~n41168;
  assign n40815 = ~n42321 ^ n38923;
  assign n37024 = ~n38142 | ~n40421;
  assign n36868 = ~n40744 | ~n39387;
  assign n36479 = ~n36456 | ~n36455;
  assign n36963 = ~P3_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n36978 = ~n36977 | ~n36976;
  assign n41259 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n41002 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n40254 = ~n40241 | ~n40820;
  assign n40531 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n40484 = ~n41145 | ~P3_REIP_REG_20__SCAN_IN;
  assign n40431 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n40421 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n40344 = ~n40337 | ~n40336;
  assign n40231 = ~n40228 | ~n40227;
  assign n40146 = ~n40143 | ~n40142;
  assign n40142 = ~n40141 | ~n40140;
  assign n40973 = ~n40963 | ~n40962;
  assign n40515 = ~n40512 | ~n40511;
  assign n40459 = ~n40457 | ~n40456;
  assign n39633 = ~n39632 | ~n39631;
  assign n39620 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n40191 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n38731 = ~n38730 & ~n38729;
  assign n36352 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n40418 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n29449 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n43992 = ~P3_STATE2_REG_3__SCAN_IN;
  assign n43577 = ~n43563 & ~n43562;
  assign n28896 = ~n28884 | ~n28883;
  assign n28880 = ~n28879 | ~n28878;
  assign n28845 = ~n29632 & ~n28844;
  assign n28844 = ~n35512 | ~n28876;
  assign n28538 = ~n28521 | ~n28520;
  assign n42191 = ~P1_REIP_REG_22__SCAN_IN | ~n42171;
  assign n27851 = ~n27839 | ~n27838;
  assign n36116 = ~n36106 | ~n36105;
  assign n35891 = ~n35888 & ~n35887;
  assign n36150 = ~n36140 | ~n36139;
  assign n28826 = ~n44023 | ~P1_EBX_REG_29__SCAN_IN;
  assign n28724 = ~n44023 | ~P1_EBX_REG_28__SCAN_IN;
  assign n28672 = ~n44023 | ~P1_EBX_REG_27__SCAN_IN;
  assign n41442 = n41441 & n41440;
  assign n26694 = ~n26693 | ~n26692;
  assign n26718 = ~n26717 | ~n26716;
  assign n26151 = ~n26150 | ~n26149;
  assign n26039 = ~n26038 | ~n26037;
  assign n25948 = ~n25947 | ~n25946;
  assign n37537 = ~n39593 | ~n43297;
  assign n43741 = ~n43740 | ~n43739;
  assign n39936 = ~n39933 | ~n39932;
  assign n37825 = ~n32242 | ~n39593;
  assign n43365 = ~n43364 | ~n43363;
  assign n43141 = ~n43140 | ~n43139;
  assign n42820 = ~n42819 | ~n42818;
  assign n43038 = ~n43037 | ~n43036;
  assign n42510 = ~n42509 | ~n42508;
  assign n41958 = ~n41957 | ~n41956;
  assign n38396 = ~n38659 | ~n43707;
  assign n35687 = ~n35686 | ~n35685;
  assign n42988 = ~n42970 | ~n42969;
  assign n42556 = ~n42542 | ~n43437;
  assign n26575 = ~n40793 | ~P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n35838 = ~n35837 & ~n35836;
  assign n37494 = ~P1_INSTQUEUE_REG_14__0__SCAN_IN | ~n38888;
  assign n34524 = ~n34522 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n34522 = ~n44098 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n39929 = ~n41934 | ~n43171;
  assign n39770 = ~n39755 & ~n39754;
  assign n40119 = ~n40113 | ~n40112;
  assign n39708 = ~n39699 | ~n39698;
  assign n36398 = ~n36397 | ~n41942;
  assign n39228 = ~n39227 & ~n39226;
  assign n40641 = ~n40640 | ~n40639;
  assign n40598 = ~n40597 | ~n40596;
  assign n40618 = ~n40617 | ~n40616;
  assign n39583 = ~n43916;
  assign n39716 = ~n39715 | ~n39714;
  assign n39296 = ~n39295 | ~n39294;
  assign n39297 = ~n39293 | ~n43523;
  assign n38138 = ~n38137 | ~n38136;
  assign n38139 = ~n38135 | ~n43523;
  assign n38982 = ~n39293 | ~n43693;
  assign n38028 = ~n38135 | ~n43693;
  assign n33424 = ~n33548 | ~P2_LWORD_REG_13__SCAN_IN;
  assign n33428 = ~n33548 | ~P2_LWORD_REG_12__SCAN_IN;
  assign n33432 = ~n33548 | ~P2_LWORD_REG_11__SCAN_IN;
  assign n33436 = ~n33548 | ~P2_LWORD_REG_10__SCAN_IN;
  assign n33440 = ~n33548 | ~P2_LWORD_REG_9__SCAN_IN;
  assign n33444 = ~n33548 | ~P2_LWORD_REG_8__SCAN_IN;
  assign n33448 = ~n33548 | ~P2_LWORD_REG_7__SCAN_IN;
  assign n33452 = ~n33548 | ~P2_LWORD_REG_6__SCAN_IN;
  assign n33456 = ~n33548 | ~P2_LWORD_REG_5__SCAN_IN;
  assign n33460 = ~n33548 | ~P2_LWORD_REG_4__SCAN_IN;
  assign n33477 = ~n33548 | ~P2_LWORD_REG_3__SCAN_IN;
  assign n33464 = ~n33548 | ~P2_LWORD_REG_2__SCAN_IN;
  assign n33468 = ~n33548 | ~P2_LWORD_REG_1__SCAN_IN;
  assign n33472 = ~n33548 | ~P2_LWORD_REG_0__SCAN_IN;
  assign n43909 = ~n43908 & ~n43907;
  assign n42479 = ~n42478 | ~n42477;
  assign n42446 = n42445 & n42444;
  assign n42268 = ~n42267 | ~n42266;
  assign n42396 = ~n42395 | ~n42394;
  assign n42149 = ~n42148 | ~n42147;
  assign n40164 = ~n40163 | ~n40162;
  assign n42125 = ~n42124 | ~n42648;
  assign n39668 = ~n39667 | ~n43748;
  assign n37605 = ~P2_INSTQUEUE_REG_1__4__SCAN_IN | ~n37604;
  assign n37529 = ~P2_INSTQUEUE_REG_1__6__SCAN_IN | ~n37604;
  assign n37917 = ~n37915 & ~n37914;
  assign n37909 = ~n37907 & ~n37906;
  assign n39613 = ~P2_INSTQUEUE_REG_4__7__SCAN_IN | ~n39612;
  assign n37549 = ~n37546 & ~n37545;
  assign n37433 = ~n37431 & ~n37430;
  assign n37414 = ~P2_INSTQUEUE_REG_9__1__SCAN_IN | ~n37423;
  assign n37424 = ~P2_INSTQUEUE_REG_9__2__SCAN_IN | ~n37423;
  assign n37406 = ~P2_INSTQUEUE_REG_9__7__SCAN_IN | ~n37423;
  assign n38939 = ~P2_INSTQUEUE_REG_11__0__SCAN_IN | ~n38938;
  assign n38635 = ~n38624 & ~n38623;
  assign n38314 = ~P2_INSTQUEUE_REG_12__4__SCAN_IN | ~n38313;
  assign n38275 = ~P2_INSTQUEUE_REG_12__6__SCAN_IN | ~n38313;
  assign n38751 = ~P2_INSTQUEUE_REG_14__2__SCAN_IN | ~n38778;
  assign n38743 = ~P2_INSTQUEUE_REG_14__3__SCAN_IN | ~n38778;
  assign n38779 = ~P2_INSTQUEUE_REG_14__4__SCAN_IN | ~n38778;
  assign n38759 = ~P2_INSTQUEUE_REG_14__6__SCAN_IN | ~n38778;
  assign n38767 = ~P2_INSTQUEUE_REG_14__7__SCAN_IN | ~n38778;
  assign n40916 = ~P2_INSTQUEUE_REG_15__2__SCAN_IN | ~n41309;
  assign n40904 = ~P2_INSTQUEUE_REG_15__3__SCAN_IN | ~n41309;
  assign n40892 = ~P2_INSTQUEUE_REG_15__5__SCAN_IN | ~n41309;
  assign n40893 = ~n40890 & ~n40889;
  assign n41306 = ~n41300 & ~n41299;
  assign n41294 = ~n41288 & ~n41287;
  assign n35781 = ~n35816 | ~P2_STATE2_REG_3__SCAN_IN;
  assign n35958 = ~n35957 | ~n35956;
  assign n35660 = ~n35659 | ~n35940;
  assign n40546 = ~n40543 | ~n40545;
  assign n39744 = ~n39742 | ~n39741;
  assign n39504 = ~n39501 | ~n39503;
  assign n37922 = ~n37920 | ~n37919;
  assign n37327 = ~n37326 | ~n37919;
  assign n36405 = ~n36404 | ~n37325;
  assign n36179 = ~n36178 | ~n36401;
  assign n35555 = ~n35554 | ~n36177;
  assign n41421 = ~P3_PHYADDRPOINTER_REG_31__SCAN_IN | ~n41420;
  assign n41167 = ~n42341;
  assign n39438 = ~n40747 | ~n41002;
  assign n37778 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~n37777;
  assign n37777 = ~n37776 | ~n37775;
  assign n38169 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~n38188;
  assign n38189 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN | ~n38188;
  assign n37594 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN | ~n38047;
  assign n38048 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN | ~n38047;
  assign n36887 = ~n39410 | ~n40857;
  assign n36673 = ~n36672 | ~n36671;
  assign n27820 = ~n27819 | ~n41410;
  assign n28105 = ~n28104 | ~n41527;
  assign n28771 = ~n28770 | ~n41104;
  assign n40986 = ~n41257 | ~n40985;
  assign n38610 = ~n38609 | ~n41257;
  assign n42026 = ~n42025 | ~n42024;
  assign U215 = P2_ADDRESS_REG_29__SCAN_IN | n23017;
  assign n27152 = ~n36320;
  assign n28191 = ~n43061 & ~P2_STATE2_REG_3__SCAN_IN;
  assign n22929 = n23846 & n23845;
  assign n22930 = n24217 & n24727;
  assign n22931 = n23414 & n23413;
  assign n22932 = n24220 & n24219;
  assign n43540 = ~n43917;
  assign n23127 = ~n43061;
  assign n22934 = ~n29580 | ~n29579;
  assign n34812 = ~n34814 & ~n34813;
  assign n22935 = n32672 | n32860;
  assign n22936 = n33487 | n27604;
  assign n22937 = n27346 | n27345;
  assign n27697 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n34858 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n26859 = ~n26808;
  assign n28062 = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n26522 = ~P2_REIP_REG_4__SCAN_IN;
  assign n28316 = ~P2_REIP_REG_24__SCAN_IN;
  assign n22938 = n25887 | n25886;
  assign n22939 = n26441 | n23322;
  assign n22940 = n23887 & n23886;
  assign n22941 = n23351 & n23350;
  assign n23758 = ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n27696 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n22942 = n24874 | n24873;
  assign n25556 = ~n25758;
  assign n25758 = ~n25494 & ~n23322;
  assign n26849 = ~n26789;
  assign n28236 = ~P2_REIP_REG_12__SCAN_IN;
  assign n24862 = ~P1_EAX_REG_7__SCAN_IN;
  assign n28249 = ~P2_REIP_REG_14__SCAN_IN;
  assign n29669 = ~P1_REIP_REG_31__SCAN_IN;
  assign n28229 = ~P2_REIP_REG_11__SCAN_IN;
  assign n28331 = ~P2_REIP_REG_26__SCAN_IN;
  assign n25724 = ~P2_EAX_REG_9__SCAN_IN;
  assign n22943 = n23402 & n23401;
  assign n35543 = ~P3_REIP_REG_28__SCAN_IN;
  assign n33191 = ~n35392;
  assign n24804 = ~P1_EAX_REG_0__SCAN_IN;
  assign n28345 = ~P2_REIP_REG_28__SCAN_IN;
  assign n26537 = ~P2_REIP_REG_6__SCAN_IN;
  assign n27915 = ~P2_REIP_REG_10__SCAN_IN;
  assign n29493 = ~P2_REIP_REG_19__SCAN_IN;
  assign n29749 = ~NA;
  assign n24818 = ~P1_EAX_REG_3__SCAN_IN;
  assign n24788 = ~P1_EAX_REG_2__SCAN_IN;
  assign n29506 = ~P2_REIP_REG_17__SCAN_IN;
  assign n28324 = ~P2_REIP_REG_25__SCAN_IN;
  assign n23636 = ~P2_REIP_REG_2__SCAN_IN;
  assign n28262 = ~P2_REIP_REG_16__SCAN_IN;
  assign n27901 = ~P2_REIP_REG_8__SCAN_IN;
  assign n26530 = ~P2_REIP_REG_5__SCAN_IN;
  assign n25671 = ~P2_EAX_REG_6__SCAN_IN;
  assign n25738 = ~P2_EAX_REG_11__SCAN_IN;
  assign n29462 = ~n29226;
  assign n22945 = n24948 | n24947;
  assign n28289 = ~P2_REIP_REG_20__SCAN_IN;
  assign n43850 = ~n43879;
  assign n25583 = ~n25574 & ~n25573;
  assign n24283 = ~P1_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n24537 = ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n23225 = ~n23223;
  assign n26302 = ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n24287 = ~P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n24351 = ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n24665 = ~n24732;
  assign n38489 = ~n38562;
  assign n25644 = ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n27625 = ~n40471;
  assign n24039 = ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n24018 = ~P1_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n24432 = ~n24429;
  assign n42783 = ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n26806 = ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n23618 = ~n23630;
  assign n27094 = ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n28648 = ~P1_EAX_REG_27__SCAN_IN;
  assign n24435 = ~n24226 | ~n24225;
  assign n24565 = ~n24568;
  assign n24335 = ~n24334;
  assign n40672 = ~n42847;
  assign n23467 = ~n43408 & ~n35715;
  assign n43833 = ~n43832;
  assign n26479 = ~n40570;
  assign n39772 = ~n39775;
  assign n24422 = ~n24421;
  assign n28354 = ~P2_REIP_REG_29__SCAN_IN;
  assign n28302 = ~P2_REIP_REG_22__SCAN_IN;
  assign n42754 = ~n42753;
  assign n25626 = ~P2_EAX_REG_5__SCAN_IN;
  assign n42465 = ~n42716;
  assign n26283 = ~n26282;
  assign n27301 = ~n36311;
  assign n26179 = ~n35801;
  assign n40312 = ~n26460;
  assign n42206 = ~n42664;
  assign n26486 = ~n26485;
  assign n43660 = ~n43657;
  assign n42096 = ~n42307;
  assign n35439 = ~n35435;
  assign n26063 = ~n43712;
  assign n42546 = ~n42002 | ~n42001;
  assign n35366 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n42801 = ~BUF2_REG_27__SCAN_IN;
  assign n37271 = ~n36373 & ~n26913;
  assign n42657 = ~n42656;
  assign n41173 = ~n41172;
  assign n43605 = ~n43191 | ~n43190;
  assign n42255 = ~n42251 | ~n42250;
  assign n27867 = ~n27860 & ~n27859;
  assign n36562 = ~n37132;
  assign n38325 = ~n38336;
  assign n37374 = ~n37372;
  assign n35711 = ~n35708;
  assign n37577 = ~P3_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n40441 = ~n40371;
  assign n25065 = ~n37536 & ~n37535;
  assign n41191 = ~n27826 | ~n27825;
  assign n26570 = ~n40695;
  assign n34679 = ~n34576;
  assign n26910 = ~n26909;
  assign n43539 = ~P2_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n28123 = ~P2_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n36918 = ~P3_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n40748 = ~n41230;
  assign n37694 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n36661 = ~P3_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n30837 = ~n30861;
  assign n28928 = ~P3_STATE_REG_2__SCAN_IN;
  assign n26046 = ~n31276;
  assign n32136 = ~n32336;
  assign n28822 = ~n43720;
  assign n37846 = ~n37551;
  assign n31989 = ~P1_EAX_REG_16__SCAN_IN;
  assign n34243 = ~n39894;
  assign n43351 = ~P1_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n40089 = ~P1_REIP_REG_13__SCAN_IN;
  assign n39710 = ~n37469 & ~n37468;
  assign n41785 = ~n41568 | ~n41567;
  assign n38969 = ~n25487 | ~n25488;
  assign n43390 = ~n43058 & ~n43057;
  assign n32271 = ~n37303;
  assign n31252 = ~P2_EAX_REG_28__SCAN_IN;
  assign n28144 = ~P2_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n27852 = ~n27855 ^ n27853;
  assign n37286 = ~P2_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n43599 = ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n42303 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n39600 = ~n38332;
  assign n29471 = ~P2_REIP_REG_15__SCAN_IN;
  assign n39502 = ~P3_EBX_REG_22__SCAN_IN;
  assign n41391 = ~n41393;
  assign n34402 = ~n34404;
  assign n33527 = ~P3_EBX_REG_7__SCAN_IN;
  assign n31633 = ~P3_EAX_REG_16__SCAN_IN;
  assign n32499 = ~P3_EAX_REG_5__SCAN_IN;
  assign n34844 = ~BUF2_REG_12__SCAN_IN;
  assign n36220 = ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n40820 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n38732 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n36966 = ~P3_REIP_REG_4__SCAN_IN;
  assign n29381 = ~P3_REIP_REG_20__SCAN_IN;
  assign n44105 = ~n44098;
  assign n39741 = ~n39743;
  assign n35551 = ~n35553;
  assign n43931 = ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n36283 = ~n36237;
  assign n43967 = ~P3_EAX_REG_21__SCAN_IN;
  assign n22981 = n22980 | n22979;
  assign U214 = n39896 | n22988;
  assign n36557 = ~n23016 & ~n29171;
  assign n27891 = ~P2_STATE2_REG_0__SCAN_IN & ~n39522;
  assign n32176 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_STATE2_REG_2__SCAN_IN;
  assign n31487 = ~n32176;
  assign n35800 = ~P2_STATE2_REG_0__SCAN_IN | ~n31487;
  assign n23018 = ~n35800;
  assign n23541 = ~P2_FLUSH_REG_SCAN_IN | ~n23018;
  assign n23021 = ~n43499 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n23045 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n35718 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23036 = ~n23028 & ~n23027;
  assign n23464 = ~n43408 & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23035 = ~n23034 & ~n23033;
  assign n25645 = n43514 | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n26832 = ~n43094 & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n25652 = n26877 | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23051 = ~n23043 & ~n23042;
  assign n23044 = ~n43092 & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n25656 = ~n23044;
  assign n26726 = ~n25656;
  assign n23047 = ~n26726 | ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n26878 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23048 = ~n22905 & ~n41597;
  assign n23050 = ~n23049 & ~n23048;
  assign n23055 = ~n43499 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n23070 = ~n23062 & ~n23061;
  assign n23069 = ~n23068 & ~n23067;
  assign n23084 = ~n23070 | ~n23069;
  assign n23082 = ~n23076 & ~n23075;
  assign n26828 = ~n25656;
  assign n23079 = ~n22905 & ~n37629;
  assign n23081 = ~n23080 & ~n23079;
  assign n23088 = ~n26807 & ~n37739;
  assign n26789 = ~n35755 | ~n23105;
  assign n23086 = ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n23087 = ~n26789 & ~n23086;
  assign n23090 = ~n23088 & ~n23087;
  assign n25495 = ~n23467;
  assign n23095 = ~n22926 | ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n25440 = ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n23107 = ~n26791 & ~n25440;
  assign n26808 = ~n23105 | ~n23104;
  assign n23106 = ~n26808 & ~n41631;
  assign n23111 = ~n26838 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n25641 = ~n23468;
  assign n23114 = ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n23115 = ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n23129 = ~n26153 & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n26154 = P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ^ P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n39534 = ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n23138 = ~n26791 & ~n39534;
  assign n23137 = ~n26808 & ~n23136;
  assign n23140 = ~n23138 & ~n23137;
  assign n23139 = ~n22906 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n23142 = ~n26852 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n23141 = ~n26832 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n23146 = ~n26831 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n23145 = ~n26837 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n23148 = ~n26827 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n23147 = ~n26841 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n23153 = ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n23157 = ~n25652 & ~n23153;
  assign n23154 = ~n23481 | ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n23159 = ~n26828 | ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n23158 = ~n26838 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n23160 = n23159 & n23158;
  assign n23162 = ~n22926 | ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n34885 = ~n23167 | ~n23166;
  assign n23171 = ~n26154;
  assign n23267 = ~n23184 | ~n23183;
  assign n26317 = ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n23187 = ~n26789 & ~n26317;
  assign n23186 = ~n26807 & ~n37796;
  assign n23189 = ~n23187 & ~n23186;
  assign n23188 = ~n26848 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n23195 = ~n26837 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n23194 = ~n26832 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n23197 = ~n22926 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n23196 = ~n26841 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n23203 = ~n26791 & ~n26301;
  assign n23202 = ~n26808 & ~n26298;
  assign n23207 = ~n26828 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n23206 = ~n26838 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n23211 = ~n25645 & ~n26302;
  assign n23564 = ~n31498;
  assign n23281 = ~n23228 | ~n26505;
  assign n23231 = ~n26807 & ~n42782;
  assign n23229 = ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n23230 = ~n26789 & ~n23229;
  assign n26780 = ~n22926;
  assign n26737 = ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n23244 = ~n26791 & ~n26737;
  assign n23242 = ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n23243 = ~n26808 & ~n23242;
  assign n26341 = ~n23260 & ~n23259;
  assign n23270 = ~n32075 & ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n23282 = ~n23262 | ~n23261;
  assign n23274 = ~n23265 | ~n23264;
  assign n23276 = ~n23269 | ~n23268;
  assign n26168 = ~n23276 & ~n23275;
  assign n23280 = ~n23274 | ~n23273;
  assign n23285 = ~n32075 | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n23512 = ~n23277 | ~n23285;
  assign n23288 = ~n23280 | ~n23279;
  assign n23286 = ~n23284 | ~n23283;
  assign n26192 = ~n23286 | ~n23285;
  assign n23287 = ~n26192 | ~n23564;
  assign n31493 = ~n28196 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n25653 = ~n26838;
  assign n23291 = ~n25653 & ~n23289;
  assign n23295 = ~n23291 & ~n23290;
  assign n23292 = ~n26820 & ~n26779;
  assign n23294 = ~n23293 & ~n23292;
  assign n23297 = ~n25656 & ~n43099;
  assign n23299 = ~n23297 & ~n23296;
  assign n23302 = ~n43092 & ~n25285;
  assign n23308 = ~n25687 & ~n26345;
  assign n23307 = ~n26780 & ~n43082;
  assign n23309 = ~n23308 & ~n23307;
  assign n23319 = ~n23310 | ~n23309;
  assign n23311 = ~n25634 & ~n43097;
  assign n23315 = ~n25641 & ~n23313;
  assign n23314 = ~n25495 & ~n26346;
  assign n23320 = ~n23319 & ~n23318;
  assign n23322 = ~n23501;
  assign n23339 = n23328 | n23327;
  assign n23330 = ~n43499 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n23352 = ~n23339 & ~n23338;
  assign n23342 = ~n26858 | ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n23347 = ~n26828 | ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n23349 = ~n23347 | ~n23346;
  assign n23348 = ~n22905 & ~n42782;
  assign n23350 = ~n23349 & ~n23348;
  assign n36779 = ~n23352 | ~n22941;
  assign n23385 = ~n23322 & ~n36779;
  assign n23354 = ~n43499 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n23372 = ~n22906 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n23373 = ~n26858 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n23382 = ~n23376 & ~n23375;
  assign n23378 = ~n26726 | ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n23380 = ~n23378 | ~n23377;
  assign n23379 = ~n22905 & ~n35254;
  assign n23381 = ~n23380 & ~n23379;
  assign n23448 = ~n23385 | ~n23724;
  assign n23387 = ~n43499 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n23404 = ~n26726 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n23417 = ~n43499 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n23444 = ~n23438 & ~n23437;
  assign n23440 = ~n26726 | ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n23441 = ~n22905 & ~n37739;
  assign n23443 = ~n23442 & ~n23441;
  assign n36688 = n23490;
  assign n26184 = ~n36779;
  assign n23585 = ~n36688 | ~n26184;
  assign n23450 = ~n23493 | ~n23585;
  assign n23451 = ~n23450 | ~n23449;
  assign n23544 = ~n23452 | ~n23451;
  assign n23454 = ~n43499 | ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n23489 = ~n23474 | ~n23473;
  assign n23483 = ~n26726 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n23484 = ~n22905 & ~n37796;
  assign n23488 = ~n23487 | ~n23486;
  assign n23520 = ~n23415 | ~n23575;
  assign n23495 = ~n23493;
  assign n23494 = ~n25093 & ~n36779;
  assign n23496 = ~n23495 | ~n23494;
  assign n26200 = ~n23496 & ~n23520;
  assign n23498 = ~n23523 | ~n23497;
  assign n23502 = ~n23415 | ~n23501;
  assign n23505 = n23502 & n37289;
  assign n23711 = ~n23505 & ~n23504;
  assign n23730 = ~n37289 | ~n36795;
  assign n23706 = ~n23730 & ~n36688;
  assign n31058 = ~n23711 | ~n23706;
  assign n23506 = ~n23571 & ~n26507;
  assign n23508 = ~n26167;
  assign n31770 = ~n23513 | ~n26177;
  assign n25099 = ~n23516 | ~n23515;
  assign n32148 = ~n31779 & ~n31777;
  assign n31057 = ~n26546 & ~n31770;
  assign n29085 = ~P2_STATE_REG_1__SCAN_IN & ~P2_STATE_REG_2__SCAN_IN;
  assign n23518 = ~n29085 & ~P2_STATE_REG_0__SCAN_IN;
  assign n23517 = ~P2_STATE_REG_1__SCAN_IN | ~P2_STATE_REG_2__SCAN_IN;
  assign n31819 = ~n23518 | ~n23517;
  assign n23532 = n26180 | n31819;
  assign n23519 = ~n26184 & ~n23127;
  assign n23521 = ~n23519 & ~n23728;
  assign n23522 = ~n23521 & ~n23520;
  assign n23527 = ~n23522 & ~n25093;
  assign n23562 = ~n23523;
  assign n23554 = ~n23524 & ~n23562;
  assign n23525 = ~n32217 | ~n28196;
  assign n23526 = ~n23554 | ~n23525;
  assign n23530 = n23527 | n23526;
  assign n23553 = ~n25491 & ~n26184;
  assign n23528 = ~n23553 & ~n25093;
  assign n23529 = ~n23733 & ~n23528;
  assign n23533 = ~n32148 & ~n26189;
  assign n31766 = ~n23733 | ~n23127;
  assign n28197 = ~n35802 & ~n31819;
  assign n23535 = ~n28197;
  assign n23536 = ~n31766 & ~n23535;
  assign n23701 = ~n23546 & ~n23545;
  assign n23550 = ~n23547 & ~n33357;
  assign n23555 = ~n23553 & ~n22904;
  assign n23715 = ~n23556 | ~n23575;
  assign n23557 = ~n23415 & ~n36779;
  assign n25096 = ~n23557 | ~n23562;
  assign n23702 = ~n25096 | ~n36795;
  assign n23593 = ~n23715 | ~n23702;
  assign n23561 = ~n23560 | ~n23559;
  assign n23574 = ~n23630 & ~n23684;
  assign n25532 = ~n22900 & ~n22904;
  assign n23563 = n25532 & n36561;
  assign n23731 = ~n23563 | ~n23562;
  assign n23569 = ~n23567 & ~n23566;
  assign n35707 = ~n23729 | ~n23568;
  assign n23572 = ~n23583 & ~n23570;
  assign n23573 = ~n23572 | ~n23635;
  assign n23582 = ~n28346 & ~n29550;
  assign n23598 = ~n23578 & ~n25096;
  assign n23580 = ~n23598 | ~P2_EBX_REG_1__SCAN_IN;
  assign n23590 = ~n23582 & ~n23581;
  assign n41873 = ~n23322;
  assign n23584 = ~n25093 & ~n41873;
  assign n23659 = ~n23724 & ~n36357;
  assign n23610 = ~n23723 | ~n23659;
  assign n27912 = ~n23588 | ~n23610;
  assign n23589 = ~n27912 | ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n23614 = ~n23590 | ~n23589;
  assign n23597 = ~n23635 & ~n23592;
  assign n39573 = n23598;
  assign n23601 = ~n39573 | ~P2_EBX_REG_0__SCAN_IN;
  assign n23599 = P2_STATE2_REG_1__SCAN_IN & P2_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n23602 = ~n23601 | ~n23600;
  assign n23604 = ~n23603 & ~n23602;
  assign n26527 = ~n27912;
  assign n23606 = ~n26527 & ~n33579;
  assign n23675 = ~n23607 & ~n23606;
  assign n23612 = ~n23630 & ~n26153;
  assign n23609 = ~n39573 & ~n23608;
  assign n23676 = ~n23675 & ~n23674;
  assign n23616 = ~n23615 & ~n23614;
  assign n23623 = ~n23634;
  assign n23633 = ~n23621 | ~n23620;
  assign n23666 = ~n23623 | ~n23622;
  assign n26512 = ~n23666;
  assign n23625 = ~n27912 | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n23624 = ~n23591 | ~P2_REIP_REG_3__SCAN_IN;
  assign n23627 = ~n39573 | ~P2_EBX_REG_3__SCAN_IN;
  assign n26518 = ~n23632 & ~n23631;
  assign n23646 = ~n26512 | ~n23644;
  assign n23643 = ~n23665;
  assign n28361 = n23635;
  assign n23640 = ~n23635 & ~n23636;
  assign n23638 = ~n39573 | ~P2_EBX_REG_2__SCAN_IN;
  assign n23641 = ~n27912 | ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n26513 = ~n23643 & ~n23667;
  assign n23650 = ~n23646 | ~n23645;
  assign n23648 = ~n23666 | ~n23647;
  assign n23651 = ~n23650 & ~n23649;
  assign n36607 = ~n23651;
  assign n38820 = ~n36607;
  assign n31816 = ~n39511 & ~P2_STATE2_REG_0__SCAN_IN;
  assign n23658 = ~n38820 & ~n27927;
  assign n23685 = ~n23652 & ~P2_STATE2_REG_3__SCAN_IN;
  assign n23653 = ~n37634 & ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n39508 = ~P2_STATE2_REG_3__SCAN_IN & ~P2_STATE2_REG_2__SCAN_IN;
  assign n42796 = ~n23660 & ~n43061;
  assign n25105 = ~n23661 | ~n23662;
  assign n25107 = ~n23664 | ~n23663;
  assign n23699 = ~n25105 | ~n25107;
  assign n23668 = ~n23666 | ~n23665;
  assign n23669 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n23672 = ~n23671 & ~n23670;
  assign n23677 = ~n23675 | ~n23674;
  assign n23683 = ~n23676;
  assign n23682 = ~n37279 & ~n27927;
  assign n23690 = ~n23682 & ~n23681;
  assign n32143 = n23690 ^ n23691;
  assign n37852 = n37635 ^ P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n32892 = ~n23694 | ~n23693;
  assign n32896 = ~n32891 | ~n32892;
  assign n25106 = ~n32896 | ~n23698;
  assign n36533 = ~n31779 | ~P2_STATE2_REG_3__SCAN_IN;
  assign n23744 = ~n37131 & ~n36533;
  assign n23710 = ~n23701;
  assign n23704 = ~n23702;
  assign n23705 = ~n23704 | ~n23703;
  assign n23707 = ~n23706;
  assign n23713 = ~n23711;
  assign n23712 = ~n28196;
  assign n31522 = ~n23127 | ~n37289;
  assign n26506 = ~n26200;
  assign n35750 = ~n26209;
  assign n23742 = ~n38820 & ~n35750;
  assign n23718 = ~n44000;
  assign n35725 = ~n23719 | ~n23718;
  assign n35721 = ~n23720 & ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23721 = ~n35721 ^ n35715;
  assign n23740 = n35725 | n23721;
  assign n26509 = ~n23723;
  assign n23725 = ~n26509 & ~n23724;
  assign n35722 = ~n32147 & ~n23725;
  assign n43484 = ~n43514;
  assign n23726 = ~n43484 & ~n35715;
  assign n23727 = ~n22906 & ~n23726;
  assign n23738 = ~n35722 & ~n23727;
  assign n26508 = ~n23729 | ~n23728;
  assign n23732 = ~n23731 & ~n23730;
  assign n23734 = ~n23733 & ~n23732;
  assign n35752 = ~n26508 | ~n23734;
  assign n23736 = ~n35752;
  assign n35729 = ~n32506;
  assign n23735 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ n35729;
  assign n23737 = ~n23736 & ~n23735;
  assign n23739 = ~n23738 & ~n23737;
  assign n23741 = ~n23740 | ~n23739;
  assign n35714 = ~n23742 & ~n23741;
  assign n23743 = ~n36532 & ~n35714;
  assign n23745 = ~n23744 & ~n23743;
  assign n23747 = ~n36543 & ~n23745;
  assign n23746 = ~n36542 & ~n35715;
  assign P2_U3596 = n23747 | n23746;
  assign n35113 = ~P1_INSTADDRPOINTER_REG_6__SCAN_IN | ~P1_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n23748 = ~n35113;
  assign n35112 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN | ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n34283 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN | ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n35099 = ~n35112 & ~n34283;
  assign n25950 = ~n23748 | ~n35099;
  assign n33721 = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23772 = ~n33721 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n24795 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n24515 = ~n32127 | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n31922 = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n24517 = ~n32127 | ~n31922;
  assign n32084 = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n32118 = ~n32084;
  assign n32121 = ~n32118 | ~n22928;
  assign n23769 = ~n33721 & ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n24539 = ~n23769 | ~n33727;
  assign n26095 = ~n31938 | ~n23769;
  assign n24526 = ~n23769 | ~n32118;
  assign n24527 = ~n32118 | ~n32119;
  assign n23788 = ~n23768 & ~n23767;
  assign n27006 = ~n31938 | ~n32119;
  assign n23771 = ~n43260 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n31937 = ~n24795 & ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n28585 = ~n23769 | ~n31937;
  assign n23770 = ~n43274 | ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n27004 = ~n31938 | ~n23777;
  assign n23774 = ~n43245 | ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n28591 = ~n31937 | ~n22928;
  assign n23773 = ~n43275 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n27011 = ~n23777 | ~n33727;
  assign n23779 = ~n43265 | ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n26659 = ~n31937 | ~n32119;
  assign n23778 = ~n43264 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n28593 = ~n22928 | ~n33727;
  assign n27009 = ~n31938 | ~n22928;
  assign n23780 = ~n22908 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n23786 = ~n23785 | ~n23784;
  assign n39891 = ~n23788 | ~n23787;
  assign n23790 = ~n24515 & ~n24341;
  assign n23789 = ~n24517 & ~n24373;
  assign n23794 = ~n23790 & ~n23789;
  assign n23793 = ~n23792 & ~n23791;
  assign n23802 = ~n23794 | ~n23793;
  assign n23795 = ~n32121 & ~n24367;
  assign n23800 = ~n23796 & ~n23795;
  assign n23798 = ~n26095 & ~n24356;
  assign n23797 = ~n27006 & ~n24374;
  assign n23799 = ~n23798 & ~n23797;
  assign n23801 = ~n23800 | ~n23799;
  assign n23818 = ~n23802 & ~n23801;
  assign n23804 = ~n27009 & ~n24378;
  assign n23803 = ~n27011 & ~n24346;
  assign n23808 = ~n23804 & ~n23803;
  assign n23806 = ~n28591 & ~n24351;
  assign n23807 = ~n23806 & ~n23805;
  assign n23816 = ~n23808 | ~n23807;
  assign n23812 = ~n28593 & ~n24345;
  assign n23813 = ~n23812 & ~n23811;
  assign n23817 = ~n23816 & ~n23815;
  assign n31382 = ~n22947;
  assign n23847 = ~n23832 & ~n23831;
  assign n23834 = ~n43260 | ~P1_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n43270 = ~n26095;
  assign n23833 = ~n43270 | ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n23836 = ~n43274 | ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n23835 = ~n43261 | ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n23840 = ~n43245 | ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n23839 = ~n43242 | ~P1_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n23842 = ~n43251 | ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n23841 = ~n43246 | ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n23845 = ~n23844 & ~n23843;
  assign n23875 = ~n43265 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n23874 = ~n43264 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n43271 = ~n28587;
  assign n23876 = ~n43270 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n23887 = ~n23879 & ~n23878;
  assign n23881 = ~n43260 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n23883 = ~n43261 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n23882 = ~n22908 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n23886 = ~n23885 & ~n23884;
  assign n24122 = ~n31382 | ~n24392;
  assign n23895 = n23889 | n24706;
  assign n24394 = ~n24122;
  assign n24872 = ~n24394 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n23945 = ~n24872 & ~n24745;
  assign n24655 = ~n24872;
  assign n23923 = n23945 | n23903;
  assign n23906 = n31922 ^ P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n24200 = ~n34097 & ~n24392;
  assign n23907 = ~n23906;
  assign n35466 = ~n22947 | ~n34187;
  assign n23941 = ~n23932 | ~n23931;
  assign n23940 = n23935 | n23934;
  assign n23939 = ~n23938 & ~n23937;
  assign n23947 = ~n23940 | ~n23939;
  assign n24101 = ~n23944 | ~n23943;
  assign n23949 = ~n23947 | ~n23946;
  assign n23948 = ~n24101 | ~n24654;
  assign n23950 = ~n22907 | ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n23952 = ~n43265 | ~P1_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n23967 = ~n43245 | ~P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n23966 = ~n43242 | ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n23973 = ~n43274 | ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n23978 = ~n23977 | ~n23976;
  assign n24002 = ~n43260 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n24001 = ~n43270 | ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n24004 = ~n43274 | ~P1_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n24003 = ~n43261 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n24014 = ~n24006 & ~n24005;
  assign n24008 = ~n43245 | ~P1_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n24007 = ~n43242 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n24012 = ~n24008 | ~n24007;
  assign n24010 = ~n43251 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n24009 = ~n43246 | ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n24011 = ~n24010 | ~n24009;
  assign n24013 = ~n24012 & ~n24011;
  assign n24061 = ~n24037 & ~n24036;
  assign n24060 = ~n24059 & ~n24058;
  assign n24092 = ~n24406 | ~n32238;
  assign n25069 = ~n24392 & ~n39891;
  assign n24062 = ~n22907 | ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n24091 = ~n24075 | ~n24074;
  assign n24090 = ~n24089 | ~n24088;
  assign n24093 = ~n31721 & ~n34515;
  assign n31478 = ~READY11_REG_SCAN_IN | ~READY1;
  assign n39895 = ~n39892 & ~n34149;
  assign n24094 = ~n39895 & ~n22947;
  assign n24107 = ~n24096 | ~n34226;
  assign n31374 = ~n34515;
  assign n24104 = ~n31721 | ~n31374;
  assign n24106 = ~n24105 | ~n31891;
  assign n32239 = ~n34149 | ~n39891;
  assign n24149 = ~n24392 | ~n32238;
  assign n24110 = ~n24200 | ~n31891;
  assign n24113 = ~n24112 & ~n39892;
  assign n24120 = ~n24199 | ~n24208;
  assign n24134 = ~n24118 | ~n32238;
  assign n24123 = ~n32239;
  assign n24124 = ~n24123 & ~n24122;
  assign n31715 = ~n34187 | ~n31382;
  assign n24509 = ~n33714 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n44102 = ~n24509 & ~n33710;
  assign n35474 = ~n34187 & ~n31382;
  assign n31892 = ~n35474;
  assign n24131 = ~n24130 & ~n31892;
  assign n32080 = ~n24216 | ~n24131;
  assign n42922 = ~n24132 | ~n32131;
  assign n24148 = ~n24246;
  assign n31477 = ~n31715;
  assign n24136 = ~n24134 | ~n31477;
  assign n24240 = ~n24136 | ~n24135;
  assign n40073 = ~n34187 & ~n34164;
  assign n28825 = ~n40073;
  assign n24235 = ~n34164 | ~n31382;
  assign n24138 = ~n24165 | ~n24137;
  assign n24206 = ~n24139 | ~n24138;
  assign n24146 = ~n24206;
  assign n24144 = ~n24222 & ~n28825;
  assign n24140 = ~n26568 | ~n34134;
  assign n24141 = ~n24140 | ~n35474;
  assign n24143 = ~n24142 | ~n24141;
  assign n24145 = ~n24144 & ~n24143;
  assign n24147 = ~n24146 | ~n24145;
  assign n24151 = ~n24802 & ~n24149;
  assign n25068 = ~n24150 & ~n31891;
  assign n32123 = ~n24151 | ~n25068;
  assign n24152 = n31920 & n32123;
  assign n42924 = ~n24205 & ~n24152;
  assign n24154 = ~n25950 & ~n34279;
  assign n36891 = ~n31447 & ~n24205;
  assign n24420 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n32540 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN | ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n34290 = n24420 & n32540;
  assign n35100 = n35112 | n34290;
  assign n25952 = ~n35100 & ~n35113;
  assign n24153 = n36891 & n25952;
  assign n24155 = ~P1_INSTADDRPOINTER_REG_8__SCAN_IN & ~P1_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n24752 = ~P1_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n24738 = ~P1_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n25951 = ~n24752 & ~n24738;
  assign n24156 = n24155 | n25951;
  assign n24762 = ~n36890 & ~n24156;
  assign n24158 = ~n25952 & ~n41976;
  assign n39315 = ~P1_STATE2_REG_2__SCAN_IN & ~P1_STATE2_REG_3__SCAN_IN;
  assign n32552 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n24160 = ~n24158 & ~n38650;
  assign n24159 = ~n41979 | ~n25950;
  assign n35833 = ~n24160 | ~n24159;
  assign n24760 = ~n35833 | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n32232 = ~n24161 & ~n35466;
  assign n24163 = ~n24425 & ~n24392;
  assign n31358 = ~n31916 & ~n31715;
  assign n24164 = ~n24163 & ~n31358;
  assign n43344 = ~n24205 & ~n24164;
  assign n31705 = ~P1_EBX_REG_0__SCAN_IN;
  assign n37246 = ~n35821 ^ n25076;
  assign n24758 = ~n43441 & ~n37246;
  assign n24198 = ~n24425 & ~n34134;
  assign n24197 = ~n31916 & ~n40081;
  assign n24202 = ~n24198 & ~n24197;
  assign n24201 = ~n39895 | ~n24200;
  assign n31449 = ~n31907 & ~n34498;
  assign n36906 = ~n24205 & ~n24204;
  assign n24213 = ~n24206 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n31898 = ~n31451 | ~n32238;
  assign n24424 = ~n31898 & ~n24211;
  assign n24212 = ~n24424 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n24217 = ~n24216 | ~n34187;
  assign n24727 = ~n31382 & ~n33710;
  assign n24218 = ~n39895 | ~n40073;
  assign n24241 = ~n32123 | ~n24218;
  assign n24231 = ~n24222 | ~n24221;
  assign n24224 = ~n22932 | ~n24223;
  assign n24225 = ~n22930 & ~n24224;
  assign n24230 = ~n24435 | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n24338 = ~n24247 | ~n24246;
  assign n31936 = ~n24340 | ~n24338;
  assign n24429 = ~n24252 | ~n24251;
  assign n24253 = n31936 ^ n24429;
  assign n24298 = ~n24253 & ~P1_STATE2_REG_0__SCAN_IN;
  assign n24477 = ~n34134 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n24254 = ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n24257 = ~n24515 & ~n24254;
  assign n24256 = ~n24517 & ~n24255;
  assign n24258 = ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n24260 = ~n28591 & ~n24258;
  assign n24259 = ~n32121 & ~n26099;
  assign n24263 = ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n24266 = ~n27011 & ~n24263;
  assign n24265 = ~n27006 & ~n24264;
  assign n24269 = ~n27009 & ~n24267;
  assign n24268 = ~n24527 & ~n26096;
  assign n24274 = ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n24277 = ~n28585 & ~n24274;
  assign n24276 = ~n27004 & ~n24275;
  assign n24279 = ~n24526 & ~n26094;
  assign n24278 = ~n26659 & ~n26100;
  assign n24282 = ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n24285 = ~n26095 & ~n24282;
  assign n24284 = ~n28587 & ~n24283;
  assign n24286 = ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n24289 = ~n24539 & ~n24286;
  assign n24288 = ~n28593 & ~n24287;
  assign n24749 = ~n24328 & ~n24327;
  assign n24399 = ~n24485 & ~n24337;
  assign n24390 = ~n34552 | ~n33710;
  assign n24344 = ~n24517 & ~n24341;
  assign n24343 = ~n24515 & ~n24342;
  assign n24350 = ~n24344 & ~n24343;
  assign n24348 = ~n24526 & ~n24345;
  assign n24347 = ~n24527 & ~n24346;
  assign n24349 = ~n24348 & ~n24347;
  assign n24354 = ~n27009 & ~n24351;
  assign n24353 = ~n26659 & ~n24352;
  assign n24360 = ~n24354 & ~n24353;
  assign n24358 = ~n32121 & ~n24355;
  assign n24357 = ~n24539 & ~n24356;
  assign n24359 = ~n24358 & ~n24357;
  assign n24366 = ~n28585 & ~n24363;
  assign n24365 = ~n26095 & ~n24364;
  assign n24372 = ~n24366 & ~n24365;
  assign n24370 = ~n28591 & ~n24367;
  assign n24369 = ~n27006 & ~n24368;
  assign n24371 = ~n24370 & ~n24369;
  assign n24376 = ~n27004 & ~n24373;
  assign n24375 = ~n28587 & ~n24374;
  assign n24382 = ~n24376 & ~n24375;
  assign n24380 = ~n27011 & ~n24377;
  assign n24379 = ~n28593 & ~n24378;
  assign n24381 = ~n24380 & ~n24379;
  assign n24412 = ~n24390 | ~n24389;
  assign n24397 = ~n24749 & ~n24392;
  assign n24398 = ~n24412 | ~n24411;
  assign n25895 = ~n24397 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n24400 = ~n24398 | ~n25895;
  assign n24403 = ~n24399 & ~n24400;
  assign n24402 = ~n24399;
  assign n24484 = ~n24402 & ~n24401;
  assign n34560 = ~n24403 & ~n24484;
  assign n24410 = ~n34560 | ~n26568;
  assign n24404 = ~n24489 ^ n24488;
  assign n24408 = ~n24404 & ~n31715;
  assign n24407 = ~n24406 | ~n24405;
  assign n24409 = ~n24408 & ~n24407;
  assign n24416 = ~n24410 | ~n24409;
  assign n34551 = n24412 ^ n24411;
  assign n24415 = ~n34551 | ~n26568;
  assign n24413 = ~n31715 & ~n24488;
  assign n24491 = ~n34164 & ~n31382;
  assign n24414 = ~n24413 & ~n24491;
  assign n31687 = ~n24415 | ~n24414;
  assign n24417 = ~n31687 | ~P1_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n32062 = n24416 ^ n24417;
  assign n32556 = ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n32061 = ~n32062 & ~n32556;
  assign n24421 = ~n32061 & ~n24419;
  assign n24495 = ~n24421 & ~n24420;
  assign n24423 = ~n24422 & ~P1_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n32546 = ~n24495 & ~n24423;
  assign n24428 = ~n32337 & ~n24427;
  assign n35165 = ~n24429 ^ n24430;
  assign n24446 = ~n24442 | ~n24443;
  assign n36136 = ~n24446 | ~n32334;
  assign n24563 = ~n24476 & ~n24475;
  assign n24478 = ~n24477 & ~n24563;
  assign n24499 = n24500 ^ n24483;
  assign n24487 = ~n24484;
  assign n24497 = ~n24487 | ~n24486;
  assign n24564 = ~n24489 | ~n24488;
  assign n24490 = n24564 ^ n24563;
  assign n24492 = ~n24490 & ~n31715;
  assign n24493 = ~n24492 & ~n24491;
  assign n32547 = ~n32546 | ~n32545;
  assign n34057 = ~n32547 | ~n24496;
  assign n24498 = ~n24497;
  assign n24502 = ~n24499 | ~n24498;
  assign n24513 = ~n24503 & ~n33721;
  assign n24514 = ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n24519 = ~n24515 & ~n24514;
  assign n24516 = ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n24518 = ~n24517 & ~n24516;
  assign n24520 = ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n24522 = ~n27004 & ~n24520;
  assign n24521 = ~n32121 & ~n28592;
  assign n24525 = ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n24529 = ~n24526 & ~n24525;
  assign n24528 = ~n24527 & ~n28586;
  assign n26662 = ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n24532 = ~n26659 & ~n26662;
  assign n24530 = ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n24531 = ~n28587 & ~n24530;
  assign n24541 = ~n28591 & ~n24537;
  assign n24538 = ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n24540 = ~n24539 & ~n24538;
  assign n24542 = ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n24544 = ~n26095 & ~n24542;
  assign n28590 = ~P1_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n24543 = ~n27006 & ~n28590;
  assign n24547 = ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n24549 = ~n28585 & ~n24547;
  assign n28584 = ~P1_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n24548 = ~n27009 & ~n28584;
  assign n26658 = ~P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n24552 = ~n27011 & ~n26658;
  assign n24550 = ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n24551 = ~n28593 & ~n24550;
  assign n24561 = ~n24560 & ~n24559;
  assign n24573 = ~n22916 & ~n24745;
  assign n24569 = ~n24564 | ~n24563;
  assign n24566 = ~n24569;
  assign n24567 = ~n24566 | ~n24565;
  assign n24571 = ~n24567 | ~n31477;
  assign n24570 = ~n24659;
  assign n24572 = ~n24571 & ~n24570;
  assign n35322 = ~n24573 & ~n24572;
  assign n34055 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n24574 = ~n35322 | ~n34055;
  assign n24622 = ~n34057 | ~n24574;
  assign n24616 = ~n24659 ^ n24658;
  assign n24617 = ~n24616 & ~n31715;
  assign n35332 = ~n24618 & ~n24617;
  assign n24619 = ~n35322 & ~n34055;
  assign n24621 = ~n24620 & ~n24619;
  assign n24674 = ~n24622 | ~n24621;
  assign n24664 = n24653 | n24652;
  assign n24712 = ~n24657 | ~n24656;
  assign n24668 = ~n24841 & ~n24745;
  assign n24661 = ~n24664;
  assign n24663 = ~n24659 & ~n24658;
  assign n24660 = ~n24663;
  assign n24662 = ~n24661 | ~n24660;
  assign n24666 = ~n24662 | ~n31477;
  assign n24667 = ~n24666 & ~n24665;
  assign n24669 = ~n24668 & ~n24667;
  assign n36128 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n24671 = ~n24669 | ~n36128;
  assign n24675 = ~n24670 | ~P1_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n36086 = ~n24671 | ~n24675;
  assign n24673 = ~n36086 & ~n24672;
  assign n36091 = ~n24674 | ~n24673;
  assign n35109 = ~n36091 | ~n24675;
  assign n24691 = ~n43275 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n24690 = ~n43264 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n24693 = ~n43274 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n24692 = ~n43265 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n24697 = ~n22908 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n24696 = ~n43261 | ~P1_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n24699 = ~n43260 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n24698 = ~n43271 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n24714 = n24713 & n24712;
  assign n24719 = ~n24718 | ~n31477;
  assign n35104 = ~P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n24724 = ~n24721 & ~n35104;
  assign n35108 = ~n24724 & ~n24723;
  assign n35110 = ~n35109 | ~n35108;
  assign n35831 = ~n35110 | ~n24725;
  assign n24747 = ~n24733 & ~n24732;
  assign n24736 = ~n24735 & ~n31715;
  assign n24744 = ~n35831 | ~n35832;
  assign n25962 = ~n24744 | ~n24743;
  assign n24748 = ~n24747;
  assign n24750 = ~n24749 & ~n24748;
  assign n24755 = ~n25965 | ~n25963;
  assign n43469 = ~n43033;
  assign n37006 = ~n43469 | ~P1_REIP_REG_8__SCAN_IN;
  assign P1_U3023 = n24762 | n24761;
  assign n24764 = ~P2_STATE2_REG_0__SCAN_IN & ~n37286;
  assign n24763 = ~n36357 & ~n33579;
  assign n37285 = ~n24764 & ~n24763;
  assign n24767 = ~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n28146 = ~P2_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n28122 = ~P2_PHYADDRPOINTER_REG_2__SCAN_IN | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n28118 = ~n28123 & ~n28122;
  assign n24769 = ~n37285 | ~n41718;
  assign n24768 = ~n41204 | ~n33579;
  assign n24774 = ~P2_STATE2_REG_1__SCAN_IN | ~n36500;
  assign n36365 = ~n36532;
  assign n24770 = ~n34876 | ~n26209;
  assign n35756 = ~n35722 | ~n35725;
  assign n35751 = ~n35756 | ~n26153;
  assign n24772 = n24770 & n35751;
  assign n24771 = ~n35752 | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n35749 = ~n24772 | ~n24771;
  assign n24773 = ~n36365 | ~n35749;
  assign n24783 = ~n24774 | ~n24773;
  assign n24776 = ~n36357 & ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n24782 = ~n38279 & ~n36533;
  assign n24784 = ~n24783 & ~n24782;
  assign n24786 = ~n36543 & ~n24784;
  assign n24785 = ~n36542 & ~n26153;
  assign P2_U3601 = n24786 | n24785;
  assign n24873 = ~n34149 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n43722 = ~P1_STATE2_REG_2__SCAN_IN;
  assign n24815 = ~n24787 | ~n24864;
  assign n24792 = ~n28810 & ~n24788;
  assign n24790 = ~n28608 | ~P1_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n43294 = ~P1_STATE2_REG_2__SCAN_IN & ~P1_STATEBS16_REG_SCAN_IN;
  assign n36144 = ~P1_PHYADDRPOINTER_REG_1__SCAN_IN ^ P1_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n24789 = ~n43294 | ~n36144;
  assign n32630 = n24815 ^ n24814;
  assign n24799 = ~n24831 & ~n24795;
  assign n24796 = ~n43722 | ~P1_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n24806 = ~n24831 & ~n31922;
  assign n24805 = ~n28810 & ~n24804;
  assign n24809 = ~P1_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n24810 = ~n24809 & ~P1_STATE2_REG_2__SCAN_IN;
  assign n32631 = ~n32630 | ~n32629;
  assign n33313 = ~n32631 | ~n24816;
  assign n24827 = ~n34270 | ~n25932;
  assign n35889 = P1_PHYADDRPOINTER_REG_3__SCAN_IN ^ n24829;
  assign n43725 = ~n43294;
  assign n24821 = ~n28810 & ~n24818;
  assign n24819 = ~P1_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n24820 = ~n24864 & ~n24819;
  assign n33314 = ~n24827 | ~n24826;
  assign n33794 = ~n33313 | ~n33314;
  assign n24832 = P1_PHYADDRPOINTER_REG_4__SCAN_IN & n43722;
  assign n24850 = n24841 | n24873;
  assign n24844 = ~P1_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n35820 = ~n34812 ^ n24860;
  assign n36992 = P1_PHYADDRPOINTER_REG_7__SCAN_IN ^ n24906;
  assign n24868 = n36992 | n43725;
  assign n24863 = ~P1_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n24865 = ~n24864 & ~n24863;
  assign n24870 = ~n35820 & ~n35819;
  assign n36273 = ~n24870 & ~n24869;
  assign n24876 = ~n43274 | ~P1_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n24875 = ~n22915 | ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n24880 = ~n24876 | ~n24875;
  assign n24878 = ~n43270 | ~P1_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n24877 = ~n22908 | ~P1_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n24879 = ~n24878 | ~n24877;
  assign n24888 = ~n24880 & ~n24879;
  assign n24882 = ~n43260 | ~P1_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n24881 = ~n43261 | ~P1_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n24886 = ~n24882 | ~n24881;
  assign n24884 = ~n43245 | ~P1_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n24883 = ~n43275 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n24885 = ~n24884 | ~n24883;
  assign n24887 = ~n24886 & ~n24885;
  assign n24890 = ~n43246 | ~P1_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n24889 = ~n43251 | ~P1_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n24894 = ~n24890 | ~n24889;
  assign n24892 = ~n43264 | ~P1_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n24891 = ~n43242 | ~P1_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n24893 = ~n24892 | ~n24891;
  assign n24902 = ~n24894 & ~n24893;
  assign n24896 = ~n22907 | ~P1_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n24895 = ~n43241 | ~P1_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n24900 = ~n24896 | ~n24895;
  assign n24898 = ~n43265 | ~P1_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n24897 = ~n43271 | ~P1_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n24899 = ~n24898 | ~n24897;
  assign n24901 = ~n24900 & ~n24899;
  assign n24912 = n22942 | n24905;
  assign n24914 = ~n43270 | ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n24913 = ~n43271 | ~P1_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n24918 = ~n24914 | ~n24913;
  assign n24916 = ~n43245 | ~P1_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n24915 = ~n43275 | ~P1_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n24917 = ~n24916 | ~n24915;
  assign n24926 = ~n24918 & ~n24917;
  assign n24920 = ~n43260 | ~P1_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n24919 = ~n43261 | ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n24924 = ~n24920 | ~n24919;
  assign n24922 = ~n43264 | ~P1_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n24921 = ~n43265 | ~P1_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n24923 = ~n24922 | ~n24921;
  assign n24925 = ~n24924 & ~n24923;
  assign n24942 = ~n24926 | ~n24925;
  assign n24928 = ~n22907 | ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n24927 = ~n43251 | ~P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n24932 = ~n24928 | ~n24927;
  assign n24930 = ~n28775 | ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n24929 = ~n22915 | ~P1_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n24931 = ~n24930 | ~n24929;
  assign n24940 = ~n24932 & ~n24931;
  assign n24934 = ~n43246 | ~P1_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n24933 = ~n43242 | ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n24938 = ~n24934 | ~n24933;
  assign n24936 = ~n43274 | ~P1_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n24935 = ~n22908 | ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n24937 = ~n24936 | ~n24935;
  assign n24939 = ~n24938 & ~n24937;
  assign n24951 = ~n43275 | ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n24950 = ~n43265 | ~P1_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n24955 = ~n24951 | ~n24950;
  assign n24953 = ~n43245 | ~P1_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n24952 = ~n43271 | ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n24954 = ~n24953 | ~n24952;
  assign n24963 = ~n24955 & ~n24954;
  assign n24957 = ~n43270 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n24956 = ~n43264 | ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n24961 = ~n24957 | ~n24956;
  assign n24959 = ~n22908 | ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n24958 = ~n43260 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n24960 = ~n24959 | ~n24958;
  assign n24962 = ~n24961 & ~n24960;
  assign n24979 = ~n24963 | ~n24962;
  assign n24965 = ~n22907 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n24964 = ~n43246 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n24969 = ~n24965 | ~n24964;
  assign n24967 = ~n28775 | ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n24966 = ~n43274 | ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n24968 = ~n24967 | ~n24966;
  assign n24977 = ~n24969 & ~n24968;
  assign n24971 = ~n43251 | ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n24970 = ~n43242 | ~P1_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n24975 = ~n24971 | ~n24970;
  assign n24973 = ~n43261 | ~P1_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n24972 = ~n22915 | ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n24974 = ~n24973 | ~n24972;
  assign n24976 = ~n24975 & ~n24974;
  assign n24987 = n22942 | n24980;
  assign n24989 = ~n43275 | ~P1_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n24988 = ~n43261 | ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n24993 = ~n24989 | ~n24988;
  assign n24991 = ~n22915 | ~P1_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n24990 = ~n43271 | ~P1_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n24992 = ~n24991 | ~n24990;
  assign n25001 = ~n24993 & ~n24992;
  assign n24995 = ~n28775 | ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n24994 = ~n43274 | ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n24999 = ~n24995 | ~n24994;
  assign n24997 = ~n43270 | ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n24996 = ~n43265 | ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n24998 = ~n24997 | ~n24996;
  assign n25000 = ~n24999 & ~n24998;
  assign n25017 = ~n25001 | ~n25000;
  assign n25003 = ~n43246 | ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n25002 = ~n43242 | ~P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n25007 = ~n25003 | ~n25002;
  assign n25005 = ~n43245 | ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n25004 = ~n22908 | ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n25006 = ~n25005 | ~n25004;
  assign n25015 = ~n25007 & ~n25006;
  assign n25009 = ~n22907 | ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n25008 = ~n43251 | ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n25013 = ~n25009 | ~n25008;
  assign n25011 = ~n43260 | ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n25010 = ~n43264 | ~P1_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n25012 = ~n25011 | ~n25010;
  assign n25014 = ~n25013 & ~n25012;
  assign n25016 = ~n25015 | ~n25014;
  assign n25018 = ~n25017 & ~n25016;
  assign n25028 = ~n22907 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n25027 = ~n43246 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n25032 = ~n25028 | ~n25027;
  assign n25030 = ~n43274 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n25029 = ~n43265 | ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n25031 = ~n25030 | ~n25029;
  assign n25040 = ~n25032 & ~n25031;
  assign n25034 = ~n28775 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n25033 = ~n43242 | ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n25038 = ~n25034 | ~n25033;
  assign n25036 = ~n43261 | ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n25035 = ~n43264 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n25037 = ~n25036 | ~n25035;
  assign n25039 = ~n25038 & ~n25037;
  assign n25056 = ~n25040 | ~n25039;
  assign n25042 = ~n43260 | ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n25041 = ~n22915 | ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n25046 = ~n25042 | ~n25041;
  assign n25044 = ~n43270 | ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n25043 = ~n43275 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n25045 = ~n25044 | ~n25043;
  assign n25054 = ~n25046 & ~n25045;
  assign n25048 = ~n43245 | ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n25047 = ~n43251 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n25052 = ~n25048 | ~n25047;
  assign n25050 = ~n22908 | ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n25049 = ~n43271 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n25051 = ~n25050 | ~n25049;
  assign n25053 = ~n25052 & ~n25051;
  assign n25055 = ~n25054 | ~n25053;
  assign n25057 = ~n25056 & ~n25055;
  assign n25058 = ~n28608 | ~P1_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n25067 = ~n25850;
  assign n25070 = ~n34149 & ~n32238;
  assign n31904 = n31927 | n31447;
  assign n25075 = ~n25074 & ~n25073;
  assign n35626 = ~n44102;
  assign n43300 = ~n25075 & ~n35626;
  assign n43298 = ~n43300 | ~n39892;
  assign n25090 = ~n38662 | ~n44021;
  assign n25089 = ~P1_EBX_REG_12__SCAN_IN | ~n44023;
  assign n25091 = ~n25090 | ~n25089;
  assign P1_U2860 = n25092 | n25091;
  assign n25095 = ~n23127 & ~n25093;
  assign n25098 = ~n25097 & ~n25096;
  assign n25100 = ~n25099 & ~n25098;
  assign n41759 = ~n25100 & ~n32149;
  assign n25101 = ~n22904 & ~n36688;
  assign n25104 = ~BUF2_REG_19__SCAN_IN | ~n43689;
  assign n43690 = ~n25102 & ~n36558;
  assign n25103 = ~BUF1_REG_19__SCAN_IN | ~n43690;
  assign n25800 = ~n25104 | ~n25103;
  assign n25112 = ~n25106 | ~n25105;
  assign n25108 = ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n25111 = ~n25110 & ~n25109;
  assign n25117 = ~n26831 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n25116 = ~n26858 | ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n25119 = ~n26837 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n25118 = ~n26841 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n25123 = ~n26726 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n25122 = ~n26838 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n25127 = ~n25123 | ~n25122;
  assign n25125 = ~n22906 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n25124 = ~n26832 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n25126 = ~n25125 | ~n25124;
  assign n25377 = ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n25132 = ~n26807 & ~n25377;
  assign n25130 = ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n25131 = ~n26808 & ~n25130;
  assign n25136 = ~n25132 & ~n25131;
  assign n25134 = ~n26789 & ~n39534;
  assign n25133 = ~n26791 & ~n37629;
  assign n25135 = ~n25134 & ~n25133;
  assign n25138 = ~n26852 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n25137 = ~n26827 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n26891 = ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n25142 = ~n26780 & ~n26891;
  assign n25360 = ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n25141 = ~n22905 & ~n25360;
  assign n25717 = n25146 | n25145;
  assign n34646 = ~n35253 & ~n33915;
  assign n25150 = ~n26848 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n25148 = ~n26789 & ~n41578;
  assign n25147 = ~n26791 & ~n41597;
  assign n25149 = ~n25148 & ~n25147;
  assign n25154 = ~n25150 | ~n25149;
  assign n25152 = ~n26852 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n25151 = ~n22926 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n25153 = ~n25152 | ~n25151;
  assign n25156 = ~n26831 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n25155 = ~n22906 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n25158 = ~n26837 | ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n25157 = ~n26827 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n25164 = ~n25656 & ~n26257;
  assign n25499 = ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n25163 = ~n25653 & ~n25499;
  assign n25170 = ~n25164 & ~n25163;
  assign n25168 = ~n25652 & ~n41592;
  assign n25166 = ~n26859 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n25165 = ~n23481 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n25172 = ~n26832 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n25171 = ~n26841 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n25178 = ~n26831 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n25177 = ~n26726 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n25180 = ~n26852 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n25179 = ~n26838 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n25184 = ~n26837 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n25183 = ~n26841 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n25186 = ~n26849 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n25185 = ~n26859 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n25424 = ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n25192 = ~n26807 & ~n25424;
  assign n25191 = ~n26791 & ~n37739;
  assign n25194 = ~n25192 & ~n25191;
  assign n25193 = ~n26858 | ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n41648 = ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n25195 = ~n26780 & ~n41648;
  assign n25198 = ~n26848 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n25197 = ~n26827 | ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n25200 = ~n22906 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n25199 = ~n26832 | ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n25201 = ~n25200 | ~n25199;
  assign n25731 = n25206 | n25205;
  assign n41804 = ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n25208 = ~n25495 & ~n41804;
  assign n25469 = ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n25207 = ~n22905 & ~n25469;
  assign n25214 = ~n25208 & ~n25207;
  assign n41822 = ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n25212 = ~n26780 & ~n41822;
  assign n25210 = ~n26859 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n25209 = ~n23481 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n25211 = ~n25210 | ~n25209;
  assign n25213 = ~n25212 & ~n25211;
  assign n25216 = ~n26852 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n25215 = ~n26827 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n25220 = ~n25216 | ~n25215;
  assign n25218 = ~n26832 | ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n25217 = ~n22906 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n25219 = ~n25218 | ~n25217;
  assign n25221 = n25220 | n25219;
  assign n25224 = ~n26849 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n25223 = ~n26862 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n25226 = ~n25224 | ~n25223;
  assign n25225 = ~n25653 & ~n41805;
  assign n25230 = ~n25226 & ~n25225;
  assign n25228 = ~n26726 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n25227 = ~n26858 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n25229 = n25228 & n25227;
  assign n25232 = ~n26837 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n25231 = ~n26841 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n25238 = ~n22906 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n25237 = ~n26828 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n25242 = ~n25238 | ~n25237;
  assign n25240 = ~n26841 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n25239 = ~n26859 | ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n25244 = ~n26831 | ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n25243 = ~n26832 | ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n25248 = ~n25244 | ~n25243;
  assign n25246 = ~n22926 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n25245 = ~n26849 | ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n25247 = ~n25246 | ~n25245;
  assign n25252 = ~n26807 & ~n42786;
  assign n25251 = ~n26791 & ~n42782;
  assign n25254 = ~n25252 & ~n25251;
  assign n25253 = ~n26837 | ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n25256 = ~n26852 | ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n25255 = ~n26827 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n25260 = ~n26838 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n25259 = ~n26858 | ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n25262 = ~n25260 | ~n25259;
  assign n25261 = ~n22905 & ~n42783;
  assign n25263 = ~n25262 & ~n25261;
  assign n25745 = n25266 | n25265;
  assign n25268 = ~n22926 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n25267 = ~n26832 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n25272 = ~n25268 | ~n25267;
  assign n25270 = ~n22906 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n25269 = ~n26827 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n25271 = ~n25270 | ~n25269;
  assign n25282 = n25272 | n25271;
  assign n25274 = ~n26837 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n25273 = ~n26852 | ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n25280 = n25274 & n25273;
  assign n25276 = ~n26849 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n25275 = ~n23481 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n25278 = ~n25276 | ~n25275;
  assign n25277 = ~n22905 & ~n43093;
  assign n25279 = ~n25278 & ~n25277;
  assign n25284 = ~n25656 & ~n26779;
  assign n25283 = ~n25652 & ~n43099;
  assign n25291 = ~n25284 & ~n25283;
  assign n25289 = ~n25653 & ~n25285;
  assign n25287 = ~n26862 | ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n25286 = ~n26859 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n25288 = ~n25287 | ~n25286;
  assign n25290 = ~n25289 & ~n25288;
  assign n25293 = ~n26831 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n25292 = ~n26841 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n25294 = ~n25293 | ~n25292;
  assign n25299 = ~n26827 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n25298 = ~n26841 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n25303 = ~n25299 | ~n25298;
  assign n25301 = ~n26848 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n25300 = ~n22906 | ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n25302 = ~n25301 | ~n25300;
  assign n25311 = ~n25303 & ~n25302;
  assign n25305 = ~n26831 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n25304 = ~n26858 | ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n25309 = ~n25305 | ~n25304;
  assign n25307 = ~n22926 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n25306 = ~n23481 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n25308 = ~n25307 | ~n25306;
  assign n25310 = ~n25309 & ~n25308;
  assign n43425 = ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n25314 = ~n26789 & ~n43425;
  assign n25312 = ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n25313 = ~n26808 & ~n25312;
  assign n25316 = ~n25314 & ~n25313;
  assign n25315 = ~n26838 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n25320 = ~n25316 | ~n25315;
  assign n25318 = ~n26837 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n25317 = ~n26832 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n25319 = ~n25318 | ~n25317;
  assign n25326 = ~n25320 & ~n25319;
  assign n25324 = ~n25634 & ~n26396;
  assign n25322 = ~n26828 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n25321 = ~n26862 | ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n25323 = ~n25322 | ~n25321;
  assign n25325 = ~n25324 & ~n25323;
  assign n25759 = n25328 | n25327;
  assign n25330 = ~n26848 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n25329 = ~n26831 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n25334 = ~n25330 | ~n25329;
  assign n25332 = ~n26837 | ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n25331 = ~n22906 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n25333 = ~n25332 | ~n25331;
  assign n25344 = ~n25334 & ~n25333;
  assign n25336 = ~n26789 & ~n43512;
  assign n25335 = ~n26808 & ~n25676;
  assign n25338 = ~n25336 & ~n25335;
  assign n25337 = ~n26852 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n25342 = ~n25338 | ~n25337;
  assign n25340 = ~n22926 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n25339 = ~n26841 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n25341 = ~n25340 | ~n25339;
  assign n25343 = ~n25342 & ~n25341;
  assign n25359 = n25344 & n25343;
  assign n25345 = ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n25349 = ~n25656 & ~n25345;
  assign n25347 = ~n26862 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n25346 = ~n23481 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n25348 = ~n25347 | ~n25346;
  assign n25353 = ~n25349 & ~n25348;
  assign n25351 = ~n26838 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n25350 = ~n26858 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n25352 = n25351 & n25350;
  assign n25357 = ~n25353 | ~n25352;
  assign n25355 = ~n26827 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n25354 = ~n26832 | ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n25356 = ~n25355 | ~n25354;
  assign n25358 = ~n25357 & ~n25356;
  assign n25362 = ~n26807 & ~n25360;
  assign n25361 = ~n26808 & ~n39534;
  assign n25364 = ~n25362 & ~n25361;
  assign n25363 = ~n22926 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n25368 = ~n25364 | ~n25363;
  assign n25366 = ~n26848 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n25365 = ~n26841 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n25367 = ~n25366 | ~n25365;
  assign n25376 = ~n25368 & ~n25367;
  assign n25370 = ~n26852 | ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n25369 = ~n26837 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n25374 = ~n25370 | ~n25369;
  assign n25372 = ~n22906 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n25371 = ~n26827 | ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n25373 = ~n25372 | ~n25371;
  assign n25375 = ~n25374 & ~n25373;
  assign n25391 = ~n25376 | ~n25375;
  assign n25379 = ~n26789 & ~n37629;
  assign n25378 = ~n26791 & ~n25377;
  assign n25381 = ~n25379 & ~n25378;
  assign n25380 = ~n26726 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n25385 = ~n25381 | ~n25380;
  assign n25383 = ~n26838 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n25382 = ~n26858 | ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n25384 = ~n25383 | ~n25382;
  assign n25389 = ~n25385 & ~n25384;
  assign n25387 = ~n26831 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n25386 = ~n26832 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n25388 = n25387 & n25386;
  assign n25390 = ~n25389 | ~n25388;
  assign n37442 = ~n37120 & ~n37119;
  assign n25393 = ~n26837 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n25392 = ~n26831 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n25397 = ~n25393 | ~n25392;
  assign n25395 = ~n26841 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n25394 = ~n26838 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n25396 = ~n25395 | ~n25394;
  assign n25405 = ~n25397 & ~n25396;
  assign n25399 = ~n22906 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n25398 = ~n26858 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n25403 = ~n25399 | ~n25398;
  assign n25401 = ~n26827 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n25400 = ~n26726 | ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n25402 = ~n25401 | ~n25400;
  assign n25404 = ~n25403 & ~n25402;
  assign n25421 = ~n25405 | ~n25404;
  assign n41601 = ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n25407 = ~n26807 & ~n41601;
  assign n25406 = ~n26789 & ~n41597;
  assign n25411 = ~n25407 & ~n25406;
  assign n41591 = ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n25409 = ~n26791 & ~n41591;
  assign n25408 = ~n26808 & ~n41578;
  assign n25410 = ~n25409 & ~n25408;
  assign n25415 = ~n25411 | ~n25410;
  assign n25413 = ~n26852 | ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n25412 = ~n26832 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n25414 = ~n25413 | ~n25412;
  assign n25419 = ~n25415 & ~n25414;
  assign n25417 = ~n26780 & ~n26257;
  assign n25416 = ~n22905 & ~n41588;
  assign n25418 = ~n25417 & ~n25416;
  assign n25420 = ~n25419 | ~n25418;
  assign n37441 = n25421 | n25420;
  assign n25423 = ~n26848 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n25422 = ~n26831 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n25430 = ~n25423 | ~n25422;
  assign n25426 = ~n26789 & ~n37739;
  assign n25425 = ~n26791 & ~n25424;
  assign n25428 = ~n25426 & ~n25425;
  assign n25427 = ~n26852 | ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n25429 = ~n25428 | ~n25427;
  assign n25438 = ~n25430 & ~n25429;
  assign n25432 = ~n22926 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n25431 = ~n22906 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n25436 = ~n25432 | ~n25431;
  assign n25434 = ~n26827 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n25433 = ~n26832 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n25435 = ~n25434 | ~n25433;
  assign n25437 = ~n25436 & ~n25435;
  assign n25454 = ~n25438 | ~n25437;
  assign n25439 = ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n25442 = ~n26807 & ~n25439;
  assign n25441 = ~n26808 & ~n25440;
  assign n25444 = ~n25442 & ~n25441;
  assign n25443 = ~n26828 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n25448 = ~n25444 | ~n25443;
  assign n25446 = ~n26858 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n25445 = ~n26838 | ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n25447 = ~n25446 | ~n25445;
  assign n25452 = ~n25448 & ~n25447;
  assign n25450 = ~n26837 | ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n25449 = ~n26841 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n25451 = n25450 & n25449;
  assign n25453 = ~n25452 | ~n25451;
  assign n25456 = ~n26832 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n25455 = ~n26828 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n25460 = ~n25456 | ~n25455;
  assign n25458 = ~n26827 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n25457 = ~n26858 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n25459 = ~n25458 | ~n25457;
  assign n25468 = ~n25460 & ~n25459;
  assign n25462 = ~n26831 | ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n25461 = ~n22906 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n25466 = ~n25462 | ~n25461;
  assign n25464 = ~n26841 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n25463 = ~n26838 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n25465 = ~n25464 | ~n25463;
  assign n25467 = ~n25466 & ~n25465;
  assign n25486 = ~n25468 | ~n25467;
  assign n25471 = ~n26807 & ~n25469;
  assign n25470 = ~n26808 & ~n26301;
  assign n25475 = ~n25471 & ~n25470;
  assign n25473 = ~n26789 & ~n37796;
  assign n41821 = ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n25472 = ~n26791 & ~n41821;
  assign n25474 = ~n25473 & ~n25472;
  assign n25479 = ~n25475 | ~n25474;
  assign n25477 = ~n26837 | ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n25476 = ~n26852 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n25478 = ~n25477 | ~n25476;
  assign n25484 = ~n25479 & ~n25478;
  assign n26288 = ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n25482 = ~n26780 & ~n26288;
  assign n25480 = ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n25481 = ~n22905 & ~n25480;
  assign n25483 = ~n25482 & ~n25481;
  assign n25485 = ~n25484 | ~n25483;
  assign n25488 = n25486 | n25485;
  assign n25489 = ~n25488;
  assign n41754 = ~n41759 | ~n25491;
  assign n25497 = ~n25495 & ~n26232;
  assign n25496 = ~n26818 & ~n26257;
  assign n25498 = ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n25501 = ~n25641 & ~n25498;
  assign n25500 = ~n25687 & ~n25499;
  assign n25505 = ~n25634 & ~n41601;
  assign n25504 = ~n26820 & ~n41598;
  assign n25514 = ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n25516 = ~n25653 & ~n25514;
  assign n25515 = ~n25656 & ~n41602;
  assign n25520 = ~n25652 & ~n41588;
  assign n25531 = ~n41873 & ~P2_STATE2_REG_3__SCAN_IN;
  assign n25550 = ~n25532 | ~n25531;
  assign n25536 = ~n25550 & ~n29550;
  assign n25553 = ~n25540 & ~n25539;
  assign n32168 = ~n25541 & ~n25553;
  assign n25542 = ~P2_STATE2_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n26914 = ~n28191;
  assign n41473 = ~n25550;
  assign n32890 = ~n25572 | ~n25566;
  assign n25567 = ~P2_EAX_REG_2__SCAN_IN;
  assign n36831 = ~n25587 | ~n25586;
  assign n25588 = ~P2_EAX_REG_4__SCAN_IN;
  assign n25594 = ~n26807 & ~n43091;
  assign n25593 = ~n26791 & ~n26768;
  assign n25598 = ~n26838 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n25597 = ~n26858 | ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n25602 = ~n26818 & ~n26779;
  assign n25601 = ~n26820 & ~n43086;
  assign n25607 = ~n26789 & ~n25605;
  assign n43072 = ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n25606 = ~n26808 & ~n43072;
  assign n25609 = ~n25607 & ~n25606;
  assign n25608 = ~n26848 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n25610 = ~n22926 | ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n36829 = ~n25625 | ~n25624;
  assign n25633 = ~n22905 & ~n26790;
  assign n25631 = ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n25638 = ~n25634 & ~n26806;
  assign n25643 = ~n25641 & ~n26819;
  assign n43409 = ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n25642 = ~n26820 & ~n43409;
  assign n25647 = ~n26818 & ~n25644;
  assign n26817 = ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n25646 = ~n25645 & ~n26817;
  assign n25655 = ~n25652 & ~n26396;
  assign n25654 = ~n25653 & ~n43426;
  assign n43407 = ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n26552 = ~n25670 | ~n25669;
  assign n25712 = ~n26552 | ~n26551;
  assign n25679 = ~n26726 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n25694 = ~n26807 & ~n37805;
  assign n25693 = ~n26808 & ~n25692;
  assign n42353 = ~n25710 & ~n25709;
  assign n43835 = ~n42353;
  assign n32345 = ~n25712 | ~n25711;
  assign n31210 = ~P2_EAX_REG_7__SCAN_IN;
  assign n25740 = ~n26914 & ~n42104;
  assign n33784 = ~n33556 & ~n33555;
  assign n34836 = ~n33784 | ~n33783;
  assign n42100 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n25753 = ~n26914 & ~n42100;
  assign n31223 = ~P2_EAX_REG_13__SCAN_IN;
  assign n25752 = ~n26916 & ~n31223;
  assign n35378 = ~n34836 & ~n34835;
  assign n25760 = ~n28191 | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n35376 = ~n35378 | ~n35377;
  assign n25767 = ~n26914 & ~n42215;
  assign n31268 = ~P2_EAX_REG_15__SCAN_IN;
  assign n25766 = ~n26916 & ~n31268;
  assign n37124 = ~n35376 & ~n35316;
  assign n25774 = ~n26914 & ~n42628;
  assign n25772 = ~P2_EAX_REG_16__SCAN_IN;
  assign n25773 = ~n26916 & ~n25772;
  assign n37445 = ~n37124 | ~n37123;
  assign n25778 = ~n41474 | ~P2_EAX_REG_17__SCAN_IN;
  assign n25777 = ~n28191 | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n36375 = ~n37445 & ~n37444;
  assign n25783 = ~n26914 & ~n42282;
  assign n25781 = ~P2_EAX_REG_18__SCAN_IN;
  assign n25782 = ~n26916 & ~n25781;
  assign n25787 = ~n41474 | ~P2_EAX_REG_19__SCAN_IN;
  assign n25786 = ~n28191 | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n43695 = ~n41759 | ~n22904;
  assign n25790 = ~n22904 & ~n41873;
  assign n25792 = ~BUF2_REG_3__SCAN_IN | ~n36558;
  assign n25791 = ~n36557 | ~BUF1_REG_3__SCAN_IN;
  assign n36792 = ~n25792 | ~n25791;
  assign n36001 = ~n36792;
  assign n25794 = ~n43697 & ~n36001;
  assign n31214 = ~P2_EAX_REG_19__SCAN_IN;
  assign n25793 = ~n41759 & ~n31214;
  assign n25795 = ~n25794 & ~n25793;
  assign n25799 = n25798 | n25797;
  assign P2_U2900 = n25800 | n25799;
  assign n25802 = ~n43270 | ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n25801 = ~n43260 | ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n25806 = ~n25802 | ~n25801;
  assign n25804 = ~n43245 | ~P1_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n25803 = ~n22908 | ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n25805 = ~n25804 | ~n25803;
  assign n25814 = ~n25806 & ~n25805;
  assign n25808 = ~n43275 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n25807 = ~n43261 | ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n25812 = ~n25808 | ~n25807;
  assign n25810 = ~n43264 | ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n25809 = ~n43265 | ~P1_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n25811 = ~n25810 | ~n25809;
  assign n25813 = ~n25812 & ~n25811;
  assign n25830 = ~n25814 | ~n25813;
  assign n25816 = ~n43246 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n25815 = ~n43251 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n25820 = ~n25816 | ~n25815;
  assign n25818 = ~n43274 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n25817 = ~n43242 | ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n25819 = ~n25818 | ~n25817;
  assign n25828 = ~n25820 & ~n25819;
  assign n25822 = ~n22907 | ~P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n25821 = ~n43241 | ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n25826 = ~n25822 | ~n25821;
  assign n25824 = ~n22915 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n25823 = ~n43271 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n25825 = ~n25824 | ~n25823;
  assign n25827 = ~n25826 & ~n25825;
  assign n25829 = ~n25828 | ~n25827;
  assign n25831 = ~n25830 & ~n25829;
  assign n25835 = n22942 | n25831;
  assign n25832 = ~n28608 | ~P1_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n25848 = ~n40493 & ~n44019;
  assign n25846 = ~n40098 | ~n44021;
  assign n25845 = ~P1_EBX_REG_13__SCAN_IN | ~n44023;
  assign n25847 = ~n25846 | ~n25845;
  assign P1_U2859 = n25848 | n25847;
  assign n25852 = ~n43274 | ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n25851 = ~n43264 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n25856 = ~n25852 | ~n25851;
  assign n25854 = ~n43275 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n25853 = ~n22908 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n25855 = ~n25854 | ~n25853;
  assign n25864 = ~n25856 & ~n25855;
  assign n25858 = ~n43270 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n25857 = ~n22915 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n25862 = ~n25858 | ~n25857;
  assign n25860 = ~n43245 | ~P1_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n25859 = ~n43265 | ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n25861 = ~n25860 | ~n25859;
  assign n25863 = ~n25862 & ~n25861;
  assign n25880 = ~n25864 | ~n25863;
  assign n25866 = ~n43251 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n25865 = ~n43242 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n25870 = ~n25866 | ~n25865;
  assign n25868 = ~n43241 | ~P1_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n25867 = ~n43260 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n25869 = ~n25868 | ~n25867;
  assign n25878 = ~n25870 & ~n25869;
  assign n25872 = ~n22907 | ~P1_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n25871 = ~n43246 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n25876 = ~n25872 | ~n25871;
  assign n25874 = ~n43261 | ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n25873 = ~n43271 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n25875 = ~n25874 | ~n25873;
  assign n25877 = ~n25876 & ~n25875;
  assign n25879 = ~n25878 | ~n25877;
  assign n25881 = ~n25880 & ~n25879;
  assign n25888 = n22942 | n25881;
  assign n44034 = ~P1_EAX_REG_14__SCAN_IN;
  assign n25884 = ~n28810 & ~n44034;
  assign n25882 = ~P1_PHYADDRPOINTER_REG_14__SCAN_IN | ~n43722;
  assign n25883 = ~n43725 | ~n25882;
  assign n25887 = ~n25884 & ~n25883;
  assign n25886 = ~n41131 & ~n43725;
  assign n26084 = ~n25888 | ~n22938;
  assign n40709 = ~P1_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n25890 = ~P1_STATEBS16_REG_SCAN_IN | ~n40709;
  assign n25891 = ~n25890 | ~n43722;
  assign n25899 = ~n28775 | ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n25898 = ~n43251 | ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n25903 = ~n25899 | ~n25898;
  assign n25901 = ~n43274 | ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n25900 = ~n22908 | ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n25902 = ~n25901 | ~n25900;
  assign n25911 = ~n25903 & ~n25902;
  assign n25905 = ~n43246 | ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n25904 = ~n43242 | ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n25909 = ~n25905 | ~n25904;
  assign n25907 = ~n43270 | ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n25906 = ~n43265 | ~P1_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n25908 = ~n25907 | ~n25906;
  assign n25910 = ~n25909 & ~n25908;
  assign n25913 = ~n22907 | ~P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n25912 = ~n43264 | ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n25917 = ~n25913 | ~n25912;
  assign n25915 = ~n43275 | ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n25914 = ~n22915 | ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n25916 = ~n25915 | ~n25914;
  assign n25925 = ~n25917 & ~n25916;
  assign n25919 = ~n43245 | ~P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n25918 = ~n43260 | ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n25923 = ~n25919 | ~n25918;
  assign n25921 = ~n43261 | ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n25920 = ~n43271 | ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n25922 = ~n25921 | ~n25920;
  assign n25924 = ~n25923 & ~n25922;
  assign n25929 = n25927 | n25926;
  assign n26569 = ~n25931 | ~n25930;
  assign n25949 = ~n40707 & ~n44019;
  assign n25945 = n25944 & n25943;
  assign n25947 = ~n40706 | ~n44021;
  assign n25946 = ~n44023 | ~P1_EBX_REG_15__SCAN_IN;
  assign P1_U2857 = n25949 | n25948;
  assign n38642 = ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n25957 = ~n38643 & ~n38642;
  assign n38641 = ~P1_INSTADDRPOINTER_REG_9__SCAN_IN | ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n39555 = ~n38641;
  assign n36889 = ~n25951;
  assign n36894 = ~n36889 & ~n25950;
  assign n38652 = ~n39555 | ~n36894;
  assign n38645 = n34279 | n38652;
  assign n38648 = ~n25952 | ~n25951;
  assign n25958 = ~n38648 & ~n38641;
  assign n25953 = ~n36891 | ~n25958;
  assign n28539 = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN | ~P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n25981 = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n40091 = ~P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n25954 = ~n25981 | ~n40091;
  assign n25955 = ~n28539 | ~n25954;
  assign n25991 = ~n40088 & ~n25955;
  assign n25956 = ~n25957;
  assign n28545 = ~n25956 & ~n38652;
  assign n25961 = ~n36895 & ~n28545;
  assign n28541 = ~n25958 | ~n25957;
  assign n25959 = ~n36891 | ~n28541;
  assign n25960 = ~n36893 | ~n25959;
  assign n25989 = n40092 | n25981;
  assign n25964 = ~n25962;
  assign n25966 = ~n25964 | ~n25963;
  assign n25969 = ~n36904 | ~n36905;
  assign n25967 = ~P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n38799 = ~n25969 | ~n25968;
  assign n25974 = ~n38799 | ~n25970;
  assign n38384 = ~n25974 | ~n25973;
  assign n40093 = ~n38384 | ~n25976;
  assign n25980 = ~n40093 | ~n25978;
  assign n26565 = ~n25980 | ~n25979;
  assign n25982 = ~n26566 | ~n26564;
  assign n40786 = ~n43469 | ~P1_REIP_REG_14__SCAN_IN;
  assign P1_U3017 = n25991 | n25990;
  assign n25994 = ~P1_PHYADDRPOINTER_REG_16__SCAN_IN | ~n43722;
  assign n25997 = ~n43246 | ~P1_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n25996 = ~n43242 | ~P1_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n26001 = ~n25997 | ~n25996;
  assign n25999 = ~n28775 | ~P1_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n25998 = ~n43274 | ~P1_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n26000 = ~n25999 | ~n25998;
  assign n26009 = ~n26001 & ~n26000;
  assign n26003 = ~n22907 | ~P1_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n26002 = ~n43251 | ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n26007 = ~n26003 | ~n26002;
  assign n26005 = ~n22908 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n26004 = ~n22915 | ~P1_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n26006 = ~n26005 | ~n26004;
  assign n26008 = ~n26007 & ~n26006;
  assign n26025 = ~n26009 | ~n26008;
  assign n26011 = ~n43245 | ~P1_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n26010 = ~n43275 | ~P1_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n26015 = ~n26011 | ~n26010;
  assign n26013 = ~n43261 | ~P1_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n26012 = ~n43265 | ~P1_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n26014 = ~n26013 | ~n26012;
  assign n26023 = ~n26015 & ~n26014;
  assign n26017 = ~n43270 | ~P1_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n26016 = ~n43264 | ~P1_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n26021 = ~n26017 | ~n26016;
  assign n26019 = ~n43260 | ~P1_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n26018 = ~n43271 | ~P1_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n26020 = ~n26019 | ~n26018;
  assign n26022 = ~n26021 & ~n26020;
  assign n26024 = ~n26023 | ~n26022;
  assign n26026 = ~n26025 & ~n26024;
  assign n43286 = ~n31921 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n26027 = n26026 | n43286;
  assign n26037 = ~n44023 | ~P1_EBX_REG_16__SCAN_IN;
  assign P1_U2856 = n26040 | n26039;
  assign n37237 = ~P1_REIP_REG_8__SCAN_IN;
  assign n35875 = ~P1_REIP_REG_3__SCAN_IN;
  assign n35877 = ~P1_REIP_REG_1__SCAN_IN | ~P1_REIP_REG_2__SCAN_IN;
  assign n35501 = ~n35875 & ~n35877;
  assign n35502 = ~P1_REIP_REG_4__SCAN_IN | ~n35501;
  assign n26041 = ~P1_REIP_REG_6__SCAN_IN | ~P1_REIP_REG_5__SCAN_IN;
  assign n34829 = ~n35502 & ~n26041;
  assign n37235 = ~P1_REIP_REG_7__SCAN_IN | ~n34829;
  assign n26042 = ~n37237 & ~n37235;
  assign n37227 = ~P1_REIP_REG_9__SCAN_IN | ~n26042;
  assign n38256 = ~P1_REIP_REG_11__SCAN_IN | ~P1_REIP_REG_10__SCAN_IN;
  assign n26043 = ~n37227 & ~n38256;
  assign n26696 = ~P1_REIP_REG_12__SCAN_IN | ~n26043;
  assign n31717 = ~n31361 & ~n31898;
  assign n26045 = ~n26044;
  assign n42405 = ~n26065 & ~n26048;
  assign n26049 = ~n26696 & ~n42185;
  assign n26055 = ~n26049 | ~n40089;
  assign n26050 = ~P1_STATE2_REG_3__SCAN_IN | ~P1_STATE2_REG_0__SCAN_IN;
  assign n26586 = ~n33710 | ~P1_STATE2_REG_1__SCAN_IN;
  assign n44107 = n43725 | n26586;
  assign n26052 = ~n35624 & ~n26051;
  assign n26053 = ~n42405 | ~n26696;
  assign n38253 = ~n41894 | ~n26053;
  assign n26054 = ~P1_REIP_REG_13__SCAN_IN | ~n38253;
  assign n26083 = ~n26055 | ~n26054;
  assign n34514 = ~P1_STATEBS16_REG_SCAN_IN & ~n44100;
  assign n43803 = n26057 & n31793;
  assign n28885 = ~P1_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n26077 = ~n40490 | ~n43559;
  assign n26070 = ~n26065;
  assign n26066 = ~P1_EBX_REG_31__SCAN_IN;
  assign n26067 = ~n31382 | ~n26066;
  assign n26068 = ~n31715 | ~n26067;
  assign n26072 = ~n43796;
  assign n26071 = ~P1_EBX_REG_13__SCAN_IN;
  assign n26075 = ~n26072 & ~n26071;
  assign n41129 = ~n41894 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n26073 = ~P1_PHYADDRPOINTER_REG_13__SCAN_IN | ~n43797;
  assign n26074 = ~n43033 | ~n26073;
  assign n26076 = ~n26075 & ~n26074;
  assign P1_U2827 = n26083 | n26082;
  assign n26088 = ~n41127 | ~n44021;
  assign n26087 = ~n44023 | ~P1_EBX_REG_14__SCAN_IN;
  assign n26089 = ~n26088 | ~n26087;
  assign P1_U2858 = n26090 | n26089;
  assign n26098 = ~n26095 & ~n26094;
  assign n26097 = ~n27006 & ~n26096;
  assign n26104 = ~n26098 & ~n26097;
  assign n26102 = ~n27009 & ~n26099;
  assign n26101 = ~n28587 & ~n26100;
  assign n26103 = ~n26102 & ~n26101;
  assign n26108 = ~n26104 | ~n26103;
  assign n26106 = ~n43245 | ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n26105 = ~n43265 | ~P1_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n26107 = ~n26106 | ~n26105;
  assign n26128 = ~n26108 & ~n26107;
  assign n26110 = ~n43241 | ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n26109 = ~n43251 | ~P1_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n26114 = ~n26110 | ~n26109;
  assign n26112 = ~n43275 | ~P1_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n26111 = ~n43242 | ~P1_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n26113 = ~n26112 | ~n26111;
  assign n26122 = ~n26114 & ~n26113;
  assign n26116 = ~n22907 | ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n26115 = ~n43246 | ~P1_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n26120 = ~n26116 | ~n26115;
  assign n26118 = ~n43261 | ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n26117 = ~n22915 | ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n26119 = ~n26118 | ~n26117;
  assign n26121 = ~n26120 & ~n26119;
  assign n26126 = ~n26122 | ~n26121;
  assign n26124 = ~n43274 | ~P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n26123 = ~n43264 | ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n26125 = ~n26124 | ~n26123;
  assign n26127 = ~n26126 & ~n26125;
  assign n26129 = ~n26128 | ~n26127;
  assign n31983 = ~P1_EAX_REG_17__SCAN_IN;
  assign n26132 = ~n28810 & ~n31983;
  assign n26130 = ~P1_PHYADDRPOINTER_REG_17__SCAN_IN & ~n39944;
  assign n26131 = ~P1_STATE2_REG_2__SCAN_IN & ~n26130;
  assign n26133 = ~n26132 & ~n26131;
  assign n26140 = ~n26712;
  assign n26147 = ~n26142 | ~n26141;
  assign n26149 = ~n44023 | ~P1_EBX_REG_17__SCAN_IN;
  assign P1_U2855 = n26152 | n26151;
  assign n26156 = ~n26174 | ~n26153;
  assign n26155 = ~n26154 | ~n31055;
  assign n26161 = ~n26156 | ~n26155;
  assign n26158 = ~n26161 | ~n26157;
  assign n26160 = ~n26158 | ~n31055;
  assign n26166 = ~n26160 & ~n26159;
  assign n26162 = ~n26161;
  assign n26164 = ~n26162 & ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n26163 = ~n26174 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n26165 = ~n26164 & ~n26163;
  assign n26169 = n26168 | n26167;
  assign n26170 = ~n26174 | ~n35718;
  assign n26176 = n26173 | n26172;
  assign n26175 = ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n26174;
  assign n35801 = n32177 | n26178;
  assign n27870 = ~n26179 | ~n26200;
  assign n26187 = ~n36561 & ~n35802;
  assign n26186 = ~n31819 | ~n23127;
  assign n26188 = ~n26187 | ~n26186;
  assign n26190 = ~n31770 & ~n26188;
  assign n26194 = ~n26466;
  assign n31764 = ~n26200 | ~n28196;
  assign n26215 = ~n26206 | ~n35805;
  assign n26208 = ~n26207 | ~n31522;
  assign n43159 = ~n26550 | ~n26211;
  assign n42699 = ~n26550 | ~n31768;
  assign n26220 = ~n39656 & ~n39651;
  assign n26217 = ~n42600 & ~n26220;
  assign n34863 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n34859 = ~n34863 & ~n34858;
  assign n36601 = ~n34859;
  assign n26219 = ~n36840 & ~n36601;
  assign n26213 = ~n43159 & ~n26219;
  assign n35796 = ~n34863;
  assign n36600 = ~n35796 & ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n26218 = ~n36600 & ~n36840;
  assign n26212 = ~n42699 & ~n26218;
  assign n26216 = ~n26213 & ~n26212;
  assign n26561 = ~n28061 & ~n40770;
  assign n28067 = ~n26218 | ~n26220;
  assign n26222 = ~n42699 & ~n28067;
  assign n28065 = ~n26220 | ~n26219;
  assign n26221 = ~n43159 & ~n28065;
  assign n40767 = n26222 | n26221;
  assign n26272 = ~n26235 & ~n37279;
  assign n26229 = ~n38820 | ~n26272;
  assign n37654 = ~n26229 & ~n40306;
  assign n26230 = ~n37654 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n26234 = ~n26230 | ~n23127;
  assign n26231 = ~n38820 & ~n37302;
  assign n26258 = ~n40306 & ~n34876;
  assign n26364 = ~n26231 | ~n26258;
  assign n26247 = ~n26234 & ~n26233;
  assign n26236 = ~n26235;
  assign n26270 = ~n26236 & ~n37279;
  assign n26237 = ~n36607 | ~n26270;
  assign n37039 = ~n26237 & ~n40306;
  assign n26238 = ~n36607 | ~n26272;
  assign n38628 = ~n26238 & ~n40306;
  assign n26266 = ~n36607 | ~n40306;
  assign n26253 = ~n37302 | ~n37279;
  assign n26243 = ~n37965 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n26241 = ~n38820 | ~n26270;
  assign n36569 = ~n26241 & ~n40306;
  assign n26242 = ~n36569 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n26244 = ~n26243 | ~n26242;
  assign n26246 = ~n26245 & ~n26244;
  assign n26252 = ~n26247 | ~n26246;
  assign n26248 = ~n26258 | ~n38820;
  assign n37612 = ~n26248 & ~n35790;
  assign n26249 = ~n38237 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n26281 = ~n26252 & ~n26251;
  assign n26265 = n38820 & n40306;
  assign n26375 = ~n26265 | ~n26272;
  assign n26256 = ~n26375 & ~n41598;
  assign n26365 = ~n26265 | ~n26254;
  assign n26255 = ~n26365 & ~n41592;
  assign n26264 = ~n26256 & ~n26255;
  assign n26374 = ~n26265 | ~n22946;
  assign n26262 = ~n26374 & ~n26257;
  assign n26259 = ~n38820 & ~n35790;
  assign n26354 = ~n26259 | ~n26258;
  assign n26261 = ~n26354 & ~n26260;
  assign n26263 = ~n26262 & ~n26261;
  assign n26279 = ~n26264 | ~n26263;
  assign n26371 = ~n26265 | ~n26270;
  assign n26269 = ~n26371 & ~n41602;
  assign n26273 = ~n26266;
  assign n26370 = ~n26273 | ~n22946;
  assign n26267 = ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n26268 = ~n26370 & ~n26267;
  assign n26277 = ~n26269 & ~n26268;
  assign n26361 = ~n26273 | ~n26270;
  assign n26275 = ~n26361 & ~n26271;
  assign n26353 = ~n26273 | ~n26272;
  assign n26274 = ~n26353 & ~n41578;
  assign n26276 = ~n26275 & ~n26274;
  assign n26278 = ~n26277 | ~n26276;
  assign n26280 = ~n26279 & ~n26278;
  assign n26284 = ~n26281 | ~n26280;
  assign n26287 = ~n26284 | ~n26283;
  assign n26335 = ~n26287 | ~n26286;
  assign n26290 = ~n26371 & ~n41822;
  assign n26289 = ~n26374 & ~n26288;
  assign n26296 = ~n26290 & ~n26289;
  assign n26291 = ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n26294 = ~n26375 & ~n26291;
  assign n26293 = ~n26292 & ~n41805;
  assign n26295 = ~n26294 & ~n26293;
  assign n26308 = ~n26296 | ~n26295;
  assign n26297 = ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n26300 = ~n26365 & ~n26297;
  assign n26299 = ~n26361 & ~n26298;
  assign n26306 = ~n26300 & ~n26299;
  assign n26304 = ~n26353 & ~n26301;
  assign n26303 = ~n26354 & ~n26302;
  assign n26305 = ~n26304 & ~n26303;
  assign n26307 = ~n26306 | ~n26305;
  assign n26326 = ~n26308 & ~n26307;
  assign n26309 = ~n36569 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n26314 = ~n26310 | ~n26309;
  assign n26311 = ~n37654 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n26313 = ~n26312 | ~n26311;
  assign n26316 = ~n26314 & ~n26313;
  assign n26315 = ~n37612 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n26324 = ~n26316 | ~n26315;
  assign n26320 = ~n26370 & ~n26317;
  assign n26318 = ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n26319 = ~n26364 & ~n26318;
  assign n26322 = ~n26320 & ~n26319;
  assign n26321 = ~n38237 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n26325 = ~n26324 & ~n26323;
  assign n26329 = ~n26326 | ~n26325;
  assign n26333 = ~n26329 | ~n26328;
  assign n36485 = n26335 ^ n26333;
  assign n26336 = ~n26332 & ~n26331;
  assign n26334 = ~n26333;
  assign n26342 = ~n26335 | ~n26334;
  assign n26337 = ~n26342 ^ n26341;
  assign n26387 = ~n26340 | ~n36859;
  assign n26344 = ~n26392 & ~n43097;
  assign n26343 = ~n26397 & ~n43082;
  assign n39523 = ~n26353;
  assign n26357 = ~n26405 & ~n43093;
  assign n26359 = ~n26358 & ~n26357;
  assign n26366 = ~n38329 | ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n26381 = ~n26369 & ~n26368;
  assign n26372 = ~n37139 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n26377 = ~n39125 | ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n26376 = ~n36746 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n26378 = ~n26377 | ~n26376;
  assign n26380 = ~n26379 & ~n26378;
  assign n26382 = ~n26381 | ~n26380;
  assign n26386 = ~n26383 & ~n26382;
  assign n38376 = n26387 ^ n26432;
  assign n26388 = ~n26387 | ~n26432;
  assign n27855 = ~n26389 | ~n26388;
  assign n26420 = ~n36746 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n26430 = ~n26427 & ~n26426;
  assign n26433 = ~n26432;
  assign n26452 = ~n26433 & ~n43835;
  assign n26435 = ~n23322 | ~P2_EBX_REG_3__SCAN_IN;
  assign n26438 = ~n23322 | ~P2_EBX_REG_2__SCAN_IN;
  assign n26441 = ~n26440;
  assign n26442 = ~P2_EBX_REG_1__SCAN_IN & ~P2_EBX_REG_0__SCAN_IN;
  assign n26443 = ~n23322 | ~n26442;
  assign n26448 = ~n26445 & ~n23322;
  assign n26451 = ~n23322 | ~P2_EBX_REG_5__SCAN_IN;
  assign n26453 = ~n26452 & ~n40355;
  assign n26485 = ~n26453 & ~n39651;
  assign n26454 = ~n26453;
  assign n26455 = ~n26454 & ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n38373 = ~n26485 & ~n26455;
  assign n36488 = ~n26458 & ~n38821;
  assign n26473 = ~n26460 & ~n34858;
  assign n26461 = ~n40312 & ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n32943 = ~n26473 & ~n26461;
  assign n26465 = ~n26462;
  assign n26463 = ~P2_EBX_REG_0__SCAN_IN | ~P2_EBX_REG_1__SCAN_IN;
  assign n26464 = n41873 | n26463;
  assign n33569 = ~n26465 | ~n26464;
  assign n28119 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n26470 = ~n33569 & ~n28119;
  assign n26469 = ~n26466 & ~n23322;
  assign n26467 = ~P2_EBX_REG_0__SCAN_IN;
  assign n26468 = ~n41873 & ~n26467;
  assign n37290 = ~n26469 & ~n26468;
  assign n34880 = ~n37290 & ~n33579;
  assign n26472 = ~n26470 & ~n34880;
  assign n37310 = ~n33569;
  assign n26471 = ~n37310 & ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n32942 = ~n26472 & ~n26471;
  assign n26475 = ~n32943 | ~n32942;
  assign n26474 = ~n26473;
  assign n26480 = ~n26479 | ~n39656;
  assign n36853 = ~n26484 | ~n26480;
  assign n26481 = ~n36490 & ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n26482 = ~n36853 & ~n26481;
  assign n38374 = ~n38373 | ~n38372;
  assign n26491 = ~n26489 & ~n23322;
  assign n26502 = ~n27875 & ~n26501;
  assign n26504 = ~n26503 & ~n26502;
  assign n31772 = ~n26506 & ~n26505;
  assign n43755 = ~n26550 | ~n31772;
  assign n26556 = ~n40153 | ~n43876;
  assign n26510 = ~n31771 | ~n43061;
  assign n26511 = ~n26510 | ~n26509;
  assign n43886 = ~n26550 | ~n26511;
  assign n26517 = ~n26513 & ~n26512;
  assign n26524 = ~n39573 | ~P2_EBX_REG_4__SCAN_IN;
  assign n26523 = ~P2_PHYADDRPOINTER_REG_4__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n26532 = ~n39573 | ~P2_EBX_REG_5__SCAN_IN;
  assign n26531 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n26539 = ~n39573 | ~P2_EBX_REG_6__SCAN_IN;
  assign n26538 = ~P2_PHYADDRPOINTER_REG_6__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n40154 = n27894 ^ n27893;
  assign n26544 = ~n43767 | ~n40154;
  assign n40159 = ~n43880 | ~P2_REIP_REG_6__SCAN_IN;
  assign n26554 = ~n26544 | ~n40159;
  assign n26547 = ~n26546 | ~n26545;
  assign n26548 = ~n26547 | ~n23085;
  assign n26549 = ~n26548 | ~n31766;
  assign n43877 = ~n26550 | ~n26549;
  assign n39737 = ~n26552 ^ n26551;
  assign n26553 = ~n43877 & ~n39737;
  assign n26555 = ~n26554 & ~n26553;
  assign P2_U3040 = n26561 | n26560;
  assign n26562 = ~P1_INSTADDRPOINTER_REG_15__SCAN_IN & ~n28539;
  assign n26577 = ~n40795;
  assign n26563 = ~n28539 | ~n42539;
  assign n26567 = ~n26565 | ~n26564;
  assign n40704 = ~P1_REIP_REG_15__SCAN_IN;
  assign n40695 = ~n43033 & ~n40704;
  assign P1_U3016 = n26577 | n26576;
  assign n26583 = ~n26579 | ~n26578;
  assign n27822 = ~n26583 | ~n26582;
  assign n26584 = ~n43462 ^ n40798;
  assign n26597 = ~n40802 & ~n43358;
  assign n29569 = ~n26586 & ~n39944;
  assign n26595 = ~n41024 | ~n43367;
  assign n40803 = ~n43469 | ~P1_REIP_REG_16__SCAN_IN;
  assign n31468 = ~n26587 | ~n39946;
  assign n26588 = ~n31468 | ~n33710;
  assign n26589 = ~n43709 | ~P1_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n26593 = ~n40803 | ~n26589;
  assign n26590 = ~n33714 & ~P1_STATEBS16_REG_SCAN_IN;
  assign n31469 = ~P1_STATE2_REG_0__SCAN_IN & ~n43722;
  assign n31679 = ~n26590 & ~n31469;
  assign n26591 = ~n31679;
  assign n26592 = ~n43713 & ~n41025;
  assign n26594 = ~n26593 & ~n26592;
  assign P1_U2983 = n26597 | n26596;
  assign n26599 = ~P1_PHYADDRPOINTER_REG_18__SCAN_IN | ~n43722;
  assign n26602 = ~n43246 | ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n26601 = ~n43251 | ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n26606 = ~n26602 | ~n26601;
  assign n26604 = ~n43264 | ~P1_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n26603 = ~n43242 | ~P1_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n26605 = ~n26604 | ~n26603;
  assign n26614 = ~n26606 & ~n26605;
  assign n26608 = ~n22907 | ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n26607 = ~n28775 | ~P1_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n26612 = ~n26608 | ~n26607;
  assign n26610 = ~n22908 | ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n26609 = ~n43260 | ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n26611 = ~n26610 | ~n26609;
  assign n26613 = ~n26612 & ~n26611;
  assign n26630 = ~n26614 | ~n26613;
  assign n26616 = ~n43270 | ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n26615 = ~n43274 | ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n26620 = ~n26616 | ~n26615;
  assign n26618 = ~n43265 | ~P1_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n26617 = ~n43271 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n26619 = ~n26618 | ~n26617;
  assign n26628 = ~n26620 & ~n26619;
  assign n26622 = ~n43275 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n26621 = ~n22915 | ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n26626 = ~n26622 | ~n26621;
  assign n26624 = ~n43245 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n26623 = ~n43261 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n26625 = ~n26624 | ~n26623;
  assign n26627 = ~n26626 & ~n26625;
  assign n26629 = ~n26628 | ~n26627;
  assign n26631 = ~n26630 & ~n26629;
  assign n26632 = n26631 | n43286;
  assign n26635 = n26634 | n26633;
  assign n26639 = ~n43265 | ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n26638 = ~n22915 | ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n26643 = ~n26639 | ~n26638;
  assign n26641 = ~n43274 | ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n26640 = ~n43275 | ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n26642 = ~n26641 | ~n26640;
  assign n26670 = ~n26643 & ~n26642;
  assign n26645 = ~n28775 | ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n26644 = ~n43242 | ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n26649 = ~n26645 | ~n26644;
  assign n26647 = ~n22907 | ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n26646 = ~n43270 | ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n26648 = ~n26647 | ~n26646;
  assign n26657 = ~n26649 & ~n26648;
  assign n26651 = ~n43246 | ~P1_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n26650 = ~n43251 | ~P1_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n26655 = ~n26651 | ~n26650;
  assign n26653 = ~n43245 | ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n26652 = ~n43261 | ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n26654 = ~n26653 | ~n26652;
  assign n26656 = ~n26655 & ~n26654;
  assign n26668 = ~n26657 | ~n26656;
  assign n26661 = ~n27009 & ~n28592;
  assign n26660 = ~n26659 & ~n26658;
  assign n26666 = ~n26661 & ~n26660;
  assign n26664 = ~n27006 & ~n28586;
  assign n26663 = ~n28587 & ~n26662;
  assign n26665 = ~n26664 & ~n26663;
  assign n26667 = ~n26666 | ~n26665;
  assign n26669 = ~n26668 & ~n26667;
  assign n26671 = ~n26670 | ~n26669;
  assign n31973 = ~P1_EAX_REG_19__SCAN_IN;
  assign n26674 = ~n28810 & ~n31973;
  assign n26672 = ~P1_PHYADDRPOINTER_REG_19__SCAN_IN & ~n39944;
  assign n26673 = ~P1_STATE2_REG_2__SCAN_IN & ~n26672;
  assign n26675 = ~n26674 & ~n26673;
  assign n26682 = ~n28485;
  assign n26690 = ~n26715 | ~n26714;
  assign n26692 = ~n44023 | ~P1_EBX_REG_19__SCAN_IN;
  assign P1_U2853 = n26695 | n26694;
  assign n41125 = ~n40089 & ~n26696;
  assign n41020 = ~n40704 & ~n40703;
  assign n26697 = ~n42400 & ~n27836;
  assign n43566 = ~n42400 & ~n42405;
  assign n29613 = ~P1_REIP_REG_17__SCAN_IN;
  assign n26698 = ~n27836 & ~n42185;
  assign n26699 = ~P1_REIP_REG_17__SCAN_IN & ~n26698;
  assign n26710 = ~n41450 & ~n26699;
  assign n26701 = ~n43796 | ~P1_EBX_REG_17__SCAN_IN;
  assign n26700 = ~n43797 | ~P1_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n26709 = n26708 | n26707;
  assign P1_U2823 = n26710 | n26709;
  assign n26716 = ~n44023 | ~P1_EBX_REG_18__SCAN_IN;
  assign P1_U2854 = n26719 | n26718;
  assign n26721 = ~BUF2_REG_23__SCAN_IN | ~n43689;
  assign n26720 = ~BUF1_REG_23__SCAN_IN | ~n43690;
  assign n26942 = ~n26721 | ~n26720;
  assign n26723 = ~n26807 & ~n42783;
  assign n26722 = ~n26789 & ~n42782;
  assign n26725 = ~n26723 & ~n26722;
  assign n26724 = ~n26838 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n26730 = ~n26725 | ~n26724;
  assign n26728 = ~n26726 | ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n26727 = ~n26858 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n26729 = ~n26728 | ~n26727;
  assign n26734 = ~n26730 & ~n26729;
  assign n26732 = ~n26832 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n26731 = ~n26841 | ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n26733 = n26732 & n26731;
  assign n26753 = ~n26734 | ~n26733;
  assign n26736 = ~n26848 | ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n26735 = ~n26831 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n26743 = ~n26736 | ~n26735;
  assign n26739 = ~n26791 & ~n42786;
  assign n26738 = ~n26808 & ~n26737;
  assign n26741 = ~n26739 & ~n26738;
  assign n26740 = ~n22926 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n26742 = ~n26741 | ~n26740;
  assign n26751 = ~n26743 & ~n26742;
  assign n26745 = ~n26852 | ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n26744 = ~n26837 | ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n26749 = ~n26745 | ~n26744;
  assign n26747 = ~n22906 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n26746 = ~n26827 | ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n26748 = ~n26747 | ~n26746;
  assign n26750 = ~n26749 & ~n26748;
  assign n26752 = ~n26751 | ~n26750;
  assign n26755 = ~n22906 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n26754 = ~n26841 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n26759 = ~n26755 | ~n26754;
  assign n26757 = ~n26831 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n26756 = ~n26828 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n26758 = ~n26757 | ~n26756;
  assign n26767 = ~n26759 & ~n26758;
  assign n26761 = ~n26832 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n26760 = ~n26838 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n26765 = ~n26761 | ~n26760;
  assign n26763 = ~n26827 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n26762 = ~n26858 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n26764 = ~n26763 | ~n26762;
  assign n26766 = ~n26765 & ~n26764;
  assign n26786 = ~n26767 | ~n26766;
  assign n26770 = ~n26807 & ~n43093;
  assign n26769 = ~n26808 & ~n26768;
  assign n26774 = ~n26770 & ~n26769;
  assign n26772 = ~n26789 & ~n43091;
  assign n26771 = ~n26791 & ~n43097;
  assign n26773 = ~n26772 & ~n26771;
  assign n26778 = ~n26774 | ~n26773;
  assign n26776 = ~n26837 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n26775 = ~n26852 | ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n26777 = ~n26776 | ~n26775;
  assign n26784 = ~n26778 & ~n26777;
  assign n26782 = ~n26780 & ~n26779;
  assign n26781 = ~n22905 & ~n43082;
  assign n26783 = ~n26782 & ~n26781;
  assign n26785 = ~n26784 | ~n26783;
  assign n39670 = n26786 | n26785;
  assign n26788 = ~n26848 | ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n26787 = ~n26852 | ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n26797 = ~n26788 | ~n26787;
  assign n26793 = ~n26789 & ~n35254;
  assign n26792 = ~n26791 & ~n26790;
  assign n26795 = ~n26793 & ~n26792;
  assign n26794 = ~n22906 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n26796 = ~n26795 | ~n26794;
  assign n26805 = ~n26797 & ~n26796;
  assign n26799 = ~n22926 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n26798 = ~n26827 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n26803 = ~n26799 | ~n26798;
  assign n26801 = ~n26831 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n26800 = ~n26841 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n26802 = ~n26801 | ~n26800;
  assign n26804 = ~n26803 & ~n26802;
  assign n26826 = ~n26805 | ~n26804;
  assign n26810 = ~n26807 & ~n26806;
  assign n26809 = ~n26808 & ~n43425;
  assign n26812 = ~n26810 & ~n26809;
  assign n26811 = ~n26828 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n26816 = ~n26812 | ~n26811;
  assign n26814 = ~n26858 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n26813 = ~n26838 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n26815 = ~n26814 | ~n26813;
  assign n26824 = ~n26816 & ~n26815;
  assign n26822 = ~n26818 & ~n26817;
  assign n26821 = ~n26820 & ~n26819;
  assign n26823 = ~n26822 & ~n26821;
  assign n26825 = ~n26824 | ~n26823;
  assign n26830 = ~n26827 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n26829 = ~n26828 | ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n26836 = ~n26830 | ~n26829;
  assign n26834 = ~n26831 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n26833 = ~n26832 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n26835 = ~n26834 | ~n26833;
  assign n26847 = ~n26836 & ~n26835;
  assign n26840 = ~n26837 | ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n26839 = ~n26838 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n26845 = ~n26840 | ~n26839;
  assign n26843 = ~n22906 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n26842 = ~n26841 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n26844 = ~n26843 | ~n26842;
  assign n26846 = ~n26845 & ~n26844;
  assign n26870 = ~n26847 | ~n26846;
  assign n26851 = ~n26848 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n26850 = ~n26849 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n26857 = ~n26851 | ~n26850;
  assign n26855 = ~n26852 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n26854 = ~n22926 | ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n26856 = ~n26855 | ~n26854;
  assign n26868 = ~n26857 & ~n26856;
  assign n26861 = ~n26858 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n26860 = ~n26859 | ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n26866 = ~n26861 | ~n26860;
  assign n26864 = ~n26862 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n26863 = ~n23481 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n26865 = ~n26864 | ~n26863;
  assign n26867 = ~n26866 & ~n26865;
  assign n26869 = ~n26868 | ~n26867;
  assign n43500 = ~n43408;
  assign n26872 = ~n43500 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n26871 = ~n43503 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n26876 = ~n26872 | ~n26871;
  assign n26874 = ~n22911 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n43483 = ~n22927;
  assign n26873 = ~n43483 | ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n26875 = ~n26874 | ~n26873;
  assign n26885 = ~n26876 & ~n26875;
  assign n43495 = ~n26877;
  assign n26880 = ~n43495 | ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n26879 = ~n35715 | ~n35718;
  assign n43490 = ~n26879 | ~n26878;
  assign n43509 = ~n43490;
  assign n26883 = ~n26880 | ~n43509;
  assign n26881 = ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n26882 = ~n43094 & ~n26881;
  assign n26884 = ~n26883 & ~n26882;
  assign n26889 = ~n26885 | ~n26884;
  assign n26887 = ~n43484 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n26886 = ~n43499 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n26888 = ~n26887 | ~n26886;
  assign n26907 = n26889 | n26888;
  assign n26890 = ~n43499 | ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n26893 = ~n26890 | ~n43490;
  assign n26892 = ~n43408 & ~n26891;
  assign n26897 = n26893 | n26892;
  assign n26895 = ~n43484 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n26894 = ~n43503 | ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n26896 = ~n26895 | ~n26894;
  assign n26905 = ~n26897 & ~n26896;
  assign n26899 = ~n22911 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n26898 = ~n43483 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n26903 = ~n26899 | ~n26898;
  assign n26901 = ~n43495 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n26900 = ~n43496 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n26902 = ~n26901 | ~n26900;
  assign n26904 = ~n26903 & ~n26902;
  assign n26906 = ~n26905 | ~n26904;
  assign n41569 = ~n41790 & ~n43061;
  assign n41568 = ~n26908 | ~n26909;
  assign n42697 = ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n26918 = ~n26914 & ~n42697;
  assign n26915 = ~P2_EAX_REG_20__SCAN_IN;
  assign n26917 = ~n26916 & ~n26915;
  assign n26920 = ~n26918 & ~n26917;
  assign n37269 = ~n37271 | ~n37270;
  assign n29511 = ~P2_REIP_REG_21__SCAN_IN;
  assign n26922 = ~n41474 | ~P2_EAX_REG_21__SCAN_IN;
  assign n26921 = ~n28191 | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n39701 = ~n37269 & ~n37464;
  assign n26928 = ~n41473 | ~P2_REIP_REG_22__SCAN_IN;
  assign n26926 = ~n41474 | ~P2_EAX_REG_22__SCAN_IN;
  assign n26925 = ~n28191 | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n26927 = n26926 & n26925;
  assign n26932 = ~n41473 | ~P2_REIP_REG_23__SCAN_IN;
  assign n26930 = ~n41474 | ~P2_EAX_REG_23__SCAN_IN;
  assign n26929 = ~n28191 | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n26931 = n26930 & n26929;
  assign n26934 = ~BUF2_REG_7__SCAN_IN | ~n36558;
  assign n26933 = ~n36557 | ~BUF1_REG_7__SCAN_IN;
  assign n36590 = ~n26934 | ~n26933;
  assign n32348 = ~n36590;
  assign n26936 = ~n43697 & ~n32348;
  assign n31228 = ~P2_EAX_REG_23__SCAN_IN;
  assign n26935 = ~n41759 & ~n31228;
  assign n26937 = ~n26936 & ~n26935;
  assign n26941 = n26940 | n26939;
  assign P2_U2896 = n26942 | n26941;
  assign n26943 = ~P1_PHYADDRPOINTER_REG_20__SCAN_IN | ~n43722;
  assign n26946 = ~n43261 | ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n26945 = ~n43264 | ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n26950 = ~n26946 | ~n26945;
  assign n26948 = ~n43245 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n26947 = ~n43260 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n26949 = ~n26948 | ~n26947;
  assign n26958 = ~n26950 & ~n26949;
  assign n26952 = ~n43270 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n26951 = ~n43271 | ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n26956 = ~n26952 | ~n26951;
  assign n26954 = ~n43274 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n26953 = ~n22908 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n26955 = ~n26954 | ~n26953;
  assign n26957 = ~n26956 & ~n26955;
  assign n26974 = ~n26958 | ~n26957;
  assign n26960 = ~n22907 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n26959 = ~n43241 | ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n26964 = ~n26960 | ~n26959;
  assign n26962 = ~n43275 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n26961 = ~n43242 | ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n26963 = ~n26962 | ~n26961;
  assign n26972 = ~n26964 & ~n26963;
  assign n26966 = ~n43246 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n26965 = ~n43251 | ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n26970 = ~n26966 | ~n26965;
  assign n26968 = ~n43265 | ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n26967 = ~n22915 | ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n26969 = ~n26968 | ~n26967;
  assign n26971 = ~n26970 & ~n26969;
  assign n26973 = ~n26972 | ~n26971;
  assign n26975 = ~n26974 & ~n26973;
  assign n26976 = n26975 | n43286;
  assign n28484 = ~n26981 & ~n26980;
  assign n26984 = ~n22915 | ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n26983 = ~n43271 | ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n26988 = ~n26984 | ~n26983;
  assign n26986 = ~n43274 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n26985 = ~n43261 | ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n26987 = ~n26986 | ~n26985;
  assign n27019 = ~n26988 & ~n26987;
  assign n26990 = ~n43246 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n26989 = ~n43251 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n26994 = ~n26990 | ~n26989;
  assign n26992 = ~n22907 | ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n26991 = ~n43275 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n26993 = ~n26992 | ~n26991;
  assign n27002 = ~n26994 & ~n26993;
  assign n26996 = ~n43241 | ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n26995 = ~n43242 | ~P1_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n27000 = ~n26996 | ~n26995;
  assign n26998 = ~n43270 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n26997 = ~n43264 | ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n26999 = ~n26998 | ~n26997;
  assign n27001 = ~n27000 & ~n26999;
  assign n27017 = ~n27002 | ~n27001;
  assign n27008 = ~n27004 & ~n27003;
  assign n27005 = ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n27007 = ~n27006 & ~n27005;
  assign n27015 = ~n27008 & ~n27007;
  assign n27013 = ~n27009 & ~n23758;
  assign n27012 = ~n27011 & ~n27010;
  assign n27014 = ~n27013 & ~n27012;
  assign n27016 = ~n27015 | ~n27014;
  assign n27018 = ~n27017 & ~n27016;
  assign n27020 = ~n27019 | ~n27018;
  assign n27025 = ~n27020 | ~n28604;
  assign n31995 = ~P1_EAX_REG_21__SCAN_IN;
  assign n27023 = ~n28810 & ~n31995;
  assign n27021 = ~P1_PHYADDRPOINTER_REG_21__SCAN_IN & ~n39944;
  assign n27022 = ~P1_STATE2_REG_2__SCAN_IN & ~n27021;
  assign n27024 = ~n27023 & ~n27022;
  assign n27031 = ~n28512;
  assign n27039 = ~n42680 | ~n44021;
  assign n27038 = ~n44023 | ~P1_EBX_REG_21__SCAN_IN;
  assign P1_U2851 = n27041 | n27040;
  assign n40481 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n38144 = ~n40431 & ~n40481;
  assign n39786 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN | ~n38144;
  assign n27711 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN | ~P3_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n36049 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n36040 = ~n36049 & ~n41330;
  assign n27288 = ~n36040 | ~n33933;
  assign n27068 = ~n35663 & ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n36047 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n27230 = ~n27068 | ~n36047;
  assign n27069 = ~n33933 & ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n34042 = ~n27069 | ~n36048;
  assign n29442 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n36041 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n34773 = ~n27069 | ~n27068;
  assign n32515 = ~n27079 & ~n27078;
  assign n27114 = ~n36307 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n27113 = ~n36311 | ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n27121 = ~n22902 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n27135 = ~n36317 | ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n32808 = ~n27180 | ~n27179;
  assign n32208 = ~n27213 & ~n27212;
  assign n27252 = ~n36307 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n27254 = n27252 & n27251;
  assign n27316 = ~n35976;
  assign n27284 = ~n35392 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n27283 = ~n36307 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n27286 = n27284 & n27283;
  assign n27285 = ~n22903 | ~P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n27290 = ~n27286 | ~n27285;
  assign n27287 = ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n27289 = ~n27288 & ~n27287;
  assign n27298 = ~n27290 & ~n27289;
  assign n27292 = ~n36298 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n27291 = ~n22917 | ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n27296 = ~n27292 | ~n27291;
  assign n27294 = ~n36317 | ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n27293 = ~n22914 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n27295 = ~n27294 | ~n27293;
  assign n27297 = ~n27296 & ~n27295;
  assign n27300 = ~n22919 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n27299 = ~n22902 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n27305 = ~n27300 | ~n27299;
  assign n27303 = ~n22923 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n27302 = ~n36311 | ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n27304 = ~n27303 | ~n27302;
  assign n27313 = ~n27305 & ~n27304;
  assign n27307 = ~n36310 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n27306 = ~n22913 | ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n27311 = ~n27307 | ~n27306;
  assign n27309 = ~n36320 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n27308 = ~n22920 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n27310 = ~n27309 | ~n27308;
  assign n27312 = ~n27311 & ~n27310;
  assign n36526 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n36666 = n27324 | n27326;
  assign n36969 = n27331 | n27329;
  assign n27334 = n32501 | n27332;
  assign n36190 = ~n27710;
  assign n36230 = ~n40371 & ~n27748;
  assign n39395 = ~n37023 & ~n39388;
  assign n40244 = ~n40998 & ~n39785;
  assign n41541 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN | ~n27349;
  assign n28757 = ~n28755;
  assign n33487 = ~n27380 & ~n27379;
  assign n27403 = ~n36311 | ~P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n33501 = ~n27410 & ~n27409;
  assign n32672 = ~n27440 & ~n27439;
  assign n27442 = ~n22919 | ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n27441 = ~n36311 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n27448 = ~n22903 | ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n27450 = ~n36310 | ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n27455 = ~n22902 | ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n27461 = ~n36320 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n31802 = ~n27470 & ~n27469;
  assign n30706 = ~n27500 & ~n27499;
  assign n32475 = ~n27530 & ~n27529;
  assign n29940 = ~n27560 & ~n27559;
  assign n27581 = ~n36311 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n31801 = ~n27590 & ~n27589;
  assign n41542 = ~n32868 & ~n27593;
  assign n40422 = ~n31511 & ~n31807;
  assign n40141 = ~n27748;
  assign n27598 = ~n36352 & ~n40418;
  assign n36519 = ~n27598 & ~P3_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n40170 = ~n36519;
  assign n40166 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN | ~P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n40271 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN | ~P3_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n39622 = ~n40166 & ~n40271;
  assign n39624 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN | ~n39622;
  assign n40382 = ~n39620 & ~n39624;
  assign n40443 = n40170 & n40382;
  assign n39386 = ~n40141 | ~n40443;
  assign n39451 = ~n39386 & ~n39449;
  assign n40824 = ~n39772 & ~n40998;
  assign n40251 = ~n39451 | ~n40824;
  assign n27641 = ~n40251 & ~n41230;
  assign n41536 = ~n27641;
  assign n27624 = ~n40442 & ~n41536;
  assign n27793 = n27616 | n32475;
  assign n27621 = ~n38144;
  assign n40389 = ~n40382 | ~n40168;
  assign n39405 = ~n27748 & ~n40389;
  assign n39398 = ~n39405;
  assign n40471 = ~n39449 & ~n39398;
  assign n40417 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN | ~n40471;
  assign n39780 = ~n27621 & ~n40417;
  assign n40521 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~n39780;
  assign n39776 = ~n40531 & ~n40521;
  assign n27622 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~n39776;
  assign n41538 = ~n40998 & ~n27622;
  assign n27645 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~n41538;
  assign n27623 = ~n41537 & ~n27645;
  assign n27633 = ~n27624 & ~n27623;
  assign n40243 = ~n27625 & ~n27728;
  assign n40830 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~n40243;
  assign n41539 = ~n41230 & ~n40830;
  assign n32361 = ~n27630 | ~n27629;
  assign n27631 = n31805 | n42320;
  assign n27635 = ~n28093 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n27634 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n27636 = ~n41513 | ~n41005;
  assign n27652 = n27636 & P3_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n27651 = ~n42322 & ~P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n27639 = ~n41537 & ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n27637 = ~n40422 | ~n41516;
  assign n27638 = ~n28747 | ~n27637;
  assign n27649 = ~n27639 & ~n27638;
  assign n27640 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN | ~n41539;
  assign n27643 = ~n27640 | ~n40968;
  assign n27642 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN | ~n27641;
  assign n27648 = ~n27643 | ~n42323;
  assign n27644 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN | ~P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n27646 = ~n27645 & ~n27644;
  assign n27647 = ~n41537 & ~n27646;
  assign n27650 = ~n27649 | ~n28746;
  assign n27657 = ~n32284 & ~n27656;
  assign n27683 = ~n32501 | ~n27655;
  assign n27662 = ~n27658 | ~n27666;
  assign n35975 = ~n27659 & ~n40418;
  assign n36665 = ~n27665 | ~n27664;
  assign n36974 = ~n27670 | ~n27669;
  assign n27686 = ~n27682 | ~n27681;
  assign n27688 = ~n35988 | ~P3_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n36427 = ~n36429 & ~P3_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n27692 = ~n36427 & ~n41149;
  assign n27691 = ~n27690 & ~n39620;
  assign n27693 = ~n40127;
  assign n27694 = ~n27693 & ~n40403;
  assign n35859 = ~n40981 | ~n27696;
  assign n27698 = ~n27697 | ~n40403;
  assign n27699 = ~n35859 & ~n27698;
  assign n27701 = ~n27705 & ~n27700;
  assign n37107 = ~n27702 & ~n27701;
  assign n37106 = ~n37107 & ~P3_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n36192 = ~n37106 | ~n41147;
  assign n40132 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n27703 = ~n40132 & ~n27710;
  assign n36211 = ~n27707 | ~n27706;
  assign n27708 = ~n36211 & ~P3_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n27714 = ~n27708 & ~n41149;
  assign n27712 = ~n27711 & ~n27710;
  assign n37710 = ~n27714 & ~n27713;
  assign n27716 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n36885 = ~n27719 | ~n27718;
  assign n37569 = ~n36885 | ~n39440;
  assign n38147 = ~n37569 | ~n27722;
  assign n27723 = ~n40421 | ~n40431;
  assign n27725 = ~n27723 & ~P3_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n27724 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN & ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n27726 = ~n27725 | ~n27724;
  assign n27730 = ~n38147 | ~n27727;
  assign n37766 = ~n27730 | ~n27729;
  assign n39422 = ~n27732 | ~n27731;
  assign n27735 = ~n39422 | ~n27733;
  assign n27736 = ~n27735 | ~n27734;
  assign n38903 = ~n27736 & ~n42321;
  assign n27739 = ~n38903 & ~n41147;
  assign n38904 = ~n27736 | ~n42321;
  assign n40750 = ~n38904 | ~n41147;
  assign n27740 = ~n40750 | ~n41233;
  assign n41146 = ~n27737 | ~n27740;
  assign n28759 = ~n41146 & ~n41147;
  assign n27738 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN | ~P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n28099 = ~n41238 & ~n27738;
  assign n41252 = ~n27741 | ~n42337;
  assign n28760 = ~n27743 | ~n27742;
  assign n28098 = ~n28760 & ~P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n40202 = ~n32848 | ~n27747;
  assign n40451 = ~n36429 | ~n36075;
  assign n36227 = ~n40451 & ~n27748;
  assign n27806 = ~n27781 & ~n27775;
  assign n27779 = ~n27776;
  assign n27778 = ~n27790 & ~n27777;
  assign n27780 = ~n27779 & ~n27778;
  assign n31671 = ~n27806 & ~n27805;
  assign n29149 = ~P3_STATE_REG_0__SCAN_IN;
  assign n29561 = ~P3_STATE_REG_2__SCAN_IN | ~n29149;
  assign n27782 = P3_STATE_REG_1__SCAN_IN | n29561;
  assign n27783 = ~n31825 | ~n33487;
  assign n27794 = ~n27792;
  assign n27807 = n27805 & n27804;
  assign n27808 = ~n30706 & ~n31788;
  assign n41384 = ~P3_STATE2_REG_0__SCAN_IN | ~n35452;
  assign n42025 = ~n40527 & ~n41384;
  assign n41257 = n27817 & n42025;
  assign n40865 = n32966 | P3_STATE2_REG_0__SCAN_IN;
  assign n27819 = ~n40529 | ~P3_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n41410 = ~n41145 | ~P3_REIP_REG_31__SCAN_IN;
  assign P3_U2831 = n27821 | n27820;
  assign n27826 = ~n27824 | ~n27823;
  assign n41272 = ~P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n41185 = ~n43462 & ~n41272;
  assign n28477 = ~n41186 & ~n41185;
  assign n27827 = ~n43462 ^ P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n27832 = ~n41454 | ~n43367;
  assign n27830 = n43362 & n41444;
  assign n41744 = ~n43469 | ~P1_REIP_REG_18__SCAN_IN;
  assign n27828 = ~n43709 | ~P1_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n27829 = ~n41744 | ~n27828;
  assign n27831 = ~n27830 & ~n27829;
  assign P1_U2981 = n27834 | n27833;
  assign n29646 = ~P1_REIP_REG_19__SCAN_IN;
  assign n27835 = ~P1_REIP_REG_18__SCAN_IN | ~P1_REIP_REG_17__SCAN_IN;
  assign n27840 = ~n27836 & ~n27835;
  assign n27837 = ~n29646 & ~n41451;
  assign n27839 = ~n43469 & ~n27837;
  assign n27838 = ~n43797 | ~P1_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n41893 = ~n42405 | ~n41848;
  assign n27849 = ~n41893 & ~n27841;
  assign n27842 = ~n43796 | ~P1_EBX_REG_19__SCAN_IN;
  assign n27850 = n27849 | n27848;
  assign P1_U2821 = n27851 | n27850;
  assign n40759 = ~n27857 | ~n27856;
  assign n27864 = ~n40759 | ~n27861;
  assign n31714 = ~n35744 | ~n35805;
  assign n27874 = ~n42058 | ~n43809;
  assign n40760 = ~n27875;
  assign n27877 = ~n23322 | ~P2_EBX_REG_7__SCAN_IN;
  assign n42238 = n40760 & n41078;
  assign n42086 = ~n42242 | ~n42238;
  assign n27881 = ~n23322 | ~P2_EBX_REG_8__SCAN_IN;
  assign n27884 = ~n41491 | ~n41072;
  assign n27883 = ~n37329;
  assign n27886 = ~n41072 | ~n41697;
  assign n28198 = ~n23322 | ~P2_EBX_REG_10__SCAN_IN;
  assign n27890 = ~n42081 ^ P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n43913 = ~n31714 & ~n43061;
  assign n27933 = ~n28076 | ~n43913;
  assign n28158 = ~n31495 | ~n32176;
  assign n27892 = ~n28150 | ~n27891;
  assign n29199 = ~P2_REIP_REG_7__SCAN_IN;
  assign n27896 = ~n39573 | ~P2_EBX_REG_7__SCAN_IN;
  assign n27895 = ~P2_PHYADDRPOINTER_REG_7__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n27903 = ~n39573 | ~P2_EBX_REG_8__SCAN_IN;
  assign n27902 = ~P2_PHYADDRPOINTER_REG_8__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n27906 = ~n27912 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n27909 = ~n39573 | ~P2_EBX_REG_9__SCAN_IN;
  assign n27908 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n27913 = ~n27912 | ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n27917 = ~n39573 | ~P2_EBX_REG_10__SCAN_IN;
  assign n27916 = ~P2_PHYADDRPOINTER_REG_10__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n40299 = ~n28228 ^ n28226;
  assign n34920 = ~n40299;
  assign n27926 = ~n43915 & ~n34920;
  assign n32180 = ~n39508 & ~n36365;
  assign n27922 = ~n32180 & ~P2_STATE2_REG_0__SCAN_IN;
  assign n43917 = ~n27923 & ~n27922;
  assign n27924 = ~n43917 | ~P2_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n28077 = ~n43880 | ~P2_REIP_REG_10__SCAN_IN;
  assign n27925 = ~n27924 | ~n28077;
  assign n27931 = n27926 | n27925;
  assign n28159 = ~P2_STATE2_REG_1__SCAN_IN | ~n38321;
  assign n33577 = ~n27927 | ~n28159;
  assign n27928 = ~n33577;
  assign n43896 = ~n43917 & ~n27928;
  assign n40285 = ~P2_PHYADDRPOINTER_REG_10__SCAN_IN ^ n27929;
  assign n27930 = ~n43911 & ~n40285;
  assign n27932 = ~n27931 & ~n27930;
  assign P2_U3004 = n27935 | n27934;
  assign n27937 = ~n43721 | ~P1_EAX_REG_22__SCAN_IN;
  assign n27936 = ~P1_PHYADDRPOINTER_REG_22__SCAN_IN | ~n43722;
  assign n27939 = ~n43264 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n27938 = ~n43265 | ~P1_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n27943 = ~n27939 | ~n27938;
  assign n27941 = ~n22908 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n27940 = ~n43260 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n27942 = ~n27941 | ~n27940;
  assign n27951 = ~n27943 & ~n27942;
  assign n27945 = ~n43245 | ~P1_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n27944 = ~n43275 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n27949 = ~n27945 | ~n27944;
  assign n27947 = ~n43270 | ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n27946 = ~n43274 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n27948 = ~n27947 | ~n27946;
  assign n27950 = ~n27949 & ~n27948;
  assign n27967 = ~n27951 | ~n27950;
  assign n27953 = ~n22907 | ~P1_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n27952 = ~n28775 | ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n27957 = ~n27953 | ~n27952;
  assign n27955 = ~n43251 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n27954 = ~n43261 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n27956 = ~n27955 | ~n27954;
  assign n27965 = ~n27957 & ~n27956;
  assign n27959 = ~n43246 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n27958 = ~n43242 | ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n27963 = ~n27959 | ~n27958;
  assign n27961 = ~n22915 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n27960 = ~n43271 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n27962 = ~n27961 | ~n27960;
  assign n27964 = ~n27963 & ~n27962;
  assign n27966 = ~n27965 | ~n27964;
  assign n27968 = ~n27967 & ~n27966;
  assign n27969 = n27968 | n43286;
  assign n27970 = ~n27969 | ~n43725;
  assign n27976 = ~n22907 | ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n27975 = ~n43251 | ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n27980 = ~n27976 | ~n27975;
  assign n27978 = ~n43246 | ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n27977 = ~n22908 | ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n27979 = ~n27978 | ~n27977;
  assign n27988 = ~n27980 & ~n27979;
  assign n27982 = ~n28775 | ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n27981 = ~n43242 | ~P1_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n27986 = ~n27982 | ~n27981;
  assign n27984 = ~n43270 | ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n27983 = ~n43264 | ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n27985 = ~n27984 | ~n27983;
  assign n27987 = ~n27986 & ~n27985;
  assign n28004 = ~n27988 | ~n27987;
  assign n27990 = ~n43274 | ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n27989 = ~n43265 | ~P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n27994 = ~n27990 | ~n27989;
  assign n27992 = ~n43261 | ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n27991 = ~n22915 | ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n27993 = ~n27992 | ~n27991;
  assign n28002 = ~n27994 & ~n27993;
  assign n27996 = ~n43275 | ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n27995 = ~n43271 | ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n28000 = ~n27996 | ~n27995;
  assign n27998 = ~n43245 | ~P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n27997 = ~n43260 | ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n27999 = ~n27998 | ~n27997;
  assign n28001 = ~n28000 & ~n27999;
  assign n28003 = ~n28002 | ~n28001;
  assign n28378 = ~n28004 & ~n28003;
  assign n28006 = ~n22907 | ~P1_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n28005 = ~n28775 | ~P1_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n28010 = ~n28006 | ~n28005;
  assign n28008 = ~n22908 | ~P1_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n28007 = ~n43242 | ~P1_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n28009 = ~n28008 | ~n28007;
  assign n28018 = ~n28010 & ~n28009;
  assign n28012 = ~n43246 | ~P1_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n28011 = ~n43251 | ~P1_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n28016 = ~n28012 | ~n28011;
  assign n28014 = ~n43265 | ~P1_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n28013 = ~n43271 | ~P1_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n28015 = ~n28014 | ~n28013;
  assign n28017 = ~n28016 & ~n28015;
  assign n28034 = ~n28018 | ~n28017;
  assign n28020 = ~n43245 | ~P1_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n28019 = ~n43260 | ~P1_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n28024 = ~n28020 | ~n28019;
  assign n28022 = ~n43270 | ~P1_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n28021 = ~n43274 | ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n28023 = ~n28022 | ~n28021;
  assign n28032 = ~n28024 & ~n28023;
  assign n28026 = ~n43264 | ~P1_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n28025 = ~n22915 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n28030 = ~n28026 | ~n28025;
  assign n28028 = ~n43275 | ~P1_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n28027 = ~n43261 | ~P1_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n28029 = ~n28028 | ~n28027;
  assign n28031 = ~n28030 & ~n28029;
  assign n28033 = ~n28032 | ~n28031;
  assign n28377 = ~n28034 & ~n28033;
  assign n28035 = ~n28378 ^ n28377;
  assign n28042 = n28035 | n43286;
  assign n32001 = ~P1_EAX_REG_23__SCAN_IN;
  assign n28040 = ~n28810 & ~n32001;
  assign n28038 = ~n28608 | ~P1_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n28551 = ~n41435 & ~n28047;
  assign n28055 = ~n28551 | ~n28550;
  assign n28058 = ~n42408 | ~n44021;
  assign n28057 = ~n44023 | ~P1_EBX_REG_23__SCAN_IN;
  assign P1_U2849 = n28060 | n28059;
  assign n28063 = ~n41697 & ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n28064 = ~n28062 & ~n28061;
  assign n28073 = ~n28063 | ~n42558;
  assign n28066 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN | ~n28064;
  assign n42105 = ~n28066 & ~n28065;
  assign n28069 = ~n43159 & ~n42105;
  assign n42109 = ~n28067 & ~n28066;
  assign n28068 = ~n42699 & ~n42109;
  assign n28070 = ~n28069 & ~n28068;
  assign n41698 = n28070 & n42110;
  assign n42557 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN | ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n28071 = ~n42557 | ~n43165;
  assign n28072 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN | ~n42560;
  assign n28087 = ~n28073 | ~n28072;
  assign n28083 = ~n28076 | ~n43876;
  assign n28078 = ~n43767 | ~n40299;
  assign n28081 = ~n28078 | ~n28077;
  assign n28080 = ~n43877 & ~n40298;
  assign n28082 = ~n28081 & ~n28080;
  assign n28086 = n28085 | n28084;
  assign P2_U3036 = n28087 | n28086;
  assign n28089 = ~n28088 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n28094 = n28093 | P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n28104 = ~n40529 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n41527 = ~n41145 | ~P3_REIP_REG_30__SCAN_IN;
  assign P3_U2832 = n28106 | n28105;
  assign n43774 = P2_PHYADDRPOINTER_REG_28__SCAN_IN ^ n28107;
  assign n43326 = P2_PHYADDRPOINTER_REG_26__SCAN_IN ^ n28108;
  assign n43217 = P2_PHYADDRPOINTER_REG_24__SCAN_IN ^ n28109;
  assign n43000 = P2_PHYADDRPOINTER_REG_22__SCAN_IN ^ n28110;
  assign n42473 = P2_PHYADDRPOINTER_REG_20__SCAN_IN ^ n28111;
  assign n42438 = P2_PHYADDRPOINTER_REG_18__SCAN_IN ^ n28112;
  assign n42393 = ~P2_PHYADDRPOINTER_REG_16__SCAN_IN ^ n28113;
  assign n40626 = ~n42393;
  assign n42847 = ~P2_PHYADDRPOINTER_REG_14__SCAN_IN ^ n28114;
  assign n42457 = ~P2_PHYADDRPOINTER_REG_12__SCAN_IN ^ n28115;
  assign n40648 = ~n42457;
  assign n40294 = ~n40285;
  assign n41176 = P2_PHYADDRPOINTER_REG_8__SCAN_IN ^ n28116;
  assign n40157 = P2_PHYADDRPOINTER_REG_6__SCAN_IN ^ n28117;
  assign n40574 = P2_PHYADDRPOINTER_REG_4__SCAN_IN ^ n28118;
  assign n40320 = P2_PHYADDRPOINTER_REG_2__SCAN_IN ^ P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n28121 = ~n28119 & ~n36357;
  assign n28120 = ~P2_STATE2_REG_0__SCAN_IN & ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n36501 = ~n28121 & ~n28120;
  assign n40319 = ~n37285 | ~n36501;
  assign n38828 = ~n40320 & ~n40319;
  assign n38829 = ~n28123 ^ n28122;
  assign n40573 = ~n38828 | ~n38829;
  assign n40362 = ~n40574 & ~n40573;
  assign n40363 = ~n28125 ^ n28124;
  assign n39722 = ~n40362 | ~n40363;
  assign n39721 = ~n40157 & ~n39722;
  assign n40948 = ~n28127 ^ n28126;
  assign n38941 = ~n39721 | ~n40948;
  assign n39471 = ~n41176 & ~n38941;
  assign n41504 = ~n28129 ^ n28128;
  assign n40293 = ~n39471 | ~n41504;
  assign n40296 = ~n40294 & ~n40293;
  assign n42061 = ~n42070 ^ n28130;
  assign n40647 = ~n40296 | ~n42061;
  assign n40646 = ~n40648 & ~n40647;
  assign n42145 = ~n28132 ^ n28131;
  assign n40671 = ~n40646 | ~n42145;
  assign n40670 = ~n40672 & ~n40671;
  assign n42429 = ~n28134 ^ n28133;
  assign n40625 = ~n40670 | ~n42429;
  assign n40624 = ~n40626 & ~n40625;
  assign n42260 = ~n28136 ^ n28135;
  assign n39222 = ~n40624 | ~n42260;
  assign n37716 = ~n42438 & ~n39222;
  assign n42345 = ~n42354 ^ n28137;
  assign n37717 = ~n37716 | ~n42345;
  assign n37452 = ~n42473 & ~n37717;
  assign n42856 = ~n28139 ^ n28138;
  assign n39693 = ~n37452 | ~n42856;
  assign n40107 = ~n43000 & ~n39693;
  assign n42960 = ~n28141 ^ n28140;
  assign n39749 = ~n40107 | ~n42960;
  assign n39913 = ~n43217 & ~n39749;
  assign n43546 = ~n43539 ^ n28142;
  assign n40918 = ~n39913 | ~n43546;
  assign n41203 = ~n43326 & ~n40918;
  assign n43654 = ~n28144 ^ n28143;
  assign n41719 = ~n41203 | ~n43654;
  assign n41913 = ~n43774 & ~n41719;
  assign n43897 = P2_PHYADDRPOINTER_REG_30__SCAN_IN ^ n28147;
  assign n28161 = n28148 ^ n43897;
  assign n28154 = ~n36357 & ~P2_STATE2_REG_2__SCAN_IN;
  assign n28155 = ~n28154 | ~P2_STATE2_REG_3__SCAN_IN;
  assign n28157 = ~n44003 & ~n35804;
  assign n28160 = ~n28157 | ~n28156;
  assign n41919 = ~P2_STATE2_REG_1__SCAN_IN | ~n40350;
  assign n28374 = ~n28161 & ~n41919;
  assign n28164 = ~n28162;
  assign n39758 = ~n28164 | ~n28163;
  assign n28168 = ~n25550 & ~n28316;
  assign n28166 = ~n41474 | ~P2_EAX_REG_24__SCAN_IN;
  assign n28165 = ~n28191 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n28167 = ~n28166 | ~n28165;
  assign n39910 = ~n39758 & ~n39759;
  assign n28172 = ~n41473 | ~P2_REIP_REG_25__SCAN_IN;
  assign n28170 = ~n41474 | ~P2_EAX_REG_25__SCAN_IN;
  assign n28169 = ~n28191 | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n28171 = n28170 & n28169;
  assign n40923 = ~n39910 | ~n39909;
  assign n28177 = ~n40923;
  assign n28176 = ~n41473 | ~P2_REIP_REG_26__SCAN_IN;
  assign n28174 = ~n41474 | ~P2_EAX_REG_26__SCAN_IN;
  assign n28173 = ~n28191 | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n28175 = n28174 & n28173;
  assign n41209 = ~n28177 | ~n40921;
  assign n29525 = ~P2_REIP_REG_27__SCAN_IN;
  assign n28181 = ~n25550 & ~n29525;
  assign n28179 = ~n41474 | ~P2_EAX_REG_27__SCAN_IN;
  assign n28178 = ~n28191 | ~P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n28180 = ~n28179 | ~n28178;
  assign n41725 = ~n41209 & ~n41208;
  assign n28185 = ~n25550 & ~n28345;
  assign n28183 = ~n41474 | ~P2_EAX_REG_28__SCAN_IN;
  assign n28182 = ~n28191 | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n28184 = ~n28183 | ~n28182;
  assign n41724 = ~n28185 & ~n28184;
  assign n41928 = ~n41725 | ~n28186;
  assign n28190 = ~n25550 & ~n28354;
  assign n28188 = ~n41474 | ~P2_EAX_REG_29__SCAN_IN;
  assign n28187 = ~n28191 | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n28189 = ~n28188 | ~n28187;
  assign n41471 = ~n41928 & ~n41927;
  assign n29484 = ~P2_REIP_REG_30__SCAN_IN;
  assign n28195 = ~n25550 & ~n29484;
  assign n28193 = ~n41474 | ~P2_EAX_REG_30__SCAN_IN;
  assign n28192 = ~n28191 | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n28194 = ~n28193 | ~n28192;
  assign n43878 = n41471 ^ n41472;
  assign n37288 = ~n41920 & ~n39511;
  assign n40602 = ~n41879 & ~n41877;
  assign n40651 = ~n23322 | ~P2_EBX_REG_12__SCAN_IN;
  assign n40675 = ~n23322 | ~P2_EBX_REG_14__SCAN_IN;
  assign n40629 = ~n23322 | ~P2_EBX_REG_16__SCAN_IN;
  assign n39211 = ~n40630 | ~n40629;
  assign n36384 = ~n23322 | ~P2_EBX_REG_18__SCAN_IN;
  assign n37736 = ~n36385 | ~n36384;
  assign n28204 = ~P2_EBX_REG_19__SCAN_IN;
  assign n37273 = ~n23322 | ~P2_EBX_REG_20__SCAN_IN;
  assign n37469 = ~n37274 | ~n37273;
  assign n28205 = ~P2_EBX_REG_21__SCAN_IN;
  assign n39709 = ~n23322 | ~P2_EBX_REG_22__SCAN_IN;
  assign n40121 = ~n39710 | ~n39709;
  assign n40120 = ~n23322 | ~P2_EBX_REG_23__SCAN_IN;
  assign n39763 = ~n23322 | ~P2_EBX_REG_24__SCAN_IN;
  assign n39928 = ~n39764 | ~n39763;
  assign n28207 = ~P2_EBX_REG_25__SCAN_IN;
  assign n40926 = ~n39928 & ~n39927;
  assign n40925 = ~n23322 | ~P2_EBX_REG_26__SCAN_IN;
  assign n41874 = ~n40926 | ~n40925;
  assign n41213 = ~P2_EBX_REG_27__SCAN_IN;
  assign n41727 = ~n41874 & ~n41212;
  assign n41726 = ~n23322 | ~P2_EBX_REG_28__SCAN_IN;
  assign n28208 = ~P2_EBX_REG_29__SCAN_IN;
  assign n28209 = ~n23322 | ~P2_EBX_REG_30__SCAN_IN;
  assign n28369 = ~n36364 | ~n38321;
  assign n28214 = ~n23085 | ~n28369;
  assign n39482 = n28214 | n28210;
  assign n28212 = ~P2_EBX_REG_31__SCAN_IN;
  assign n28215 = n28214 | n28213;
  assign n28221 = ~n41935 | ~P2_EBX_REG_30__SCAN_IN;
  assign n28217 = ~P2_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n36390 = n41920 | n39522;
  assign n28219 = ~n28217 & ~n36390;
  assign n28218 = ~n29484 & ~n40350;
  assign n28220 = ~n28219 & ~n28218;
  assign n28224 = n28223 | n28222;
  assign n28231 = ~n39573 | ~P2_EBX_REG_11__SCAN_IN;
  assign n28230 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n28238 = ~n39573 | ~P2_EBX_REG_12__SCAN_IN;
  assign n28237 = ~P2_PHYADDRPOINTER_REG_12__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28244 = ~n39573 | ~P2_EBX_REG_13__SCAN_IN;
  assign n28243 = ~P2_PHYADDRPOINTER_REG_13__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28251 = ~n39573 | ~P2_EBX_REG_14__SCAN_IN;
  assign n28250 = ~P2_PHYADDRPOINTER_REG_14__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28256 = ~P2_PHYADDRPOINTER_REG_15__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28263 = ~P2_PHYADDRPOINTER_REG_16__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28270 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n36380 = ~P2_REIP_REG_18__SCAN_IN;
  assign n28276 = ~P2_PHYADDRPOINTER_REG_18__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28283 = ~P2_PHYADDRPOINTER_REG_19__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28290 = ~P2_PHYADDRPOINTER_REG_20__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28297 = ~n23598 | ~P2_EBX_REG_21__SCAN_IN;
  assign n28296 = ~P2_PHYADDRPOINTER_REG_21__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28306 = ~n28361 & ~n28302;
  assign n28304 = ~n23598 | ~P2_EBX_REG_22__SCAN_IN;
  assign n28303 = ~P2_PHYADDRPOINTER_REG_22__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n29520 = ~P2_REIP_REG_23__SCAN_IN;
  assign n28313 = ~n28361 & ~n29520;
  assign n28311 = ~n23598 | ~P2_EBX_REG_23__SCAN_IN;
  assign n28310 = ~P2_PHYADDRPOINTER_REG_23__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28312 = ~n28311 | ~n28310;
  assign n28320 = ~n28361 & ~n28316;
  assign n28318 = ~n23598 | ~P2_EBX_REG_24__SCAN_IN;
  assign n28317 = ~P2_PHYADDRPOINTER_REG_24__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28319 = ~n28318 | ~n28317;
  assign n28328 = ~n28361 & ~n28324;
  assign n28326 = ~n23598 | ~P2_EBX_REG_25__SCAN_IN;
  assign n28325 = ~P2_PHYADDRPOINTER_REG_25__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28327 = ~n28326 | ~n28325;
  assign n40936 = ~n39921 | ~n39920;
  assign n28335 = ~n28361 & ~n28331;
  assign n28333 = ~n23598 | ~P2_EBX_REG_26__SCAN_IN;
  assign n28332 = ~P2_PHYADDRPOINTER_REG_26__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28334 = ~n28333 | ~n28332;
  assign n28337 = ~n28335 & ~n28334;
  assign n28342 = ~n28361 & ~n29525;
  assign n28340 = ~n23598 | ~P2_EBX_REG_27__SCAN_IN;
  assign n28339 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n28341 = ~n28340 | ~n28339;
  assign n28344 = ~n28342 & ~n28341;
  assign n28343 = ~n39578 | ~P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n41733 = ~n41224 | ~n41223;
  assign n28350 = ~n28361 & ~n28345;
  assign n28348 = ~n23598 | ~P2_EBX_REG_28__SCAN_IN;
  assign n28347 = ~P2_PHYADDRPOINTER_REG_28__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28349 = ~n28348 | ~n28347;
  assign n28352 = ~n28350 & ~n28349;
  assign n28351 = ~n39578 | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n41941 = ~n41733 & ~n28353;
  assign n28358 = ~n28361 & ~n28354;
  assign n28356 = ~n23598 | ~P2_EBX_REG_29__SCAN_IN;
  assign n28355 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n28357 = ~n28356 | ~n28355;
  assign n28360 = ~n28358 & ~n28357;
  assign n28359 = ~n39578 | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n39571 = ~n41941 | ~n41940;
  assign n28365 = ~n28361 & ~n29484;
  assign n28363 = ~n23598 | ~P2_EBX_REG_30__SCAN_IN;
  assign n28362 = ~P2_PHYADDRPOINTER_REG_30__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28364 = ~n28363 | ~n28362;
  assign n28367 = ~n28365 & ~n28364;
  assign n28366 = ~n39578 | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign P2_U2825 = n28374 | n28373;
  assign n28376 = ~n43721 | ~P1_EAX_REG_24__SCAN_IN;
  assign n28375 = ~P1_PHYADDRPOINTER_REG_24__SCAN_IN | ~n43722;
  assign n28412 = ~n28376 | ~n28375;
  assign n28417 = ~n28378 & ~n28377;
  assign n28380 = ~n43251 | ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n28379 = ~n43242 | ~P1_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n28384 = ~n28380 | ~n28379;
  assign n28382 = ~n43241 | ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n28381 = ~n43270 | ~P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n28383 = ~n28382 | ~n28381;
  assign n28392 = ~n28384 & ~n28383;
  assign n28386 = ~n22907 | ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n28385 = ~n43246 | ~P1_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n28390 = ~n28386 | ~n28385;
  assign n28388 = ~n43274 | ~P1_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n28387 = ~n43275 | ~P1_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n28389 = ~n28388 | ~n28387;
  assign n28391 = ~n28390 & ~n28389;
  assign n28408 = ~n28392 | ~n28391;
  assign n28394 = ~n43260 | ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n28393 = ~n22915 | ~P1_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n28398 = ~n28394 | ~n28393;
  assign n28396 = ~n43245 | ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n28395 = ~n22908 | ~P1_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n28397 = ~n28396 | ~n28395;
  assign n28406 = ~n28398 & ~n28397;
  assign n28400 = ~n43261 | ~P1_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n28399 = ~n43265 | ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n28404 = ~n28400 | ~n28399;
  assign n28402 = ~n43264 | ~P1_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n28401 = ~n43271 | ~P1_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n28403 = ~n28402 | ~n28401;
  assign n28405 = ~n28404 & ~n28403;
  assign n28407 = ~n28406 | ~n28405;
  assign n28416 = n28408 | n28407;
  assign n28409 = ~n28417 ^ n28416;
  assign n28410 = n28409 | n43286;
  assign n28411 = ~n28410 | ~n43725;
  assign n28524 = ~n28415 & ~n28414;
  assign n28450 = ~n28417 | ~n28416;
  assign n28449 = ~n28450 | ~n28604;
  assign n28419 = ~n22907 | ~P1_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n28418 = ~n43242 | ~P1_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n28423 = ~n28419 | ~n28418;
  assign n28421 = ~n43246 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n28420 = ~n43260 | ~P1_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n28422 = ~n28421 | ~n28420;
  assign n28431 = ~n28423 & ~n28422;
  assign n28425 = ~n28775 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n28424 = ~n43251 | ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n28429 = ~n28425 | ~n28424;
  assign n28427 = ~n43261 | ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n28426 = ~n43265 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n28428 = ~n28427 | ~n28426;
  assign n28430 = ~n28429 & ~n28428;
  assign n28447 = ~n28431 | ~n28430;
  assign n28433 = ~n22915 | ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n28432 = ~n43271 | ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n28437 = ~n28433 | ~n28432;
  assign n28435 = ~n43270 | ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n28434 = ~n43274 | ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n28436 = ~n28435 | ~n28434;
  assign n28445 = ~n28437 & ~n28436;
  assign n28439 = ~n22908 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n28438 = ~n43264 | ~P1_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n28443 = ~n28439 | ~n28438;
  assign n28441 = ~n43245 | ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n28440 = ~n43275 | ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n28442 = ~n28441 | ~n28440;
  assign n28444 = ~n28443 & ~n28442;
  assign n28446 = ~n28445 | ~n28444;
  assign n28603 = ~n28447 & ~n28446;
  assign n28448 = ~n28603;
  assign n28452 = ~n28449 | ~n28448;
  assign n28602 = n28450 | n43286;
  assign n28451 = ~n28602 | ~n28603;
  assign n28458 = ~n28452 | ~n28451;
  assign n28453 = ~P1_EAX_REG_25__SCAN_IN;
  assign n28456 = ~n28810 & ~n28453;
  assign n28454 = ~P1_PHYADDRPOINTER_REG_25__SCAN_IN | ~n43722;
  assign n28455 = ~n43725 | ~n28454;
  assign n28457 = ~n28456 & ~n28455;
  assign n28462 = ~n28461 | ~n28460;
  assign n43031 = ~n28465 | ~n28464;
  assign n28467 = ~n40080 | ~P1_EBX_REG_24__SCAN_IN;
  assign n28662 = ~n28523 | ~n28522;
  assign n28470 = ~n40080 | ~P1_EBX_REG_25__SCAN_IN;
  assign n28472 = ~n44023 | ~P1_EBX_REG_25__SCAN_IN;
  assign P1_U2847 = n28475 | n28474;
  assign n42501 = ~n28477 | ~n28476;
  assign n28480 = ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n42587 = ~n43469 | ~P1_REIP_REG_20__SCAN_IN;
  assign n28486 = ~n43709 | ~P1_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n28488 = ~n42587 | ~n28486;
  assign n28487 = ~n43713 & ~n41899;
  assign n28489 = ~n28488 & ~n28487;
  assign P1_U2979 = n28492 | n28491;
  assign n41989 = ~P1_INSTADDRPOINTER_REG_19__SCAN_IN | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n42580 = ~n41989;
  assign n28493 = ~n42580 | ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n28506 = ~n41949 & ~n28493;
  assign n28496 = ~n28506 | ~P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n42579 = ~P1_INSTADDRPOINTER_REG_20__SCAN_IN & ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n28560 = ~P1_INSTADDRPOINTER_REG_22__SCAN_IN & ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n41999 = ~n42579 | ~n28560;
  assign n28495 = ~n28507 | ~n28494;
  assign n28852 = ~n28495 | ~n22933;
  assign n42372 = ~n43469 | ~P1_REIP_REG_23__SCAN_IN;
  assign n28498 = ~n43709 | ~P1_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n28500 = ~n42372 | ~n28498;
  assign n28499 = ~n43713 & ~n42410;
  assign n28501 = ~n28500 & ~n28499;
  assign P1_U2976 = n28504 | n28503;
  assign n28552 = ~n43469 | ~P1_REIP_REG_22__SCAN_IN;
  assign n28513 = ~n43709 | ~P1_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n28515 = ~n28552 | ~n28513;
  assign n28514 = ~n43713 & ~n42174;
  assign n28516 = ~n28515 & ~n28514;
  assign P1_U2977 = n28519 | n28518;
  assign n28521 = ~n43796 | ~P1_EBX_REG_24__SCAN_IN;
  assign n28520 = ~n43797 | ~P1_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n29684 = ~P1_REIP_REG_24__SCAN_IN;
  assign n42186 = ~P1_REIP_REG_22__SCAN_IN;
  assign n41896 = ~P1_REIP_REG_20__SCAN_IN;
  assign n28526 = ~n41896 & ~n41848;
  assign n42403 = ~n42186 & ~n42184;
  assign n42161 = ~n29684 & ~n42404;
  assign n28527 = ~n42404 | ~n29684;
  assign n28528 = ~n28527 | ~n42405;
  assign n28532 = n42161 | n28528;
  assign n28530 = ~n42175 & ~n28737;
  assign n28529 = ~n41894 & ~n29684;
  assign n28531 = ~n28530 & ~n28529;
  assign P1_U2816 = n28538 | n28537;
  assign n28540 = ~P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n40796 = ~n28540 & ~n28539;
  assign n28544 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN | ~n40796;
  assign n28558 = ~n28541 & ~n28544;
  assign n28542 = ~n41976 & ~n28558;
  assign n41962 = ~P1_INSTADDRPOINTER_REG_18__SCAN_IN | ~P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n41963 = ~n41962;
  assign n43335 = ~n42580 | ~n41963;
  assign n28543 = ~n36891 | ~n43335;
  assign n28546 = ~n28544;
  assign n42919 = ~n43330 & ~n43335;
  assign n28547 = ~n36895 & ~n42919;
  assign n28548 = ~n42676;
  assign n42364 = ~n28559 & ~n43333;
  assign n42826 = n42364 | n43335;
  assign n41990 = ~P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n42675 = ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n42365 = ~n41990 & ~n42675;
  assign n28561 = n28560 | n42365;
  assign n28562 = ~n42826 & ~n28561;
  assign P1_U3009 = n28563 | n28562;
  assign n28565 = ~n43245 | ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n28564 = ~n22908 | ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n28569 = ~n28565 | ~n28564;
  assign n28567 = ~n43270 | ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n28566 = ~n43264 | ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n28568 = ~n28567 | ~n28566;
  assign n28601 = ~n28569 & ~n28568;
  assign n28571 = ~n28775 | ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n28570 = ~n43242 | ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n28575 = ~n28571 | ~n28570;
  assign n28573 = ~n43246 | ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n28572 = ~n43265 | ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n28574 = ~n28573 | ~n28572;
  assign n28583 = ~n28575 & ~n28574;
  assign n28577 = ~n22907 | ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n28576 = ~n43251 | ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n28581 = ~n28577 | ~n28576;
  assign n28579 = ~n43260 | ~P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n28578 = ~n43261 | ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n28580 = ~n28579 | ~n28578;
  assign n28582 = ~n28581 & ~n28580;
  assign n28599 = ~n28583 | ~n28582;
  assign n28589 = ~n28585 & ~n28584;
  assign n28588 = ~n28587 & ~n28586;
  assign n28597 = ~n28589 & ~n28588;
  assign n28595 = ~n28591 & ~n28590;
  assign n28594 = ~n28593 & ~n28592;
  assign n28596 = ~n28595 & ~n28594;
  assign n28598 = ~n28597 | ~n28596;
  assign n28600 = ~n28599 & ~n28598;
  assign n28605 = n28616 ^ n28615;
  assign n28607 = ~n28605 | ~n28604;
  assign n28606 = ~n43721 | ~P1_EAX_REG_26__SCAN_IN;
  assign n28611 = ~n28607 | ~n28606;
  assign n28609 = ~n28608 | ~P1_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n28610 = ~n28609 | ~n43725;
  assign n28614 = ~n28611 & ~n28610;
  assign n28658 = ~n28835 | ~n28834;
  assign n28618 = ~n43251 | ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n28617 = ~n43242 | ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n28622 = ~n28618 | ~n28617;
  assign n28620 = ~n43241 | ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n28619 = ~n43271 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n28621 = ~n28620 | ~n28619;
  assign n28630 = ~n28622 & ~n28621;
  assign n28624 = ~n22907 | ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n28623 = ~n43246 | ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n28628 = ~n28624 | ~n28623;
  assign n28626 = ~n22908 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n28625 = ~n43260 | ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n28627 = ~n28626 | ~n28625;
  assign n28629 = ~n28628 & ~n28627;
  assign n28646 = ~n28630 | ~n28629;
  assign n28632 = ~n43245 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n28631 = ~n22915 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n28636 = ~n28632 | ~n28631;
  assign n28634 = ~n43270 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n28633 = ~n43275 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n28635 = ~n28634 | ~n28633;
  assign n28644 = ~n28636 & ~n28635;
  assign n28638 = ~n43261 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n28637 = ~n43264 | ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n28642 = ~n28638 | ~n28637;
  assign n28640 = ~n43274 | ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n28639 = ~n43265 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n28641 = ~n28640 | ~n28639;
  assign n28643 = ~n28642 & ~n28641;
  assign n28645 = ~n28644 | ~n28643;
  assign n28707 = ~n28646 & ~n28645;
  assign n28647 = n28706 ^ n28707;
  assign n28653 = ~n28647 | ~n28604;
  assign n28651 = ~n28810 & ~n28648;
  assign n28649 = ~P1_PHYADDRPOINTER_REG_27__SCAN_IN | ~n43722;
  assign n28650 = ~n43725 | ~n28649;
  assign n28652 = ~n28651 & ~n28650;
  assign n28774 = ~n28658 & ~n28657;
  assign n28659 = ~n28658 | ~n28657;
  assign n43377 = ~n28660 | ~n28659;
  assign n28833 = ~n28662 & ~n28661;
  assign n28664 = ~n40080 | ~P1_EBX_REG_26__SCAN_IN;
  assign n28670 = ~n28833 | ~n28832;
  assign n28667 = ~n40080 | ~P1_EBX_REG_27__SCAN_IN;
  assign n28666 = ~n40081 | ~P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n28721 = ~n28670 & ~n28669;
  assign P1_U2845 = n28675 | n28674;
  assign n28677 = ~n43274 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n28676 = ~n22915 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n28681 = ~n28677 | ~n28676;
  assign n28679 = ~n43270 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n28678 = ~n43260 | ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n28680 = ~n28679 | ~n28678;
  assign n28685 = n28681 | n28680;
  assign n28683 = ~n43261 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n28682 = ~n43271 | ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n28684 = ~n28683 | ~n28682;
  assign n28705 = ~n28685 & ~n28684;
  assign n28687 = ~n43251 | ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n28686 = ~n43242 | ~P1_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n28691 = ~n28687 | ~n28686;
  assign n28689 = ~n28775 | ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n28688 = ~n43275 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n28690 = ~n28689 | ~n28688;
  assign n28699 = ~n28691 & ~n28690;
  assign n28693 = ~n22907 | ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n28692 = ~n43246 | ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n28697 = ~n28693 | ~n28692;
  assign n28695 = ~n43245 | ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n28694 = ~n43265 | ~P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n28696 = ~n28695 | ~n28694;
  assign n28698 = ~n28697 & ~n28696;
  assign n28703 = ~n28699 | ~n28698;
  assign n28701 = ~n22908 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n28700 = ~n43264 | ~P1_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n28702 = ~n28701 | ~n28700;
  assign n28704 = ~n28703 & ~n28702;
  assign n28807 = ~n28705 | ~n28704;
  assign n28806 = ~n28707 & ~n28706;
  assign n28708 = n28807 ^ n28806;
  assign n28710 = ~n28708 | ~n28604;
  assign n28709 = ~n43721 | ~P1_EAX_REG_28__SCAN_IN;
  assign n28713 = ~n28710 | ~n28709;
  assign n28711 = ~P1_PHYADDRPOINTER_REG_28__SCAN_IN | ~n43722;
  assign n28712 = ~n43725 | ~n28711;
  assign n28716 = ~n28713 & ~n28712;
  assign n28718 = ~n40080 | ~P1_EBX_REG_28__SCAN_IN;
  assign n28717 = ~n40081 | ~P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n42979 = ~n28721 | ~n28720;
  assign P1_U2844 = n28727 | n28726;
  assign n42367 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n28730 = ~n28848 | ~n28728;
  assign n28733 = ~n28730 | ~n28729;
  assign n42828 = ~P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n43028 = ~n28733 & ~n28732;
  assign n28736 = ~n43709 | ~P1_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n28739 = ~n42834 | ~n28736;
  assign n28738 = ~n43713 & ~n28737;
  assign n28740 = ~n28739 & ~n28738;
  assign P1_U2975 = n28743 | n28742;
  assign n28750 = ~n41535 | ~n41259;
  assign n41117 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n41119 = ~n28757 | ~n41117;
  assign n28770 = ~n40529 | ~P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n41104 = ~n41145 | ~P3_REIP_REG_29__SCAN_IN;
  assign P3_U2833 = n28772 | n28771;
  assign n28777 = ~n28775 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n28776 = ~n43242 | ~P1_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n28781 = ~n28777 | ~n28776;
  assign n28779 = ~n22907 | ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n28778 = ~n22908 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n28780 = ~n28779 | ~n28778;
  assign n28789 = ~n28781 & ~n28780;
  assign n28783 = ~n43246 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n28782 = ~n43251 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n28787 = ~n28783 | ~n28782;
  assign n28785 = ~n43274 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n28784 = ~n43261 | ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n28786 = ~n28785 | ~n28784;
  assign n28788 = ~n28787 & ~n28786;
  assign n28805 = ~n28789 | ~n28788;
  assign n28791 = ~n43245 | ~P1_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n28790 = ~n22915 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n28795 = ~n28791 | ~n28790;
  assign n28793 = ~n43260 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n28792 = ~n43265 | ~P1_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n28794 = ~n28793 | ~n28792;
  assign n28803 = ~n28795 & ~n28794;
  assign n28797 = ~n43270 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n28796 = ~n43275 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n28801 = ~n28797 | ~n28796;
  assign n28799 = ~n43264 | ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n28798 = ~n43271 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n28800 = ~n28799 | ~n28798;
  assign n28802 = ~n28801 & ~n28800;
  assign n28804 = ~n28803 | ~n28802;
  assign n43240 = ~n28805 & ~n28804;
  assign n28808 = n43240 ^ n43239;
  assign n28815 = ~n28808 | ~n28604;
  assign n28809 = ~P1_EAX_REG_29__SCAN_IN;
  assign n28813 = ~n28810 & ~n28809;
  assign n28811 = ~P1_PHYADDRPOINTER_REG_29__SCAN_IN & ~n39944;
  assign n28812 = ~P1_STATE2_REG_2__SCAN_IN & ~n28811;
  assign n28814 = ~n28813 & ~n28812;
  assign n28818 = ~n28815 | ~n28814;
  assign n43720 = ~n28820 & ~n28819;
  assign n28821 = ~n28820 | ~n28819;
  assign n43120 = ~n28822 | ~n28821;
  assign n28824 = ~n40080 | ~P1_EBX_REG_29__SCAN_IN;
  assign n28823 = ~n40081 | ~P1_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign P1_U2843 = n28829 | n28828;
  assign n28831 = ~P1_EBX_REG_26__SCAN_IN | ~n43796;
  assign n29632 = ~P1_REIP_REG_26__SCAN_IN;
  assign n28830 = ~n43372 | ~n29632;
  assign n28843 = ~n28831 | ~n28830;
  assign n28837 = n42175 | n28860;
  assign n28836 = ~n43797 | ~P1_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n28846 = n28843 | n28842;
  assign n28876 = n42160 | n42400;
  assign P1_U2814 = n28846 | n28845;
  assign n41988 = ~P1_INSTADDRPOINTER_REG_25__SCAN_IN | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n28847 = ~n41988;
  assign n28849 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN & ~P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n28850 = ~n28849 | ~n43351;
  assign n28859 = ~n43709 | ~P1_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n28862 = ~n42935 | ~n28859;
  assign n28861 = ~n43713 & ~n28860;
  assign n28863 = ~n28862 & ~n28861;
  assign P1_U2973 = n28866 | n28865;
  assign n29674 = ~P1_REIP_REG_27__SCAN_IN;
  assign n28874 = ~n29674 & ~n29632;
  assign n28868 = n42175 | n43046;
  assign n28867 = ~n43797 | ~P1_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n28871 = ~n28870 & ~n28869;
  assign n28881 = n28886 | n28873;
  assign n28875 = ~n28874;
  assign n28878 = ~n43796 | ~P1_EBX_REG_28__SCAN_IN;
  assign P1_U2812 = n28881 | n28880;
  assign n28884 = ~P1_EBX_REG_29__SCAN_IN | ~n43796;
  assign n42488 = ~P1_REIP_REG_28__SCAN_IN;
  assign n43564 = ~P1_REIP_REG_29__SCAN_IN;
  assign n28883 = ~n43788 | ~n43564;
  assign n28892 = ~n43120 & ~n43794;
  assign n28888 = ~n41129 & ~n28885;
  assign n28887 = ~n43564 & ~n43567;
  assign n28890 = ~n28888 & ~n28887;
  assign n28889 = ~n43559 | ~n43138;
  assign n28893 = ~n28892 & ~n28891;
  assign P1_U2811 = n28896 | n28895;
  assign n28897 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_STATEBS16_REG_SCAN_IN;
  assign n28898 = ~n28897 | ~n39511;
  assign n28899 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_STATE2_REG_0__SCAN_IN;
  assign n28902 = ~n28898 | ~n28899;
  assign n28900 = ~n35802 & ~n28899;
  assign n28901 = ~n28900 | ~n39511;
  assign P2_U3178 = ~n28902 | ~n28901;
  assign n29541 = ~n31478 & ~n29055;
  assign n28906 = ~n29541 & ~n34515;
  assign n29750 = ~P1_STATE_REG_0__SCAN_IN | ~P1_REQUESTPENDING_REG_SCAN_IN;
  assign n29538 = ~P1_STATE_REG_1__SCAN_IN | ~HOLD;
  assign n28904 = ~n29750 | ~n29538;
  assign n28903 = ~HOLD | ~P1_STATE_REG_2__SCAN_IN;
  assign n28905 = ~n28904 | ~n28903;
  assign P1_U3195 = ~n28906 | ~n28905;
  assign n28950 = ~P2_STATE_REG_0__SCAN_IN;
  assign n29092 = ~P2_STATE_REG_1__SCAN_IN;
  assign n29095 = ~n28950 | ~n29092;
  assign n28907 = ~P2_STATE_REG_2__SCAN_IN & ~n29092;
  assign n28908 = ~P2_STATE_REG_0__SCAN_IN | ~n28907;
  assign n28937 = ~n29095 | ~n28908;
  assign n28909 = ~P2_STATE_REG_0__SCAN_IN | ~P2_ADS_N_REG_SCAN_IN;
  assign P2_U2815 = ~n28943 | ~n28909;
  assign n29150 = ~P3_STATE_REG_1__SCAN_IN;
  assign n28910 = ~n29150 & ~P3_STATE_REG_2__SCAN_IN;
  assign n28911 = ~n28910 | ~P3_STATE_REG_0__SCAN_IN;
  assign n29557 = ~n29149 | ~n29150;
  assign n28930 = ~n28911 | ~n29557;
  assign n28912 = ~P3_STATE_REG_0__SCAN_IN | ~P3_ADS_N_REG_SCAN_IN;
  assign P3_U2633 = ~n28934 | ~n28912;
  assign n29556 = ~n31667 & ~n29150;
  assign n29148 = ~n29556 & ~n29149;
  assign n28913 = ~P3_STATE_REG_1__SCAN_IN & ~n29749;
  assign n28914 = ~n29148 & ~n28913;
  assign n28920 = ~n28914 | ~P3_STATE_REG_2__SCAN_IN;
  assign n29560 = ~P3_REQUESTPENDING_REG_SCAN_IN & ~HOLD;
  assign n28918 = ~n29560 & ~n29149;
  assign n28915 = ~P3_STATE_REG_1__SCAN_IN & ~P3_REQUESTPENDING_REG_SCAN_IN;
  assign n29761 = ~HOLD;
  assign n29151 = ~n28928 & ~n29761;
  assign n29558 = ~n28915 & ~n29151;
  assign n28916 = ~n29556 | ~n29749;
  assign n28917 = ~n29558 | ~n28916;
  assign n28919 = ~n28918 | ~n28917;
  assign P3_U3031 = ~n28920 | ~n28919;
  assign n28921 = ~P2_STATE_REG_0__SCAN_IN | ~P2_REQUESTPENDING_REG_SCAN_IN;
  assign n28926 = ~HOLD & ~n28921;
  assign n29084 = ~n35802 | ~P2_STATE_REG_1__SCAN_IN;
  assign n29089 = ~P2_REQUESTPENDING_REG_SCAN_IN & ~HOLD;
  assign n28923 = ~n29089 & ~P2_STATE_REG_2__SCAN_IN;
  assign n28922 = ~n28921 | ~n29092;
  assign n28924 = ~n28923 | ~n28922;
  assign n28925 = ~n29084 | ~n28924;
  assign n28927 = ~n28926 & ~n28925;
  assign P2_U3210 = ~n28927 | ~n31819;
  assign n28932 = ~P3_DATAWIDTH_REG_0__SCAN_IN & ~n28930;
  assign n29057 = ~BS16;
  assign n29178 = ~n29150 | ~n28928;
  assign n28929 = ~n29057 | ~n29178;
  assign n28936 = ~n28930 | ~n28929;
  assign n28931 = ~n28936;
  assign P3_U3280 = ~n28932 & ~n28931;
  assign P2_U3205 = P2_DATAWIDTH_REG_5__SCAN_IN & n28943;
  assign P2_U3208 = P2_DATAWIDTH_REG_2__SCAN_IN & n28943;
  assign P2_U3204 = P2_DATAWIDTH_REG_6__SCAN_IN & n28943;
  assign P2_U3200 = P2_DATAWIDTH_REG_10__SCAN_IN & n28943;
  assign P2_U3199 = P2_DATAWIDTH_REG_11__SCAN_IN & n28943;
  assign P2_U3207 = P2_DATAWIDTH_REG_3__SCAN_IN & n28943;
  assign P2_U3197 = P2_DATAWIDTH_REG_13__SCAN_IN & n28943;
  assign P2_U3196 = P2_DATAWIDTH_REG_14__SCAN_IN & n28943;
  assign P2_U3203 = P2_DATAWIDTH_REG_7__SCAN_IN & n28943;
  assign P2_U3202 = P2_DATAWIDTH_REG_8__SCAN_IN & n28943;
  assign P2_U3201 = P2_DATAWIDTH_REG_9__SCAN_IN & n28943;
  assign P2_U3192 = P2_DATAWIDTH_REG_18__SCAN_IN & n28943;
  assign P2_U3191 = P2_DATAWIDTH_REG_19__SCAN_IN & n28943;
  assign P2_U3190 = P2_DATAWIDTH_REG_20__SCAN_IN & n28943;
  assign P2_U3206 = P2_DATAWIDTH_REG_4__SCAN_IN & n28943;
  assign P2_U3188 = P2_DATAWIDTH_REG_22__SCAN_IN & n28943;
  assign P2_U3187 = P2_DATAWIDTH_REG_23__SCAN_IN & n28943;
  assign P2_U3186 = P2_DATAWIDTH_REG_24__SCAN_IN & n28943;
  assign P2_U3185 = P2_DATAWIDTH_REG_25__SCAN_IN & n28943;
  assign P2_U3184 = P2_DATAWIDTH_REG_26__SCAN_IN & n28943;
  assign P2_U3183 = P2_DATAWIDTH_REG_27__SCAN_IN & n28943;
  assign P2_U3182 = P2_DATAWIDTH_REG_28__SCAN_IN & n28943;
  assign P2_U3181 = P2_DATAWIDTH_REG_29__SCAN_IN & n28943;
  assign P2_U3198 = P2_DATAWIDTH_REG_12__SCAN_IN & n28943;
  assign P2_U3180 = P2_DATAWIDTH_REG_30__SCAN_IN & n28943;
  assign P2_U3179 = P2_DATAWIDTH_REG_31__SCAN_IN & n28943;
  assign P2_U3195 = P2_DATAWIDTH_REG_15__SCAN_IN & n28943;
  assign P2_U3194 = P2_DATAWIDTH_REG_16__SCAN_IN & n28943;
  assign P2_U3193 = P2_DATAWIDTH_REG_17__SCAN_IN & n28943;
  assign P2_U3189 = P2_DATAWIDTH_REG_21__SCAN_IN & n28943;
  assign P3_U3000 = P3_DATAWIDTH_REG_30__SCAN_IN & n28934;
  assign P3_U3001 = P3_DATAWIDTH_REG_29__SCAN_IN & n28934;
  assign P3_U2999 = P3_DATAWIDTH_REG_31__SCAN_IN & n28934;
  assign P3_U3002 = P3_DATAWIDTH_REG_28__SCAN_IN & n28934;
  assign P3_U3003 = P3_DATAWIDTH_REG_27__SCAN_IN & n28934;
  assign P3_U3011 = P3_DATAWIDTH_REG_19__SCAN_IN & n28934;
  assign P3_U3016 = P3_DATAWIDTH_REG_14__SCAN_IN & n28934;
  assign P3_U3017 = P3_DATAWIDTH_REG_13__SCAN_IN & n28934;
  assign P3_U3018 = P3_DATAWIDTH_REG_12__SCAN_IN & n28934;
  assign P3_U3019 = P3_DATAWIDTH_REG_11__SCAN_IN & n28934;
  assign P3_U3004 = P3_DATAWIDTH_REG_26__SCAN_IN & n28934;
  assign P3_U3005 = P3_DATAWIDTH_REG_25__SCAN_IN & n28934;
  assign P3_U3022 = P3_DATAWIDTH_REG_8__SCAN_IN & n28934;
  assign P3_U3007 = P3_DATAWIDTH_REG_23__SCAN_IN & n28934;
  assign P3_U3008 = P3_DATAWIDTH_REG_22__SCAN_IN & n28934;
  assign P3_U3009 = P3_DATAWIDTH_REG_21__SCAN_IN & n28934;
  assign P3_U3010 = P3_DATAWIDTH_REG_20__SCAN_IN & n28934;
  assign P3_U3012 = P3_DATAWIDTH_REG_18__SCAN_IN & n28934;
  assign P3_U3013 = P3_DATAWIDTH_REG_17__SCAN_IN & n28934;
  assign P3_U3014 = P3_DATAWIDTH_REG_16__SCAN_IN & n28934;
  assign P3_U3015 = P3_DATAWIDTH_REG_15__SCAN_IN & n28934;
  assign P3_U3027 = P3_DATAWIDTH_REG_3__SCAN_IN & n28934;
  assign P3_U3023 = P3_DATAWIDTH_REG_7__SCAN_IN & n28934;
  assign P3_U3028 = P3_DATAWIDTH_REG_2__SCAN_IN & n28934;
  assign P3_U3025 = P3_DATAWIDTH_REG_5__SCAN_IN & n28934;
  assign P3_U3006 = P3_DATAWIDTH_REG_24__SCAN_IN & n28934;
  assign P3_U3021 = P3_DATAWIDTH_REG_9__SCAN_IN & n28934;
  assign P3_U3020 = P3_DATAWIDTH_REG_10__SCAN_IN & n28934;
  assign P3_U3024 = P3_DATAWIDTH_REG_6__SCAN_IN & n28934;
  assign P3_U3026 = P3_DATAWIDTH_REG_4__SCAN_IN & n28934;
  assign n28933 = ~P3_STATEBS16_REG_SCAN_IN | ~n28934;
  assign P3_U2636 = ~n28936 | ~n28933;
  assign n28935 = ~P3_DATAWIDTH_REG_1__SCAN_IN | ~n28934;
  assign P3_U3281 = ~n28936 | ~n28935;
  assign n28938 = ~P2_DATAWIDTH_REG_1__SCAN_IN & ~n28937;
  assign n28939 = ~n29057 | ~n28937;
  assign n28942 = ~n29085 & ~n28939;
  assign P2_U3592 = ~n28938 & ~n28942;
  assign n28940 = ~n28943 | ~n38321;
  assign n28941 = ~n28940 | ~n28939;
  assign n29164 = ~n29085 | ~n28950;
  assign P2_U2818 = ~n28941 | ~n29164;
  assign n28945 = ~n28942;
  assign n28944 = ~P2_DATAWIDTH_REG_0__SCAN_IN | ~n28943;
  assign P2_U3591 = ~n28945 | ~n28944;
  assign n41672 = ~n41671 & ~n31507;
  assign n28948 = ~n41671 & ~n42016;
  assign n28946 = ~P3_STATE2_REG_0__SCAN_IN & ~P3_STATEBS16_REG_SCAN_IN;
  assign n32843 = ~n28946 | ~n40527;
  assign n28947 = ~n32843;
  assign n41380 = ~n28948 & ~n28947;
  assign n42012 = ~n40527 | ~n35452;
  assign n28949 = ~n41380 | ~n42012;
  assign P3_U2998 = ~n41672 & ~n28949;
  assign n29175 = P2_STATE_REG_1__SCAN_IN & n28950;
  assign n28952 = ~P2_BE_N_REG_0__SCAN_IN | ~n29553;
  assign n28951 = ~P2_BYTEENABLE_REG_0__SCAN_IN | ~n29175;
  assign P2_U3588 = ~n28952 | ~n28951;
  assign n28954 = ~P2_BE_N_REG_1__SCAN_IN | ~n29553;
  assign n28953 = ~P2_BYTEENABLE_REG_1__SCAN_IN | ~n29175;
  assign P2_U3587 = ~n28954 | ~n28953;
  assign n28956 = ~P2_M_IO_N_REG_SCAN_IN | ~n29553;
  assign n28955 = ~P2_MEMORYFETCH_REG_SCAN_IN | ~n29175;
  assign P2_U3611 = ~n28956 | ~n28955;
  assign n28958 = ~n29749 & ~P2_STATE_REG_0__SCAN_IN;
  assign n28957 = ~n29761 & ~n29085;
  assign n28959 = ~n28958 & ~n28957;
  assign n28960 = ~P2_REQUESTPENDING_REG_SCAN_IN | ~n28959;
  assign n28962 = ~n28960 | ~n29553;
  assign n29093 = ~P2_STATE_REG_0__SCAN_IN | ~n29084;
  assign n29174 = ~P2_STATE_REG_2__SCAN_IN;
  assign n28961 = ~n29093 | ~n29174;
  assign P2_U3209 = ~n28962 | ~n28961;
  assign n28964 = ~P2_BE_N_REG_2__SCAN_IN | ~n29553;
  assign n28963 = ~P2_BYTEENABLE_REG_2__SCAN_IN | ~n29175;
  assign P2_U3586 = ~n28964 | ~n28963;
  assign n28966 = ~P2_BE_N_REG_3__SCAN_IN | ~n29553;
  assign n28965 = ~P2_BYTEENABLE_REG_3__SCAN_IN | ~n29175;
  assign P2_U3585 = ~n28966 | ~n28965;
  assign n28968 = ~P1_DATAWIDTH_REG_30__SCAN_IN & ~P1_DATAWIDTH_REG_31__SCAN_IN;
  assign n28967 = ~P1_DATAWIDTH_REG_28__SCAN_IN & ~P1_DATAWIDTH_REG_29__SCAN_IN;
  assign n28972 = ~n28968 | ~n28967;
  assign n28970 = ~P1_DATAWIDTH_REG_18__SCAN_IN & ~P1_DATAWIDTH_REG_19__SCAN_IN;
  assign n28969 = ~P1_DATAWIDTH_REG_16__SCAN_IN & ~P1_DATAWIDTH_REG_17__SCAN_IN;
  assign n28971 = ~n28970 | ~n28969;
  assign n28980 = ~n28972 & ~n28971;
  assign n28974 = ~P1_DATAWIDTH_REG_26__SCAN_IN & ~P1_DATAWIDTH_REG_27__SCAN_IN;
  assign n28973 = ~P1_DATAWIDTH_REG_24__SCAN_IN & ~P1_DATAWIDTH_REG_25__SCAN_IN;
  assign n28978 = ~n28974 | ~n28973;
  assign n28976 = ~P1_DATAWIDTH_REG_22__SCAN_IN & ~P1_DATAWIDTH_REG_23__SCAN_IN;
  assign n28975 = ~P1_DATAWIDTH_REG_20__SCAN_IN & ~P1_DATAWIDTH_REG_21__SCAN_IN;
  assign n28977 = ~n28976 | ~n28975;
  assign n28979 = ~n28978 & ~n28977;
  assign n28996 = ~n28980 | ~n28979;
  assign n28982 = ~P1_DATAWIDTH_REG_14__SCAN_IN & ~P1_DATAWIDTH_REG_15__SCAN_IN;
  assign n28981 = ~P1_DATAWIDTH_REG_12__SCAN_IN & ~P1_DATAWIDTH_REG_13__SCAN_IN;
  assign n28986 = ~n28982 | ~n28981;
  assign n28984 = ~P1_DATAWIDTH_REG_3__SCAN_IN & ~P1_DATAWIDTH_REG_2__SCAN_IN;
  assign n28983 = ~P1_DATAWIDTH_REG_0__SCAN_IN | ~P1_DATAWIDTH_REG_1__SCAN_IN;
  assign n28985 = ~n28984 | ~n28983;
  assign n28994 = ~n28986 & ~n28985;
  assign n28988 = ~P1_DATAWIDTH_REG_10__SCAN_IN & ~P1_DATAWIDTH_REG_11__SCAN_IN;
  assign n28987 = ~P1_DATAWIDTH_REG_8__SCAN_IN & ~P1_DATAWIDTH_REG_9__SCAN_IN;
  assign n28992 = ~n28988 | ~n28987;
  assign n28990 = ~P1_DATAWIDTH_REG_6__SCAN_IN & ~P1_DATAWIDTH_REG_7__SCAN_IN;
  assign n28989 = ~P1_DATAWIDTH_REG_4__SCAN_IN & ~P1_DATAWIDTH_REG_5__SCAN_IN;
  assign n28991 = ~n28990 | ~n28989;
  assign n28993 = ~n28992 & ~n28991;
  assign n28995 = ~n28994 | ~n28993;
  assign n29075 = ~n28996 & ~n28995;
  assign n29077 = ~n29075;
  assign n29004 = ~P1_BYTEENABLE_REG_2__SCAN_IN | ~n29077;
  assign n29001 = ~P1_REIP_REG_0__SCAN_IN | ~P1_REIP_REG_1__SCAN_IN;
  assign n31686 = ~P1_REIP_REG_0__SCAN_IN;
  assign n28998 = ~P1_DATAWIDTH_REG_0__SCAN_IN | ~n31686;
  assign n29043 = ~P1_DATAWIDTH_REG_1__SCAN_IN & ~P1_DATAWIDTH_REG_0__SCAN_IN;
  assign n28997 = ~n29043;
  assign n28999 = ~n28998 | ~n28997;
  assign n35494 = ~P1_REIP_REG_1__SCAN_IN;
  assign n29000 = ~n28999 | ~n35494;
  assign n29002 = ~n29001 | ~n29000;
  assign n29003 = ~n29002 | ~n29075;
  assign P1_U3481 = ~n29004 | ~n29003;
  assign n29006 = ~P3_DATAWIDTH_REG_30__SCAN_IN & ~P3_DATAWIDTH_REG_31__SCAN_IN;
  assign n29005 = ~P3_DATAWIDTH_REG_28__SCAN_IN & ~P3_DATAWIDTH_REG_29__SCAN_IN;
  assign n29010 = ~n29006 | ~n29005;
  assign n29008 = ~P3_DATAWIDTH_REG_18__SCAN_IN & ~P3_DATAWIDTH_REG_19__SCAN_IN;
  assign n29007 = ~P3_DATAWIDTH_REG_16__SCAN_IN & ~P3_DATAWIDTH_REG_17__SCAN_IN;
  assign n29009 = ~n29008 | ~n29007;
  assign n29018 = ~n29010 & ~n29009;
  assign n29012 = ~P3_DATAWIDTH_REG_26__SCAN_IN & ~P3_DATAWIDTH_REG_27__SCAN_IN;
  assign n29011 = ~P3_DATAWIDTH_REG_24__SCAN_IN & ~P3_DATAWIDTH_REG_25__SCAN_IN;
  assign n29016 = ~n29012 | ~n29011;
  assign n29014 = ~P3_DATAWIDTH_REG_22__SCAN_IN & ~P3_DATAWIDTH_REG_23__SCAN_IN;
  assign n29013 = ~P3_DATAWIDTH_REG_20__SCAN_IN & ~P3_DATAWIDTH_REG_21__SCAN_IN;
  assign n29015 = ~n29014 | ~n29013;
  assign n29017 = ~n29016 & ~n29015;
  assign n29034 = ~n29018 | ~n29017;
  assign n29020 = ~P3_DATAWIDTH_REG_14__SCAN_IN & ~P3_DATAWIDTH_REG_15__SCAN_IN;
  assign n29019 = ~P3_DATAWIDTH_REG_12__SCAN_IN & ~P3_DATAWIDTH_REG_13__SCAN_IN;
  assign n29024 = ~n29020 | ~n29019;
  assign n29022 = ~P3_DATAWIDTH_REG_3__SCAN_IN & ~P3_DATAWIDTH_REG_2__SCAN_IN;
  assign n29021 = ~P3_DATAWIDTH_REG_0__SCAN_IN | ~P3_DATAWIDTH_REG_1__SCAN_IN;
  assign n29023 = ~n29022 | ~n29021;
  assign n29032 = ~n29024 & ~n29023;
  assign n29026 = ~P3_DATAWIDTH_REG_10__SCAN_IN & ~P3_DATAWIDTH_REG_11__SCAN_IN;
  assign n29025 = ~P3_DATAWIDTH_REG_8__SCAN_IN & ~P3_DATAWIDTH_REG_9__SCAN_IN;
  assign n29030 = ~n29026 | ~n29025;
  assign n29028 = ~P3_DATAWIDTH_REG_6__SCAN_IN & ~P3_DATAWIDTH_REG_7__SCAN_IN;
  assign n29027 = ~P3_DATAWIDTH_REG_4__SCAN_IN & ~P3_DATAWIDTH_REG_5__SCAN_IN;
  assign n29029 = ~n29028 | ~n29027;
  assign n29031 = ~n29030 & ~n29029;
  assign n29033 = ~n29032 | ~n29031;
  assign n29070 = ~n29034 & ~n29033;
  assign n29072 = ~n29070;
  assign n29042 = ~P3_BYTEENABLE_REG_2__SCAN_IN | ~n29072;
  assign n29039 = ~P3_REIP_REG_0__SCAN_IN | ~P3_REIP_REG_1__SCAN_IN;
  assign n29069 = ~P3_REIP_REG_0__SCAN_IN;
  assign n29036 = ~P3_DATAWIDTH_REG_0__SCAN_IN | ~n29069;
  assign n29048 = ~P3_DATAWIDTH_REG_1__SCAN_IN & ~P3_DATAWIDTH_REG_0__SCAN_IN;
  assign n29035 = ~n29048;
  assign n29037 = ~n29036 | ~n29035;
  assign n35979 = ~P3_REIP_REG_1__SCAN_IN;
  assign n29038 = ~n29037 | ~n35979;
  assign n29040 = ~n29039 | ~n29038;
  assign n29041 = ~n29040 | ~n29070;
  assign P3_U3292 = ~n29042 | ~n29041;
  assign n29047 = ~P1_BYTEENABLE_REG_3__SCAN_IN | ~n29077;
  assign n29044 = P1_REIP_REG_1__SCAN_IN | P1_DATAWIDTH_REG_1__SCAN_IN;
  assign n29061 = ~n29043 | ~n31686;
  assign n29045 = ~n29044 | ~n29061;
  assign n29046 = ~n29045 | ~n29075;
  assign P1_U2808 = ~n29047 | ~n29046;
  assign n29052 = ~P3_BYTEENABLE_REG_3__SCAN_IN | ~n29072;
  assign n29049 = P3_REIP_REG_1__SCAN_IN | P3_DATAWIDTH_REG_1__SCAN_IN;
  assign n29065 = ~n29048 | ~n29069;
  assign n29050 = ~n29049 | ~n29065;
  assign n29051 = ~n29050 | ~n29070;
  assign P3_U2639 = ~n29052 | ~n29051;
  assign n29054 = ~n29055 & ~P1_STATE_REG_2__SCAN_IN;
  assign n29053 = ~P1_STATE_REG_0__SCAN_IN;
  assign n29056 = ~n29054 & ~n29053;
  assign n29058 = ~n29056 & ~n29580;
  assign n29060 = ~P1_DATAWIDTH_REG_0__SCAN_IN & ~n29058;
  assign n29059 = n29057 & n29574;
  assign n29080 = ~n29059 & ~n29461;
  assign P1_U3464 = ~n29060 & ~n29080;
  assign n29062 = ~n35494 | ~n29061;
  assign n29064 = ~n29062 | ~n29075;
  assign n29063 = ~P1_BYTEENABLE_REG_1__SCAN_IN | ~n29077;
  assign P1_U2807 = ~n29064 | ~n29063;
  assign n29066 = ~n35979 | ~n29065;
  assign n29068 = ~n29066 | ~n29070;
  assign n29067 = ~P3_BYTEENABLE_REG_1__SCAN_IN | ~n29072;
  assign P3_U2638 = ~n29068 | ~n29067;
  assign n29071 = ~n35979 | ~n29069;
  assign n29074 = ~n29071 | ~n29070;
  assign n29073 = ~P3_BYTEENABLE_REG_0__SCAN_IN | ~n29072;
  assign P3_U3293 = ~n29074 | ~n29073;
  assign n29076 = ~n35494 | ~n31686;
  assign n29079 = ~n29076 | ~n29075;
  assign n29078 = ~P1_BYTEENABLE_REG_0__SCAN_IN | ~n29077;
  assign P1_U3482 = ~n29079 | ~n29078;
  assign n29083 = ~n29080;
  assign n29081 = ~P1_DATAWIDTH_REG_1__SCAN_IN | ~n29461;
  assign P1_U3465 = ~n29083 | ~n29081;
  assign n29082 = ~P1_STATEBS16_REG_SCAN_IN | ~n29461;
  assign P1_U2805 = ~n29083 | ~n29082;
  assign P1_U3164 = P1_DATAWIDTH_REG_31__SCAN_IN & n29461;
  assign P1_U3165 = P1_DATAWIDTH_REG_30__SCAN_IN & n29461;
  assign P1_U3172 = P1_DATAWIDTH_REG_23__SCAN_IN & n29461;
  assign P1_U3171 = P1_DATAWIDTH_REG_24__SCAN_IN & n29461;
  assign P1_U3173 = P1_DATAWIDTH_REG_22__SCAN_IN & n29461;
  assign P1_U3169 = P1_DATAWIDTH_REG_26__SCAN_IN & n29461;
  assign P1_U3170 = P1_DATAWIDTH_REG_25__SCAN_IN & n29461;
  assign P1_U3174 = P1_DATAWIDTH_REG_21__SCAN_IN & n29461;
  assign P1_U3175 = P1_DATAWIDTH_REG_20__SCAN_IN & n29461;
  assign P1_U3176 = P1_DATAWIDTH_REG_19__SCAN_IN & n29461;
  assign P1_U3177 = P1_DATAWIDTH_REG_18__SCAN_IN & n29461;
  assign P1_U3166 = P1_DATAWIDTH_REG_29__SCAN_IN & n29461;
  assign P1_U3167 = P1_DATAWIDTH_REG_28__SCAN_IN & n29461;
  assign P1_U3168 = P1_DATAWIDTH_REG_27__SCAN_IN & n29461;
  assign P1_U3181 = P1_DATAWIDTH_REG_14__SCAN_IN & n29461;
  assign P1_U3182 = P1_DATAWIDTH_REG_13__SCAN_IN & n29461;
  assign P1_U3183 = P1_DATAWIDTH_REG_12__SCAN_IN & n29461;
  assign P1_U3184 = P1_DATAWIDTH_REG_11__SCAN_IN & n29461;
  assign P1_U3185 = P1_DATAWIDTH_REG_10__SCAN_IN & n29461;
  assign P1_U3186 = P1_DATAWIDTH_REG_9__SCAN_IN & n29461;
  assign P1_U3187 = P1_DATAWIDTH_REG_8__SCAN_IN & n29461;
  assign P1_U3188 = P1_DATAWIDTH_REG_7__SCAN_IN & n29461;
  assign P1_U3189 = P1_DATAWIDTH_REG_6__SCAN_IN & n29461;
  assign P1_U3190 = P1_DATAWIDTH_REG_5__SCAN_IN & n29461;
  assign P1_U3191 = P1_DATAWIDTH_REG_4__SCAN_IN & n29461;
  assign P1_U3193 = P1_DATAWIDTH_REG_2__SCAN_IN & n29461;
  assign P1_U3178 = P1_DATAWIDTH_REG_17__SCAN_IN & n29461;
  assign P1_U3179 = P1_DATAWIDTH_REG_16__SCAN_IN & n29461;
  assign P1_U3180 = P1_DATAWIDTH_REG_15__SCAN_IN & n29461;
  assign P1_U3192 = P1_DATAWIDTH_REG_3__SCAN_IN & n29461;
  assign n29088 = ~n29084 & ~NA;
  assign n29086 = ~n29085;
  assign n29087 = ~n29086 & ~P2_REQUESTPENDING_REG_SCAN_IN;
  assign n29090 = ~n29088 & ~n29087;
  assign n29091 = ~n29090 & ~n29089;
  assign n29100 = ~P2_STATE_REG_0__SCAN_IN | ~n29091;
  assign n29094 = ~NA | ~n29092;
  assign n29097 = ~n29094 | ~n29093;
  assign n29096 = ~HOLD | ~n29095;
  assign n29098 = ~n29097 | ~n29096;
  assign n29099 = ~P2_STATE_REG_2__SCAN_IN | ~n29098;
  assign P2_U3211 = ~n29100 | ~n29099;
  assign n29102 = ~P2_DATAWIDTH_REG_30__SCAN_IN & ~P2_DATAWIDTH_REG_31__SCAN_IN;
  assign n29101 = ~P2_DATAWIDTH_REG_28__SCAN_IN & ~P2_DATAWIDTH_REG_29__SCAN_IN;
  assign n29106 = ~n29102 | ~n29101;
  assign n29104 = ~P2_DATAWIDTH_REG_18__SCAN_IN & ~P2_DATAWIDTH_REG_19__SCAN_IN;
  assign n29103 = ~P2_DATAWIDTH_REG_16__SCAN_IN & ~P2_DATAWIDTH_REG_17__SCAN_IN;
  assign n29105 = ~n29104 | ~n29103;
  assign n29114 = ~n29106 & ~n29105;
  assign n29108 = ~P2_DATAWIDTH_REG_26__SCAN_IN & ~P2_DATAWIDTH_REG_27__SCAN_IN;
  assign n29107 = ~P2_DATAWIDTH_REG_24__SCAN_IN & ~P2_DATAWIDTH_REG_25__SCAN_IN;
  assign n29112 = ~n29108 | ~n29107;
  assign n29110 = ~P2_DATAWIDTH_REG_22__SCAN_IN & ~P2_DATAWIDTH_REG_23__SCAN_IN;
  assign n29109 = ~P2_DATAWIDTH_REG_20__SCAN_IN & ~P2_DATAWIDTH_REG_21__SCAN_IN;
  assign n29111 = ~n29110 | ~n29109;
  assign n29113 = ~n29112 & ~n29111;
  assign n29130 = ~n29114 | ~n29113;
  assign n29116 = ~P2_DATAWIDTH_REG_14__SCAN_IN & ~P2_DATAWIDTH_REG_15__SCAN_IN;
  assign n29115 = ~P2_DATAWIDTH_REG_12__SCAN_IN & ~P2_DATAWIDTH_REG_13__SCAN_IN;
  assign n29120 = ~n29116 | ~n29115;
  assign n29118 = ~P2_DATAWIDTH_REG_3__SCAN_IN & ~P2_DATAWIDTH_REG_2__SCAN_IN;
  assign n29117 = ~P2_DATAWIDTH_REG_0__SCAN_IN | ~P2_DATAWIDTH_REG_1__SCAN_IN;
  assign n29119 = ~n29118 | ~n29117;
  assign n29128 = ~n29120 & ~n29119;
  assign n29122 = ~P2_DATAWIDTH_REG_10__SCAN_IN & ~P2_DATAWIDTH_REG_11__SCAN_IN;
  assign n29121 = ~P2_DATAWIDTH_REG_8__SCAN_IN & ~P2_DATAWIDTH_REG_9__SCAN_IN;
  assign n29126 = ~n29122 | ~n29121;
  assign n29124 = ~P2_DATAWIDTH_REG_6__SCAN_IN & ~P2_DATAWIDTH_REG_7__SCAN_IN;
  assign n29123 = ~P2_DATAWIDTH_REG_4__SCAN_IN & ~P2_DATAWIDTH_REG_5__SCAN_IN;
  assign n29125 = ~n29124 | ~n29123;
  assign n29127 = ~n29126 & ~n29125;
  assign n29129 = ~n29128 | ~n29127;
  assign n29233 = ~n29130 & ~n29129;
  assign n29133 = ~n29233 & ~P2_BYTEENABLE_REG_1__SCAN_IN;
  assign n29166 = ~n29233 | ~n29550;
  assign n29131 = P2_DATAWIDTH_REG_1__SCAN_IN | P2_DATAWIDTH_REG_0__SCAN_IN;
  assign n29168 = ~P2_REIP_REG_0__SCAN_IN & ~n29131;
  assign n29132 = ~n29166 & ~n29168;
  assign P2_U2821 = ~n29133 & ~n29132;
  assign n29135 = ~n29233 & ~P2_BYTEENABLE_REG_0__SCAN_IN;
  assign n29134 = ~n29166 & ~P2_REIP_REG_0__SCAN_IN;
  assign P2_U2820 = ~n29135 & ~n29134;
  assign n29137 = ~P2_W_R_N_REG_SCAN_IN | ~n29553;
  assign n29136 = P2_READREQUEST_REG_SCAN_IN | n29553;
  assign P2_U3608 = ~n29137 | ~n29136;
  assign n29139 = ~P3_BE_N_REG_2__SCAN_IN | ~n29439;
  assign n29138 = ~n29308 | ~P3_BYTEENABLE_REG_2__SCAN_IN;
  assign P3_U3275 = ~n29139 | ~n29138;
  assign n29141 = ~P3_BE_N_REG_1__SCAN_IN | ~n29439;
  assign n29140 = ~n29308 | ~P3_BYTEENABLE_REG_1__SCAN_IN;
  assign P3_U3276 = ~n29141 | ~n29140;
  assign n29143 = ~P3_BE_N_REG_0__SCAN_IN | ~n29439;
  assign n29142 = ~n29308 | ~P3_BYTEENABLE_REG_0__SCAN_IN;
  assign P3_U3277 = ~n29143 | ~n29142;
  assign n29145 = ~P3_M_IO_N_REG_SCAN_IN | ~n29439;
  assign n29144 = ~n29308 | ~P3_MEMORYFETCH_REG_SCAN_IN;
  assign P3_U3297 = ~n29145 | ~n29144;
  assign n29147 = ~P3_BE_N_REG_3__SCAN_IN | ~n29439;
  assign n29146 = ~n29308 | ~P3_BYTEENABLE_REG_3__SCAN_IN;
  assign P3_U3274 = ~n29147 | ~n29146;
  assign n29159 = P3_STATE_REG_2__SCAN_IN | n29148;
  assign n29156 = ~NA | ~n29149;
  assign n29154 = ~n29150 & ~n29761;
  assign n29152 = ~n29151;
  assign n29153 = ~P3_REQUESTPENDING_REG_SCAN_IN | ~n29152;
  assign n29155 = ~n29154 & ~n29153;
  assign n29157 = ~n29156 | ~n29155;
  assign n29158 = ~n29157 | ~n29439;
  assign P3_U3029 = ~n29159 | ~n29158;
  assign n29161 = ~P3_W_R_N_REG_SCAN_IN | ~n29439;
  assign n29160 = P3_READREQUEST_REG_SCAN_IN | n29439;
  assign P3_U3294 = ~n29161 | ~n29160;
  assign n29163 = ~P2_CODEFETCH_REG_SCAN_IN & ~n29553;
  assign n29162 = P2_D_C_N_REG_SCAN_IN & n29553;
  assign n29165 = ~n29163 & ~n29162;
  assign P2_U2817 = ~n29165 | ~n29164;
  assign n29235 = ~n29233;
  assign n29167 = P2_BYTEENABLE_REG_3__SCAN_IN & n29235;
  assign n29231 = ~P2_DATAWIDTH_REG_1__SCAN_IN & ~n29166;
  assign n29170 = ~n29167 & ~n29231;
  assign n29169 = ~n29233 | ~n29168;
  assign P2_U2823 = ~n29170 | ~n29169;
  assign n29173 = ~n29171 & ~n29175;
  assign n29549 = ~P2_STATE_REG_2__SCAN_IN | ~n29175;
  assign n29172 = ~n29484 & ~n29549;
  assign n29177 = ~n29173 & ~n29172;
  assign n29226 = ~n29175 | ~n29174;
  assign n29176 = ~P2_REIP_REG_31__SCAN_IN | ~n29462;
  assign P2_U3241 = ~n29177 | ~n29176;
  assign n29180 = ~n29178 & ~P3_STATE_REG_0__SCAN_IN;
  assign n29179 = ~n29439 & ~P3_CODEFETCH_REG_SCAN_IN;
  assign n29182 = ~n29180 & ~n29179;
  assign n29181 = ~P3_D_C_N_REG_SCAN_IN | ~n29439;
  assign P3_U2635 = ~n29182 | ~n29181;
  assign n29184 = ~n27915 & ~n29226;
  assign n29183 = ~n29204 & ~n29549;
  assign n29186 = ~n29184 & ~n29183;
  assign n29185 = ~P2_ADDRESS_REG_8__SCAN_IN | ~n29553;
  assign P2_U3220 = ~n29186 | ~n29185;
  assign n29188 = ~n28229 & ~n29226;
  assign n29187 = ~n27915 & ~n29549;
  assign n29190 = ~n29188 & ~n29187;
  assign n29189 = ~P2_ADDRESS_REG_9__SCAN_IN | ~n29553;
  assign P2_U3221 = ~n29190 | ~n29189;
  assign n29192 = ~n27901 & ~n29226;
  assign n29191 = ~n29199 & ~n29549;
  assign n29194 = ~n29192 & ~n29191;
  assign n29193 = ~P2_ADDRESS_REG_6__SCAN_IN | ~n29553;
  assign P2_U3218 = ~n29194 | ~n29193;
  assign n29196 = ~n26522 & ~n29226;
  assign n29195 = ~n38814 & ~n29549;
  assign n29198 = ~n29196 & ~n29195;
  assign n29197 = ~P2_ADDRESS_REG_2__SCAN_IN | ~n29553;
  assign P2_U3214 = ~n29198 | ~n29197;
  assign n29201 = ~n29199 & ~n29226;
  assign n29200 = ~n26537 & ~n29549;
  assign n29203 = ~n29201 & ~n29200;
  assign n29202 = ~P2_ADDRESS_REG_5__SCAN_IN | ~n29553;
  assign P2_U3217 = ~n29203 | ~n29202;
  assign n29206 = ~n29204 & ~n29226;
  assign n29205 = ~n27901 & ~n29549;
  assign n29208 = ~n29206 & ~n29205;
  assign n29207 = ~P2_ADDRESS_REG_7__SCAN_IN | ~n29553;
  assign P2_U3219 = ~n29208 | ~n29207;
  assign n29210 = ~n28249 & ~n29226;
  assign n29209 = ~n29221 & ~n29549;
  assign n29212 = ~n29210 & ~n29209;
  assign n29211 = ~P2_ADDRESS_REG_12__SCAN_IN | ~n29553;
  assign P2_U3224 = ~n29212 | ~n29211;
  assign n29214 = ~n28236 & ~n29226;
  assign n29213 = ~n28229 & ~n29549;
  assign n29216 = ~n29214 & ~n29213;
  assign n29215 = ~P2_ADDRESS_REG_10__SCAN_IN | ~n29553;
  assign P2_U3222 = ~n29216 | ~n29215;
  assign n29218 = ~n26530 & ~n29226;
  assign n29217 = ~n26522 & ~n29549;
  assign n29220 = ~n29218 & ~n29217;
  assign n29219 = ~P2_ADDRESS_REG_3__SCAN_IN | ~n29553;
  assign P2_U3215 = ~n29220 | ~n29219;
  assign n29223 = ~n29221 & ~n29226;
  assign n29222 = ~n28236 & ~n29549;
  assign n29225 = ~n29223 & ~n29222;
  assign n29224 = ~P2_ADDRESS_REG_11__SCAN_IN | ~n29553;
  assign P2_U3223 = ~n29225 | ~n29224;
  assign n29228 = ~n26537 & ~n29226;
  assign n29227 = ~n26530 & ~n29549;
  assign n29230 = ~n29228 & ~n29227;
  assign n29229 = ~P2_ADDRESS_REG_4__SCAN_IN | ~n29553;
  assign P2_U3216 = ~n29230 | ~n29229;
  assign n29232 = ~P2_REIP_REG_0__SCAN_IN | ~P2_DATAWIDTH_REG_0__SCAN_IN;
  assign n29239 = ~n29232 | ~n29231;
  assign n29234 = ~P2_REIP_REG_0__SCAN_IN | ~n29233;
  assign n29237 = ~n29550 & ~n29234;
  assign n29236 = P2_BYTEENABLE_REG_2__SCAN_IN & n29235;
  assign n29238 = ~n29237 & ~n29236;
  assign P2_U2822 = ~n29239 | ~n29238;
  assign n29240 = ~P3_DATAO_REG_30__SCAN_IN;
  assign n29243 = ~n29240 & ~P3_DATAO_REG_31__SCAN_IN;
  assign n29241 = ~P1_DATAO_REG_30__SCAN_IN;
  assign n29242 = ~n29241 & ~P1_DATAO_REG_31__SCAN_IN;
  assign n29245 = ~n29243 & ~n29242;
  assign n31168 = ~P2_DATAO_REG_31__SCAN_IN;
  assign n29244 = ~P2_DATAO_REG_30__SCAN_IN | ~n31168;
  assign n29247 = ~P2_ADDRESS_REG_21__SCAN_IN | ~n29304;
  assign n29246 = ~n29305 | ~P3_ADDRESS_REG_21__SCAN_IN;
  assign U363 = ~n29247 | ~n29246;
  assign n29249 = ~P2_ADDRESS_REG_18__SCAN_IN | ~n29304;
  assign n29248 = ~n29305 | ~P3_ADDRESS_REG_18__SCAN_IN;
  assign U367 = ~n29249 | ~n29248;
  assign n29251 = ~P2_ADDRESS_REG_19__SCAN_IN | ~n29304;
  assign n29250 = ~n29305 | ~P3_ADDRESS_REG_19__SCAN_IN;
  assign U366 = ~n29251 | ~n29250;
  assign n29253 = ~P2_ADDRESS_REG_22__SCAN_IN | ~n29304;
  assign n29252 = ~n29305 | ~P3_ADDRESS_REG_22__SCAN_IN;
  assign U362 = ~n29253 | ~n29252;
  assign n29255 = ~P2_ADDRESS_REG_20__SCAN_IN | ~n29304;
  assign n29254 = ~n29305 | ~P3_ADDRESS_REG_20__SCAN_IN;
  assign U364 = ~n29255 | ~n29254;
  assign n29257 = ~P2_ADDRESS_REG_25__SCAN_IN | ~n29304;
  assign n29256 = ~n29305 | ~P3_ADDRESS_REG_25__SCAN_IN;
  assign U359 = ~n29257 | ~n29256;
  assign n29259 = ~P2_ADDRESS_REG_9__SCAN_IN | ~n29304;
  assign n29258 = ~n29305 | ~P3_ADDRESS_REG_9__SCAN_IN;
  assign U347 = ~n29259 | ~n29258;
  assign n29261 = ~P2_ADDRESS_REG_8__SCAN_IN | ~n29304;
  assign n29260 = ~n29305 | ~P3_ADDRESS_REG_8__SCAN_IN;
  assign U348 = ~n29261 | ~n29260;
  assign n29263 = ~P2_ADDRESS_REG_17__SCAN_IN | ~n29304;
  assign n29262 = ~n29305 | ~P3_ADDRESS_REG_17__SCAN_IN;
  assign U368 = ~n29263 | ~n29262;
  assign n29265 = ~P2_ADDRESS_REG_11__SCAN_IN | ~n29304;
  assign n29264 = ~n29305 | ~P3_ADDRESS_REG_11__SCAN_IN;
  assign U374 = ~n29265 | ~n29264;
  assign n29267 = ~P2_ADDRESS_REG_10__SCAN_IN | ~n29304;
  assign n29266 = ~n29305 | ~P3_ADDRESS_REG_10__SCAN_IN;
  assign U375 = ~n29267 | ~n29266;
  assign n29269 = ~P2_ADDRESS_REG_28__SCAN_IN | ~n29304;
  assign n29268 = ~n29305 | ~P3_ADDRESS_REG_28__SCAN_IN;
  assign U356 = ~n29269 | ~n29268;
  assign n29271 = ~P2_ADDRESS_REG_27__SCAN_IN | ~n29304;
  assign n29270 = ~n29305 | ~P3_ADDRESS_REG_27__SCAN_IN;
  assign U357 = ~n29271 | ~n29270;
  assign n29273 = ~P2_ADDRESS_REG_26__SCAN_IN | ~n29304;
  assign n29272 = ~n29305 | ~P3_ADDRESS_REG_26__SCAN_IN;
  assign U358 = ~n29273 | ~n29272;
  assign n29275 = ~P2_ADDRESS_REG_7__SCAN_IN | ~n29304;
  assign n29274 = ~n29305 | ~P3_ADDRESS_REG_7__SCAN_IN;
  assign U349 = ~n29275 | ~n29274;
  assign n29277 = ~P2_ADDRESS_REG_24__SCAN_IN | ~n29304;
  assign n29276 = ~n29305 | ~P3_ADDRESS_REG_24__SCAN_IN;
  assign U360 = ~n29277 | ~n29276;
  assign n29279 = ~P2_ADDRESS_REG_23__SCAN_IN | ~n29304;
  assign n29278 = ~n29305 | ~P3_ADDRESS_REG_23__SCAN_IN;
  assign U361 = ~n29279 | ~n29278;
  assign n29281 = ~P2_ADDRESS_REG_6__SCAN_IN | ~n29304;
  assign n29280 = ~n29305 | ~P3_ADDRESS_REG_6__SCAN_IN;
  assign U350 = ~n29281 | ~n29280;
  assign n29283 = ~P2_ADDRESS_REG_5__SCAN_IN | ~n29304;
  assign n29282 = ~n29305 | ~P3_ADDRESS_REG_5__SCAN_IN;
  assign U351 = ~n29283 | ~n29282;
  assign n29285 = ~P2_ADDRESS_REG_4__SCAN_IN | ~n29304;
  assign n29284 = ~n29305 | ~P3_ADDRESS_REG_4__SCAN_IN;
  assign U352 = ~n29285 | ~n29284;
  assign n29287 = ~P2_ADDRESS_REG_3__SCAN_IN | ~n29304;
  assign n29286 = ~n29305 | ~P3_ADDRESS_REG_3__SCAN_IN;
  assign U353 = ~n29287 | ~n29286;
  assign n29289 = ~P2_ADDRESS_REG_2__SCAN_IN | ~n29304;
  assign n29288 = ~n29305 | ~P3_ADDRESS_REG_2__SCAN_IN;
  assign U354 = ~n29289 | ~n29288;
  assign n29291 = ~P2_ADDRESS_REG_1__SCAN_IN | ~n29304;
  assign n29290 = ~n29305 | ~P3_ADDRESS_REG_1__SCAN_IN;
  assign U365 = ~n29291 | ~n29290;
  assign n29293 = ~P2_ADDRESS_REG_16__SCAN_IN | ~n29304;
  assign n29292 = ~n29305 | ~P3_ADDRESS_REG_16__SCAN_IN;
  assign U369 = ~n29293 | ~n29292;
  assign n29295 = ~P2_ADDRESS_REG_15__SCAN_IN | ~n29304;
  assign n29294 = ~n29305 | ~P3_ADDRESS_REG_15__SCAN_IN;
  assign U370 = ~n29295 | ~n29294;
  assign n29297 = ~P2_ADDRESS_REG_29__SCAN_IN | ~n29304;
  assign n29296 = ~n29305 | ~P3_ADDRESS_REG_29__SCAN_IN;
  assign U355 = ~n29297 | ~n29296;
  assign n29299 = ~P2_ADDRESS_REG_14__SCAN_IN | ~n29304;
  assign n29298 = ~n29305 | ~P3_ADDRESS_REG_14__SCAN_IN;
  assign U371 = ~n29299 | ~n29298;
  assign n29301 = ~P2_ADDRESS_REG_13__SCAN_IN | ~n29304;
  assign n29300 = ~n29305 | ~P3_ADDRESS_REG_13__SCAN_IN;
  assign U372 = ~n29301 | ~n29300;
  assign n29303 = ~P2_ADDRESS_REG_12__SCAN_IN | ~n29304;
  assign n29302 = ~n29305 | ~P3_ADDRESS_REG_12__SCAN_IN;
  assign U373 = ~n29303 | ~n29302;
  assign n29307 = ~P2_ADDRESS_REG_0__SCAN_IN | ~n29304;
  assign n29306 = ~n29305 | ~P3_ADDRESS_REG_0__SCAN_IN;
  assign U376 = ~n29307 | ~n29306;
  assign n29313 = ~P3_REIP_REG_25__SCAN_IN;
  assign n29434 = ~n29308 | ~P3_STATE_REG_2__SCAN_IN;
  assign n29310 = ~n29313 & ~n29434;
  assign n40723 = ~P3_REIP_REG_26__SCAN_IN;
  assign n29309 = ~n29436 & ~n40723;
  assign n29312 = ~n29310 & ~n29309;
  assign n29311 = ~P3_ADDRESS_REG_24__SCAN_IN | ~n29439;
  assign P3_U3056 = ~n29312 | ~n29311;
  assign n33900 = ~P3_REIP_REG_24__SCAN_IN;
  assign n29315 = ~n33900 & ~n29434;
  assign n29314 = ~n29436 & ~n29313;
  assign n29317 = ~n29315 & ~n29314;
  assign n29316 = ~P3_ADDRESS_REG_23__SCAN_IN | ~n29439;
  assign P3_U3055 = ~n29317 | ~n29316;
  assign n37757 = ~P3_REIP_REG_23__SCAN_IN;
  assign n29319 = ~n37757 & ~n29434;
  assign n29318 = ~n29436 & ~n33900;
  assign n29321 = ~n29319 & ~n29318;
  assign n29320 = ~P3_ADDRESS_REG_22__SCAN_IN | ~n29439;
  assign P3_U3054 = ~n29321 | ~n29320;
  assign n29326 = ~P3_REIP_REG_22__SCAN_IN;
  assign n29323 = ~n29326 & ~n29434;
  assign n29322 = ~n29436 & ~n37757;
  assign n29325 = ~n29323 & ~n29322;
  assign n29324 = ~P3_ADDRESS_REG_21__SCAN_IN | ~n29439;
  assign P3_U3053 = ~n29325 | ~n29324;
  assign n33821 = ~P3_REIP_REG_21__SCAN_IN;
  assign n29328 = ~n33821 & ~n29434;
  assign n29327 = ~n29436 & ~n29326;
  assign n29330 = ~n29328 & ~n29327;
  assign n29329 = ~P3_ADDRESS_REG_20__SCAN_IN | ~n29439;
  assign P3_U3052 = ~n29330 | ~n29329;
  assign n29332 = ~n35979 & ~n29434;
  assign n35904 = ~P3_REIP_REG_2__SCAN_IN;
  assign n29331 = ~n29436 & ~n35904;
  assign n29334 = ~n29332 & ~n29331;
  assign n29333 = ~P3_ADDRESS_REG_0__SCAN_IN | ~n29439;
  assign P3_U3032 = ~n29334 | ~n29333;
  assign n29336 = ~n35904 & ~n29434;
  assign n29339 = ~P3_REIP_REG_3__SCAN_IN;
  assign n29335 = ~n29436 & ~n29339;
  assign n29338 = ~n29336 & ~n29335;
  assign n29337 = ~P3_ADDRESS_REG_1__SCAN_IN | ~n29439;
  assign P3_U3033 = ~n29338 | ~n29337;
  assign n29341 = ~n29339 & ~n29434;
  assign n29340 = ~n29436 & ~n36966;
  assign n29343 = ~n29341 & ~n29340;
  assign n29342 = ~P3_ADDRESS_REG_2__SCAN_IN | ~n29439;
  assign P3_U3034 = ~n29343 | ~n29342;
  assign n34547 = ~P3_REIP_REG_17__SCAN_IN;
  assign n29345 = ~n34547 & ~n29434;
  assign n32853 = ~P3_REIP_REG_18__SCAN_IN;
  assign n29344 = ~n29436 & ~n32853;
  assign n29347 = ~n29345 & ~n29344;
  assign n29346 = ~P3_ADDRESS_REG_16__SCAN_IN | ~n29439;
  assign P3_U3048 = ~n29347 | ~n29346;
  assign n29352 = ~P3_REIP_REG_16__SCAN_IN;
  assign n29349 = ~n29352 & ~n29434;
  assign n29348 = ~n29436 & ~n34547;
  assign n29351 = ~n29349 & ~n29348;
  assign n29350 = ~P3_ADDRESS_REG_15__SCAN_IN | ~n29439;
  assign P3_U3047 = ~n29351 | ~n29350;
  assign n33662 = ~P3_REIP_REG_15__SCAN_IN;
  assign n29354 = ~n33662 & ~n29434;
  assign n29353 = ~n29436 & ~n29352;
  assign n29356 = ~n29354 & ~n29353;
  assign n29355 = ~P3_ADDRESS_REG_14__SCAN_IN | ~n29439;
  assign P3_U3046 = ~n29356 | ~n29355;
  assign n33646 = ~P3_REIP_REG_14__SCAN_IN;
  assign n29358 = ~n33646 & ~n29434;
  assign n29357 = ~n29436 & ~n33662;
  assign n29360 = ~n29358 & ~n29357;
  assign n29359 = ~P3_ADDRESS_REG_13__SCAN_IN | ~n29439;
  assign P3_U3045 = ~n29360 | ~n29359;
  assign n37088 = ~P3_REIP_REG_13__SCAN_IN;
  assign n29362 = ~n37088 & ~n29434;
  assign n29361 = ~n29436 & ~n33646;
  assign n29364 = ~n29362 & ~n29361;
  assign n29363 = ~P3_ADDRESS_REG_12__SCAN_IN | ~n29439;
  assign P3_U3044 = ~n29364 | ~n29363;
  assign n35542 = ~P3_REIP_REG_27__SCAN_IN;
  assign n29366 = ~n35542 & ~n29434;
  assign n29365 = ~n29436 & ~n35543;
  assign n29368 = ~n29366 & ~n29365;
  assign n29367 = ~P3_ADDRESS_REG_26__SCAN_IN | ~n29439;
  assign P3_U3058 = ~n29368 | ~n29367;
  assign n29370 = ~n40723 & ~n29434;
  assign n29369 = ~n29436 & ~n35542;
  assign n29372 = ~n29370 & ~n29369;
  assign n29371 = ~P3_ADDRESS_REG_25__SCAN_IN | ~n29439;
  assign P3_U3057 = ~n29372 | ~n29371;
  assign n32969 = ~P3_REIP_REG_9__SCAN_IN;
  assign n29374 = ~n32969 & ~n29434;
  assign n33074 = ~P3_REIP_REG_10__SCAN_IN;
  assign n29373 = ~n29436 & ~n33074;
  assign n29376 = ~n29374 & ~n29373;
  assign n29375 = ~P3_ADDRESS_REG_8__SCAN_IN | ~n29439;
  assign P3_U3040 = ~n29376 | ~n29375;
  assign n29378 = ~n29381 & ~n29434;
  assign n29377 = ~n29436 & ~n33821;
  assign n29380 = ~n29378 & ~n29377;
  assign n29379 = ~P3_ADDRESS_REG_19__SCAN_IN | ~n29439;
  assign P3_U3051 = ~n29380 | ~n29379;
  assign n29386 = ~P3_REIP_REG_19__SCAN_IN;
  assign n29383 = ~n29386 & ~n29434;
  assign n29382 = ~n29436 & ~n29381;
  assign n29385 = ~n29383 & ~n29382;
  assign n29384 = ~P3_ADDRESS_REG_18__SCAN_IN | ~n29439;
  assign P3_U3050 = ~n29385 | ~n29384;
  assign n29388 = ~n32853 & ~n29434;
  assign n29387 = ~n29436 & ~n29386;
  assign n29390 = ~n29388 & ~n29387;
  assign n29389 = ~P3_ADDRESS_REG_17__SCAN_IN | ~n29439;
  assign P3_U3049 = ~n29390 | ~n29389;
  assign n29403 = ~P3_REIP_REG_30__SCAN_IN;
  assign n29392 = ~n29403 & ~n29434;
  assign n36159 = ~P3_REIP_REG_31__SCAN_IN;
  assign n29391 = ~n29436 & ~n36159;
  assign n29394 = ~n29392 & ~n29391;
  assign n29393 = ~P3_ADDRESS_REG_29__SCAN_IN | ~n29439;
  assign P3_U3061 = ~n29394 | ~n29393;
  assign n29396 = ~n36966 & ~n29434;
  assign n29412 = ~P3_REIP_REG_5__SCAN_IN;
  assign n29395 = ~n29436 & ~n29412;
  assign n29398 = ~n29396 & ~n29395;
  assign n29397 = ~P3_ADDRESS_REG_3__SCAN_IN | ~n29439;
  assign P3_U3035 = ~n29398 | ~n29397;
  assign n29400 = ~n35543 & ~n29434;
  assign n35645 = ~P3_REIP_REG_29__SCAN_IN;
  assign n29399 = ~n29436 & ~n35645;
  assign n29402 = ~n29400 & ~n29399;
  assign n29401 = ~P3_ADDRESS_REG_27__SCAN_IN | ~n29439;
  assign P3_U3059 = ~n29402 | ~n29401;
  assign n29405 = ~n35645 & ~n29434;
  assign n29404 = ~n29436 & ~n29403;
  assign n29407 = ~n29405 & ~n29404;
  assign n29406 = ~P3_ADDRESS_REG_28__SCAN_IN | ~n29439;
  assign P3_U3060 = ~n29407 | ~n29406;
  assign n32968 = ~P3_REIP_REG_8__SCAN_IN;
  assign n29409 = ~n32968 & ~n29434;
  assign n29408 = ~n29436 & ~n32969;
  assign n29411 = ~n29409 & ~n29408;
  assign n29410 = ~P3_ADDRESS_REG_7__SCAN_IN | ~n29439;
  assign P3_U3039 = ~n29411 | ~n29410;
  assign n29414 = ~n29412 & ~n29434;
  assign n33757 = ~P3_REIP_REG_6__SCAN_IN;
  assign n29413 = ~n29436 & ~n33757;
  assign n29416 = ~n29414 & ~n29413;
  assign n29415 = ~P3_ADDRESS_REG_4__SCAN_IN | ~n29439;
  assign P3_U3036 = ~n29416 | ~n29415;
  assign n29418 = ~n33757 & ~n29434;
  assign n33515 = ~P3_REIP_REG_7__SCAN_IN;
  assign n29417 = ~n29436 & ~n33515;
  assign n29420 = ~n29418 & ~n29417;
  assign n29419 = ~P3_ADDRESS_REG_5__SCAN_IN | ~n29439;
  assign P3_U3037 = ~n29420 | ~n29419;
  assign n29425 = ~P3_REIP_REG_11__SCAN_IN;
  assign n29422 = ~n29425 & ~n29434;
  assign n29435 = ~P3_REIP_REG_12__SCAN_IN;
  assign n29421 = ~n29436 & ~n29435;
  assign n29424 = ~n29422 & ~n29421;
  assign n29423 = ~P3_ADDRESS_REG_10__SCAN_IN | ~n29439;
  assign P3_U3042 = ~n29424 | ~n29423;
  assign n29427 = ~n33074 & ~n29434;
  assign n29426 = ~n29436 & ~n29425;
  assign n29429 = ~n29427 & ~n29426;
  assign n29428 = ~P3_ADDRESS_REG_9__SCAN_IN | ~n29439;
  assign P3_U3041 = ~n29429 | ~n29428;
  assign n29431 = ~n33515 & ~n29434;
  assign n29430 = ~n29436 & ~n32968;
  assign n29433 = ~n29431 & ~n29430;
  assign n29432 = ~P3_ADDRESS_REG_6__SCAN_IN | ~n29439;
  assign P3_U3038 = ~n29433 | ~n29432;
  assign n29438 = ~n29435 & ~n29434;
  assign n29437 = ~n29436 & ~n37088;
  assign n29441 = ~n29438 & ~n29437;
  assign n29440 = ~P3_ADDRESS_REG_11__SCAN_IN | ~n29439;
  assign P3_U3043 = ~n29441 | ~n29440;
  assign n29443 = ~n33502;
  assign n29444 = ~n29443 & ~n29442;
  assign n29690 = ~n29444 & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n29445 = ~P3_FLUSH_REG_SCAN_IN;
  assign n29446 = ~n29690 | ~n29445;
  assign n29448 = ~n29446 | ~n41672;
  assign n32362 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n29447 = ~n42012 | ~n31507;
  assign n30030 = ~n41671 | ~n29841;
  assign n43994 = ~n29448 | ~n30030;
  assign P3_U2867 = ~n29449 & ~n43994;
  assign n29451 = ~n29721 | ~P1_BE_N_REG_2__SCAN_IN;
  assign n29450 = ~n29580 | ~P1_BYTEENABLE_REG_2__SCAN_IN;
  assign P1_U3459 = ~n29451 | ~n29450;
  assign n29453 = ~n29721 | ~P1_BE_N_REG_3__SCAN_IN;
  assign n29452 = ~n29580 | ~P1_BYTEENABLE_REG_3__SCAN_IN;
  assign P1_U3458 = ~n29453 | ~n29452;
  assign n29455 = ~n29721 | ~P1_M_IO_N_REG_SCAN_IN;
  assign n29454 = ~n29580 | ~P1_MEMORYFETCH_REG_SCAN_IN;
  assign P1_U3486 = ~n29455 | ~n29454;
  assign n29457 = ~n29721 | ~P1_BE_N_REG_1__SCAN_IN;
  assign n29456 = ~n29580 | ~P1_BYTEENABLE_REG_1__SCAN_IN;
  assign P1_U3460 = ~n29457 | ~n29456;
  assign n29459 = ~n29721 | ~P1_BE_N_REG_0__SCAN_IN;
  assign n29458 = ~n29580 | ~P1_BYTEENABLE_REG_0__SCAN_IN;
  assign P1_U3461 = ~n29459 | ~n29458;
  assign n29460 = ~n29721 | ~P1_ADS_N_REG_SCAN_IN;
  assign P1_U2802 = ~n29461 | ~n29460;
  assign n29464 = ~n29471 & ~n29226;
  assign n29463 = ~n28249 & ~n29549;
  assign n29466 = ~n29464 & ~n29463;
  assign n29465 = ~P2_ADDRESS_REG_13__SCAN_IN | ~n29553;
  assign P2_U3225 = ~n29466 | ~n29465;
  assign n29468 = ~n29506 & ~n29226;
  assign n29467 = ~n28262 & ~n29549;
  assign n29470 = ~n29468 & ~n29467;
  assign n29469 = ~P2_ADDRESS_REG_15__SCAN_IN | ~n29553;
  assign P2_U3227 = ~n29470 | ~n29469;
  assign n29473 = ~n28262 & ~n29226;
  assign n29472 = ~n29471 & ~n29549;
  assign n29475 = ~n29473 & ~n29472;
  assign n29474 = ~P2_ADDRESS_REG_14__SCAN_IN | ~n29553;
  assign P2_U3226 = ~n29475 | ~n29474;
  assign n29477 = ~n28289 & ~n29226;
  assign n29476 = ~n29493 & ~n29549;
  assign n29479 = ~n29477 & ~n29476;
  assign n29478 = ~P2_ADDRESS_REG_18__SCAN_IN | ~n29553;
  assign P2_U3230 = ~n29479 | ~n29478;
  assign n29481 = ~n28345 & ~n29226;
  assign n29480 = ~n29525 & ~n29549;
  assign n29483 = ~n29481 & ~n29480;
  assign n29482 = ~P2_ADDRESS_REG_26__SCAN_IN | ~n29553;
  assign P2_U3238 = ~n29483 | ~n29482;
  assign n29486 = ~n29484 & ~n29226;
  assign n29485 = ~n28354 & ~n29549;
  assign n29488 = ~n29486 & ~n29485;
  assign n29487 = ~P2_ADDRESS_REG_28__SCAN_IN | ~n29553;
  assign P2_U3240 = ~n29488 | ~n29487;
  assign n29490 = ~n28331 & ~n29226;
  assign n29489 = ~n28324 & ~n29549;
  assign n29492 = ~n29490 & ~n29489;
  assign n29491 = ~P2_ADDRESS_REG_24__SCAN_IN | ~n29553;
  assign P2_U3236 = ~n29492 | ~n29491;
  assign n29495 = ~n29493 & ~n29226;
  assign n29494 = ~n36380 & ~n29549;
  assign n29497 = ~n29495 & ~n29494;
  assign n29496 = ~P2_ADDRESS_REG_17__SCAN_IN | ~n29553;
  assign P2_U3229 = ~n29497 | ~n29496;
  assign n29499 = ~n29511 & ~n29226;
  assign n29498 = ~n28289 & ~n29549;
  assign n29501 = ~n29499 & ~n29498;
  assign n29500 = ~P2_ADDRESS_REG_19__SCAN_IN | ~n29553;
  assign P2_U3231 = ~n29501 | ~n29500;
  assign n29503 = ~n29520 & ~n29226;
  assign n29502 = ~n28302 & ~n29549;
  assign n29505 = ~n29503 & ~n29502;
  assign n29504 = ~P2_ADDRESS_REG_21__SCAN_IN | ~n29553;
  assign P2_U3233 = ~n29505 | ~n29504;
  assign n29508 = ~n36380 & ~n29226;
  assign n29507 = ~n29506 & ~n29549;
  assign n29510 = ~n29508 & ~n29507;
  assign n29509 = ~P2_ADDRESS_REG_16__SCAN_IN | ~n29553;
  assign P2_U3228 = ~n29510 | ~n29509;
  assign n29513 = ~n28302 & ~n29226;
  assign n29512 = ~n29511 & ~n29549;
  assign n29515 = ~n29513 & ~n29512;
  assign n29514 = ~P2_ADDRESS_REG_20__SCAN_IN | ~n29553;
  assign P2_U3232 = ~n29515 | ~n29514;
  assign n29517 = ~n28324 & ~n29226;
  assign n29516 = ~n28316 & ~n29549;
  assign n29519 = ~n29517 & ~n29516;
  assign n29518 = ~P2_ADDRESS_REG_23__SCAN_IN | ~n29553;
  assign P2_U3235 = ~n29519 | ~n29518;
  assign n29522 = ~n28316 & ~n29226;
  assign n29521 = ~n29520 & ~n29549;
  assign n29524 = ~n29522 & ~n29521;
  assign n29523 = ~P2_ADDRESS_REG_22__SCAN_IN | ~n29553;
  assign P2_U3234 = ~n29524 | ~n29523;
  assign n29527 = ~n29525 & ~n29226;
  assign n29526 = ~n28331 & ~n29549;
  assign n29529 = ~n29527 & ~n29526;
  assign n29528 = ~P2_ADDRESS_REG_25__SCAN_IN | ~n29553;
  assign P2_U3237 = ~n29529 | ~n29528;
  assign n29531 = ~n28354 & ~n29226;
  assign n29530 = ~n28345 & ~n29549;
  assign n29533 = ~n29531 & ~n29530;
  assign n29532 = ~P2_ADDRESS_REG_27__SCAN_IN | ~n29553;
  assign P2_U3239 = ~n29533 | ~n29532;
  assign n29535 = ~n38814 & ~n29226;
  assign n29534 = ~n23636 & ~n29549;
  assign n29537 = ~n29535 & ~n29534;
  assign n29536 = ~P2_ADDRESS_REG_1__SCAN_IN | ~n29553;
  assign P2_U3213 = ~n29537 | ~n29536;
  assign n29539 = ~P1_REQUESTPENDING_REG_SCAN_IN | ~n29538;
  assign n29548 = ~n29539 | ~n29721;
  assign n29540 = n29541 | P1_STATE_REG_2__SCAN_IN;
  assign n29542 = ~n29540 | ~n29752;
  assign n29753 = ~n29541 & ~HOLD;
  assign n29546 = ~n29542 & ~n29753;
  assign n29718 = ~n29580 | ~P1_STATE_REG_2__SCAN_IN;
  assign n29543 = ~n29579 & ~P1_STATE_REG_0__SCAN_IN;
  assign n29544 = ~n29543 | ~n29749;
  assign n29754 = ~n29718 | ~n29544;
  assign n29545 = ~P1_STATE_REG_0__SCAN_IN & ~n29754;
  assign n29547 = ~n29546 & ~n29545;
  assign P1_U3194 = ~n29548 | ~n29547;
  assign n29552 = ~n29550 & ~n29549;
  assign n29551 = ~n23636 & ~n29226;
  assign n29555 = ~n29552 & ~n29551;
  assign n29554 = ~P2_ADDRESS_REG_0__SCAN_IN | ~n29553;
  assign P2_U3212 = ~n29555 | ~n29554;
  assign n29564 = ~n29556 & ~n32867;
  assign n29559 = ~n29558 | ~n29557;
  assign n29562 = ~n29560 & ~n29559;
  assign n29563 = ~n29562 | ~n29561;
  assign P3_U3030 = ~n29564 | ~n29563;
  assign n34518 = ~n33714 & ~n44100;
  assign n29565 = ~n33710 & ~P1_STATE2_REG_2__SCAN_IN;
  assign n29567 = n34518 & n29565;
  assign n29566 = ~n34550;
  assign n34512 = ~n29566 | ~n33710;
  assign n44093 = ~n34512;
  assign n29571 = ~n29567 & ~n44093;
  assign n29570 = ~n29569 & ~n29568;
  assign P1_U3163 = ~n29571 | ~n29570;
  assign n29573 = ~n29721 | ~P1_W_R_N_REG_SCAN_IN;
  assign n29572 = n29721 | P1_READREQUEST_REG_SCAN_IN;
  assign P1_U3483 = ~n29573 | ~n29572;
  assign n29576 = ~n29721 & ~P1_CODEFETCH_REG_SCAN_IN;
  assign n29575 = ~n29574 & ~P1_STATE_REG_0__SCAN_IN;
  assign n29578 = ~n29576 & ~n29575;
  assign n29577 = ~n29721 | ~P1_D_C_N_REG_SCAN_IN;
  assign P1_U2804 = ~n29578 | ~n29577;
  assign n37228 = ~P1_REIP_REG_10__SCAN_IN;
  assign n29582 = ~n22934 & ~n37228;
  assign n37508 = ~P1_REIP_REG_9__SCAN_IN;
  assign n29581 = ~n37508 & ~n29718;
  assign n29584 = ~n29582 & ~n29581;
  assign n29583 = ~n29721 | ~P1_ADDRESS_REG_8__SCAN_IN;
  assign P1_U3205 = ~n29584 | ~n29583;
  assign n29586 = ~n22934 & ~n42186;
  assign n29627 = ~P1_REIP_REG_21__SCAN_IN;
  assign n29585 = ~n29627 & ~n29718;
  assign n29588 = ~n29586 & ~n29585;
  assign n29587 = ~n29721 | ~P1_ADDRESS_REG_20__SCAN_IN;
  assign P1_U3217 = ~n29588 | ~n29587;
  assign n29679 = ~P1_REIP_REG_14__SCAN_IN;
  assign n29590 = ~n29679 & ~n29718;
  assign n29589 = ~n22934 & ~n40704;
  assign n29592 = ~n29590 & ~n29589;
  assign n29591 = ~n29721 | ~P1_ADDRESS_REG_13__SCAN_IN;
  assign P1_U3210 = ~n29592 | ~n29591;
  assign n29622 = ~P1_REIP_REG_23__SCAN_IN;
  assign n29594 = ~n29622 & ~n29718;
  assign n29593 = ~n22934 & ~n29684;
  assign n29596 = ~n29594 & ~n29593;
  assign n29595 = ~n29721 | ~P1_ADDRESS_REG_22__SCAN_IN;
  assign P1_U3219 = ~n29596 | ~n29595;
  assign n29598 = ~n42488 & ~n29718;
  assign n29597 = ~n22934 & ~n43564;
  assign n29600 = ~n29598 & ~n29597;
  assign n29599 = ~n29721 | ~P1_ADDRESS_REG_27__SCAN_IN;
  assign P1_U3224 = ~n29600 | ~n29599;
  assign n43032 = ~P1_REIP_REG_25__SCAN_IN;
  assign n29602 = ~n43032 & ~n29718;
  assign n29601 = ~n22934 & ~n29632;
  assign n29604 = ~n29602 & ~n29601;
  assign n29603 = ~n29721 | ~P1_ADDRESS_REG_24__SCAN_IN;
  assign P1_U3221 = ~n29604 | ~n29603;
  assign n29656 = ~P1_REIP_REG_16__SCAN_IN;
  assign n29606 = ~n29656 & ~n29718;
  assign n29605 = ~n22934 & ~n29613;
  assign n29608 = ~n29606 & ~n29605;
  assign n29607 = ~n29721 | ~P1_ADDRESS_REG_15__SCAN_IN;
  assign P1_U3212 = ~n29608 | ~n29607;
  assign n38791 = ~P1_REIP_REG_11__SCAN_IN;
  assign n29610 = ~n38791 & ~n29718;
  assign n29651 = ~P1_REIP_REG_12__SCAN_IN;
  assign n29609 = ~n22934 & ~n29651;
  assign n29612 = ~n29610 & ~n29609;
  assign n29611 = ~n29721 | ~P1_ADDRESS_REG_10__SCAN_IN;
  assign P1_U3207 = ~n29612 | ~n29611;
  assign n29615 = ~n29613 & ~n29718;
  assign n29645 = ~P1_REIP_REG_18__SCAN_IN;
  assign n29614 = ~n22934 & ~n29645;
  assign n29617 = ~n29615 & ~n29614;
  assign n29616 = ~n29721 | ~P1_ADDRESS_REG_16__SCAN_IN;
  assign P1_U3213 = ~n29617 | ~n29616;
  assign n29619 = ~n29646 & ~n29718;
  assign n29618 = ~n22934 & ~n41896;
  assign n29621 = ~n29619 & ~n29618;
  assign n29620 = ~n29721 | ~P1_ADDRESS_REG_18__SCAN_IN;
  assign P1_U3215 = ~n29621 | ~n29620;
  assign n29624 = ~n42186 & ~n29718;
  assign n29623 = ~n22934 & ~n29622;
  assign n29626 = ~n29624 & ~n29623;
  assign n29625 = ~n29721 | ~P1_ADDRESS_REG_21__SCAN_IN;
  assign P1_U3218 = ~n29626 | ~n29625;
  assign n29629 = ~n41896 & ~n29718;
  assign n29628 = ~n22934 & ~n29627;
  assign n29631 = ~n29629 & ~n29628;
  assign n29630 = ~n29721 | ~P1_ADDRESS_REG_19__SCAN_IN;
  assign P1_U3216 = ~n29631 | ~n29630;
  assign n29634 = ~n29632 & ~n29718;
  assign n29633 = ~n22934 & ~n29674;
  assign n29636 = ~n29634 & ~n29633;
  assign n29635 = ~n29721 | ~P1_ADDRESS_REG_25__SCAN_IN;
  assign P1_U3222 = ~n29636 | ~n29635;
  assign n29638 = ~n37237 & ~n29718;
  assign n29637 = ~n22934 & ~n37508;
  assign n29640 = ~n29638 & ~n29637;
  assign n29639 = ~n29721 | ~P1_ADDRESS_REG_7__SCAN_IN;
  assign P1_U3204 = ~n29640 | ~n29639;
  assign n29642 = ~n43564 & ~n29718;
  assign n43565 = ~P1_REIP_REG_30__SCAN_IN;
  assign n29641 = ~n22934 & ~n43565;
  assign n29644 = ~n29642 & ~n29641;
  assign n29643 = ~n29721 | ~P1_ADDRESS_REG_28__SCAN_IN;
  assign P1_U3225 = ~n29644 | ~n29643;
  assign n29648 = ~n29645 & ~n29718;
  assign n29647 = ~n22934 & ~n29646;
  assign n29650 = ~n29648 & ~n29647;
  assign n29649 = ~n29721 | ~P1_ADDRESS_REG_17__SCAN_IN;
  assign P1_U3214 = ~n29650 | ~n29649;
  assign n29653 = ~n29651 & ~n29718;
  assign n29652 = ~n22934 & ~n40089;
  assign n29655 = ~n29653 & ~n29652;
  assign n29654 = ~n29721 | ~P1_ADDRESS_REG_11__SCAN_IN;
  assign P1_U3208 = ~n29655 | ~n29654;
  assign n29658 = ~n40704 & ~n29718;
  assign n29657 = ~n22934 & ~n29656;
  assign n29660 = ~n29658 & ~n29657;
  assign n29659 = ~n29721 | ~P1_ADDRESS_REG_14__SCAN_IN;
  assign P1_U3211 = ~n29660 | ~n29659;
  assign n29662 = ~n37228 & ~n29718;
  assign n29661 = ~n22934 & ~n38791;
  assign n29664 = ~n29662 & ~n29661;
  assign n29663 = ~n29721 | ~P1_ADDRESS_REG_9__SCAN_IN;
  assign P1_U3206 = ~n29664 | ~n29663;
  assign n36991 = ~P1_REIP_REG_7__SCAN_IN;
  assign n29666 = ~n36991 & ~n29718;
  assign n29665 = ~n22934 & ~n37237;
  assign n29668 = ~n29666 & ~n29665;
  assign n29667 = ~n29721 | ~P1_ADDRESS_REG_6__SCAN_IN;
  assign P1_U3203 = ~n29668 | ~n29667;
  assign n29671 = ~n43565 & ~n29718;
  assign n29670 = ~n22934 & ~n29669;
  assign n29673 = ~n29671 & ~n29670;
  assign n29672 = ~n29721 | ~P1_ADDRESS_REG_29__SCAN_IN;
  assign P1_U3226 = ~n29673 | ~n29672;
  assign n29676 = ~n29674 & ~n29718;
  assign n29675 = ~n22934 & ~n42488;
  assign n29678 = ~n29676 & ~n29675;
  assign n29677 = ~n29721 | ~P1_ADDRESS_REG_26__SCAN_IN;
  assign P1_U3223 = ~n29678 | ~n29677;
  assign n29681 = ~n40089 & ~n29718;
  assign n29680 = ~n22934 & ~n29679;
  assign n29683 = ~n29681 & ~n29680;
  assign n29682 = ~n29721 | ~P1_ADDRESS_REG_12__SCAN_IN;
  assign P1_U3209 = ~n29683 | ~n29682;
  assign n29686 = ~n29684 & ~n29718;
  assign n29685 = ~n22934 & ~n43032;
  assign n29688 = ~n29686 & ~n29685;
  assign n29687 = ~n29721 | ~P1_ADDRESS_REG_23__SCAN_IN;
  assign P1_U3220 = ~n29688 | ~n29687;
  assign n36057 = ~P3_STATE2_REG_1__SCAN_IN & ~P3_STATE2_REG_3__SCAN_IN;
  assign n35442 = ~n29726 & ~n36057;
  assign n29689 = ~n35442 | ~n43994;
  assign n29695 = ~n29689 | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n29691 = ~P3_FLUSH_REG_SCAN_IN & ~n29690;
  assign n42018 = ~n29691 & ~n31507;
  assign n29692 = ~n42018;
  assign n30873 = ~P3_STATE2_REG_3__SCAN_IN | ~n29997;
  assign n29693 = ~n29692 | ~n30873;
  assign n29694 = ~n29693 | ~n43994;
  assign P3_U2863 = ~n29695 | ~n29694;
  assign n29713 = ~P1_REIP_REG_2__SCAN_IN;
  assign n29697 = ~n29713 & ~n22934;
  assign n29696 = ~n35494 & ~n29718;
  assign n29699 = ~n29697 & ~n29696;
  assign n29698 = ~n29721 | ~P1_ADDRESS_REG_0__SCAN_IN;
  assign P1_U3197 = ~n29699 | ~n29698;
  assign n36103 = ~P1_REIP_REG_5__SCAN_IN;
  assign n29701 = ~n36103 & ~n29718;
  assign n34830 = ~P1_REIP_REG_6__SCAN_IN;
  assign n29700 = ~n34830 & ~n22934;
  assign n29703 = ~n29701 & ~n29700;
  assign n29702 = ~n29721 | ~P1_ADDRESS_REG_4__SCAN_IN;
  assign P1_U3201 = ~n29703 | ~n29702;
  assign n29705 = ~n35875 & ~n29718;
  assign n29708 = ~P1_REIP_REG_4__SCAN_IN;
  assign n29704 = ~n29708 & ~n22934;
  assign n29707 = ~n29705 & ~n29704;
  assign n29706 = ~n29721 | ~P1_ADDRESS_REG_2__SCAN_IN;
  assign P1_U3199 = ~n29707 | ~n29706;
  assign n29710 = ~n29708 & ~n29718;
  assign n29709 = ~n36103 & ~n22934;
  assign n29712 = ~n29710 & ~n29709;
  assign n29711 = ~n29721 | ~P1_ADDRESS_REG_3__SCAN_IN;
  assign P1_U3200 = ~n29712 | ~n29711;
  assign n29715 = ~n29713 & ~n29718;
  assign n29714 = ~n35875 & ~n22934;
  assign n29717 = ~n29715 & ~n29714;
  assign n29716 = ~n29721 | ~P1_ADDRESS_REG_1__SCAN_IN;
  assign P1_U3198 = ~n29717 | ~n29716;
  assign n29720 = ~n34830 & ~n29718;
  assign n29719 = ~n36991 & ~n22934;
  assign n29723 = ~n29720 & ~n29719;
  assign n29722 = ~n29721 | ~P1_ADDRESS_REG_5__SCAN_IN;
  assign P1_U3202 = ~n29723 | ~n29722;
  assign n29995 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n30048 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~n29995;
  assign n29870 = ~n30048;
  assign n29724 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n29995;
  assign n29725 = ~n29870 | ~n29724;
  assign n31370 = ~n29726;
  assign n29843 = ~P3_STATEBS16_REG_SCAN_IN & ~n31370;
  assign n29738 = n36057 | n29843;
  assign n29731 = ~n29725 | ~n29738;
  assign n30560 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n29844 = ~n30560;
  assign n30870 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n29727 = ~n29844 | ~n30870;
  assign n29729 = ~n43990 & ~n29727;
  assign n30777 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n30048;
  assign n29728 = ~n43992 & ~n30777;
  assign n29730 = ~n29729 & ~n29728;
  assign n29732 = ~n29731 | ~n29730;
  assign n29737 = ~n29732 | ~n43994;
  assign n29734 = ~P3_STATE2_REG_3__SCAN_IN | ~n41354;
  assign n41344 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n30559 = P3_STATE2_REG_3__SCAN_IN & n41344;
  assign n29733 = ~n43994;
  assign n29740 = ~n30559 & ~n29733;
  assign n29735 = ~n29734 | ~n29740;
  assign n29736 = ~n29735 | ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign P3_U2866 = ~n29737 | ~n29736;
  assign n43989 = ~n43994 | ~n29738;
  assign n29996 = ~n41354 | ~n41341;
  assign n29739 = ~n29995 | ~n29996;
  assign n29742 = ~n43989 & ~n29739;
  assign n29741 = ~n29740 & ~n41354;
  assign n29748 = ~n29742 & ~n29741;
  assign n29744 = ~n43990;
  assign n29743 = ~n41344 & ~n43992;
  assign n29745 = ~n29744 & ~n29743;
  assign n29746 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~n29745;
  assign n29747 = ~n29746 | ~n43994;
  assign P3_U2865 = ~n29748 | ~n29747;
  assign n29758 = ~n29749 | ~n44100;
  assign n29751 = ~n29758 & ~n29750;
  assign n29757 = ~n29751 | ~P1_STATE_REG_1__SCAN_IN;
  assign n29755 = ~n29753 & ~n29752;
  assign n29756 = ~n29755 & ~n29754;
  assign n29765 = n29757 & n29756;
  assign n29759 = n29758 & P1_STATE_REG_1__SCAN_IN;
  assign n29760 = ~n29759 & ~P1_REQUESTPENDING_REG_SCAN_IN;
  assign n29762 = ~P1_STATE_REG_2__SCAN_IN & ~n29760;
  assign n29763 = ~n29762 & ~n29761;
  assign n29764 = ~P1_STATE_REG_0__SCAN_IN | ~n29763;
  assign P1_U3196 = ~n29765 | ~n29764;
  assign n29772 = ~n29835 & ~P3_BE_N_REG_3__SCAN_IN;
  assign n29769 = ~P3_D_C_N_REG_SCAN_IN & ~P3_W_R_N_REG_SCAN_IN;
  assign n29766 = ~P3_BE_N_REG_0__SCAN_IN & ~P3_BE_N_REG_1__SCAN_IN;
  assign n29767 = ~P3_M_IO_N_REG_SCAN_IN | ~n29766;
  assign n29768 = ~n29767 & ~P3_ADS_N_REG_SCAN_IN;
  assign n29770 = ~n29769 | ~n29768;
  assign n29771 = ~n29770 & ~P3_BE_N_REG_2__SCAN_IN;
  assign U213 = ~n29772 | ~n29771;
  assign n29774 = ~BUF2_REG_12__SCAN_IN | ~U215;
  assign n29773 = ~P2_DATAO_REG_12__SCAN_IN | ~n29835;
  assign U263 = ~n29774 | ~n29773;
  assign n29776 = ~BUF2_REG_10__SCAN_IN | ~U215;
  assign n29775 = ~P2_DATAO_REG_10__SCAN_IN | ~n29835;
  assign U261 = ~n29776 | ~n29775;
  assign n29778 = ~BUF2_REG_13__SCAN_IN | ~U215;
  assign n29777 = ~P2_DATAO_REG_13__SCAN_IN | ~n29835;
  assign U264 = ~n29778 | ~n29777;
  assign n29780 = ~BUF2_REG_14__SCAN_IN | ~U215;
  assign n29779 = ~P2_DATAO_REG_14__SCAN_IN | ~n29835;
  assign U265 = ~n29780 | ~n29779;
  assign n29782 = ~BUF2_REG_15__SCAN_IN | ~U215;
  assign n29781 = ~P2_DATAO_REG_15__SCAN_IN | ~n29835;
  assign U266 = ~n29782 | ~n29781;
  assign n29784 = ~BUF2_REG_16__SCAN_IN | ~U215;
  assign n29783 = ~P2_DATAO_REG_16__SCAN_IN | ~n29835;
  assign U267 = ~n29784 | ~n29783;
  assign n29786 = ~BUF2_REG_17__SCAN_IN | ~U215;
  assign n29785 = ~P2_DATAO_REG_17__SCAN_IN | ~n29835;
  assign U268 = ~n29786 | ~n29785;
  assign n29788 = ~BUF2_REG_18__SCAN_IN | ~U215;
  assign n29787 = ~P2_DATAO_REG_18__SCAN_IN | ~n29835;
  assign U269 = ~n29788 | ~n29787;
  assign n29790 = ~BUF2_REG_19__SCAN_IN | ~U215;
  assign n29789 = ~P2_DATAO_REG_19__SCAN_IN | ~n29835;
  assign U270 = ~n29790 | ~n29789;
  assign n29792 = ~BUF2_REG_20__SCAN_IN | ~U215;
  assign n29791 = ~P2_DATAO_REG_20__SCAN_IN | ~n29835;
  assign U271 = ~n29792 | ~n29791;
  assign n29794 = ~BUF2_REG_21__SCAN_IN | ~U215;
  assign n29793 = ~P2_DATAO_REG_21__SCAN_IN | ~n29835;
  assign U272 = ~n29794 | ~n29793;
  assign n29796 = ~BUF2_REG_22__SCAN_IN | ~U215;
  assign n29795 = ~P2_DATAO_REG_22__SCAN_IN | ~n29835;
  assign U273 = ~n29796 | ~n29795;
  assign n29798 = ~BUF2_REG_23__SCAN_IN | ~U215;
  assign n29797 = ~P2_DATAO_REG_23__SCAN_IN | ~n29835;
  assign U274 = ~n29798 | ~n29797;
  assign n29800 = ~BUF2_REG_24__SCAN_IN | ~U215;
  assign n29799 = ~P2_DATAO_REG_24__SCAN_IN | ~n29835;
  assign U275 = ~n29800 | ~n29799;
  assign n29802 = ~BUF2_REG_25__SCAN_IN | ~U215;
  assign n29801 = ~P2_DATAO_REG_25__SCAN_IN | ~n29835;
  assign U276 = ~n29802 | ~n29801;
  assign n29804 = ~BUF2_REG_26__SCAN_IN | ~U215;
  assign n29803 = ~P2_DATAO_REG_26__SCAN_IN | ~n29835;
  assign U277 = ~n29804 | ~n29803;
  assign n29806 = ~BUF2_REG_27__SCAN_IN | ~U215;
  assign n29805 = ~P2_DATAO_REG_27__SCAN_IN | ~n29835;
  assign U278 = ~n29806 | ~n29805;
  assign n29808 = ~BUF2_REG_9__SCAN_IN | ~U215;
  assign n29807 = ~P2_DATAO_REG_9__SCAN_IN | ~n29835;
  assign U260 = ~n29808 | ~n29807;
  assign n29810 = ~BUF2_REG_8__SCAN_IN | ~U215;
  assign n29809 = ~P2_DATAO_REG_8__SCAN_IN | ~n29835;
  assign U259 = ~n29810 | ~n29809;
  assign n29812 = ~BUF2_REG_7__SCAN_IN | ~U215;
  assign n29811 = ~P2_DATAO_REG_7__SCAN_IN | ~n29835;
  assign U258 = ~n29812 | ~n29811;
  assign n29814 = ~BUF2_REG_6__SCAN_IN | ~U215;
  assign n29813 = ~P2_DATAO_REG_6__SCAN_IN | ~n29835;
  assign U257 = ~n29814 | ~n29813;
  assign n29816 = ~BUF2_REG_5__SCAN_IN | ~U215;
  assign n29815 = ~P2_DATAO_REG_5__SCAN_IN | ~n29835;
  assign U256 = ~n29816 | ~n29815;
  assign n29818 = ~BUF2_REG_28__SCAN_IN | ~U215;
  assign n29817 = ~P2_DATAO_REG_28__SCAN_IN | ~n29835;
  assign U279 = ~n29818 | ~n29817;
  assign n29820 = ~BUF2_REG_29__SCAN_IN | ~U215;
  assign n29819 = ~P2_DATAO_REG_29__SCAN_IN | ~n29835;
  assign U280 = ~n29820 | ~n29819;
  assign n29822 = ~BUF2_REG_30__SCAN_IN | ~U215;
  assign n29821 = ~P2_DATAO_REG_30__SCAN_IN | ~n29835;
  assign U281 = ~n29822 | ~n29821;
  assign n29824 = ~BUF2_REG_31__SCAN_IN | ~U215;
  assign n29823 = ~P2_DATAO_REG_31__SCAN_IN | ~n29835;
  assign U282 = ~n29824 | ~n29823;
  assign n29826 = ~BUF2_REG_4__SCAN_IN | ~U215;
  assign n29825 = ~P2_DATAO_REG_4__SCAN_IN | ~n29835;
  assign U255 = ~n29826 | ~n29825;
  assign n29828 = ~BUF2_REG_3__SCAN_IN | ~U215;
  assign n29827 = ~P2_DATAO_REG_3__SCAN_IN | ~n29835;
  assign U254 = ~n29828 | ~n29827;
  assign n29830 = ~BUF2_REG_2__SCAN_IN | ~U215;
  assign n29829 = ~P2_DATAO_REG_2__SCAN_IN | ~n29835;
  assign U253 = ~n29830 | ~n29829;
  assign n29832 = ~BUF2_REG_1__SCAN_IN | ~U215;
  assign n29831 = ~P2_DATAO_REG_1__SCAN_IN | ~n29835;
  assign U252 = ~n29832 | ~n29831;
  assign n29834 = ~BUF2_REG_0__SCAN_IN | ~U215;
  assign n29833 = ~P2_DATAO_REG_0__SCAN_IN | ~n29835;
  assign U251 = ~n29834 | ~n29833;
  assign n29837 = ~BUF2_REG_11__SCAN_IN | ~U215;
  assign n29836 = ~P2_DATAO_REG_11__SCAN_IN | ~n29835;
  assign U262 = ~n29837 | ~n29836;
  assign n31014 = ~BUF2_REG_4__SCAN_IN | ~n30874;
  assign n29838 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ n29997;
  assign n29923 = ~n41341 | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n29881 = ~n29997 | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n43993 = n29923 & n29881;
  assign n29884 = ~n29838 | ~n43993;
  assign n29845 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~n29884;
  assign n41382 = ~P3_STATE2_REG_3__SCAN_IN | ~n40527;
  assign n30809 = ~n29845 | ~n41382;
  assign n29840 = ~n31014 & ~n30809;
  assign n30900 = ~n41341 & ~n29844;
  assign n31045 = ~n29997 | ~n30900;
  assign n41095 = ~n43990 & ~n30030;
  assign n31015 = ~BUF2_REG_20__SCAN_IN | ~n41095;
  assign n29839 = ~n31045 & ~n31015;
  assign n29854 = ~n29840 & ~n29839;
  assign n30862 = ~n29923 & ~n29844;
  assign n30812 = ~n30862;
  assign n31018 = ~BUF2_REG_28__SCAN_IN | ~n41095;
  assign n29852 = ~n30812 & ~n31018;
  assign n32374 = ~P3_STATE2_REG_0__SCAN_IN & ~n43992;
  assign n30705 = ~n32374 | ~n29841;
  assign n31019 = ~n31801 & ~n30705;
  assign n41350 = ~n41341 | ~n29997;
  assign n30894 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~n41337;
  assign n30813 = ~n41350 & ~n30894;
  assign n29850 = ~n31019 | ~n30813;
  assign n29842 = ~n30813 & ~n43992;
  assign n29848 = ~n29842 & ~n30030;
  assign n30027 = ~P3_STATE2_REG_2__SCAN_IN & ~n29843;
  assign n30011 = ~n43993 & ~n29844;
  assign n29846 = ~n30027 | ~n30011;
  assign n29857 = ~n29845;
  assign n29847 = ~n29846 | ~n29857;
  assign n30814 = ~n29848 | ~n29847;
  assign n29849 = ~P3_INSTQUEUE_REG_4__4__SCAN_IN | ~n30814;
  assign n29851 = ~n29850 | ~n29849;
  assign n29853 = ~n29852 & ~n29851;
  assign P3_U2904 = ~n29854 | ~n29853;
  assign n29927 = ~n43993 & ~n30894;
  assign n30797 = ~n29927 | ~n41382;
  assign n29856 = ~n31014 & ~n30797;
  assign n30800 = ~n30813;
  assign n29855 = ~n31015 & ~n30800;
  assign n29867 = ~n29856 & ~n29855;
  assign n31040 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n30900;
  assign n29865 = ~n31018 & ~n31040;
  assign n30801 = ~n29881 & ~n30894;
  assign n29863 = ~n31019 | ~n30801;
  assign n30049 = ~n30027;
  assign n29858 = ~n29857 & ~n30049;
  assign n29859 = ~n29858 & ~n29927;
  assign n29861 = ~n29859 & ~n30030;
  assign n30773 = ~n30801;
  assign n29860 = ~P3_STATE2_REG_3__SCAN_IN | ~n30773;
  assign n30802 = ~n29861 | ~n29860;
  assign n29862 = ~P3_INSTQUEUE_REG_6__4__SCAN_IN | ~n30802;
  assign n29864 = ~n29863 | ~n29862;
  assign n29866 = ~n29865 & ~n29864;
  assign P3_U2920 = ~n29867 | ~n29866;
  assign n29897 = ~n41337 & ~n29996;
  assign n30774 = ~n29897 | ~n41382;
  assign n29869 = ~n31014 & ~n30774;
  assign n29868 = ~n31015 & ~n30777;
  assign n29880 = ~n29869 & ~n29868;
  assign n29878 = ~n31018 & ~n30773;
  assign n30750 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n29897;
  assign n30778 = ~n30750;
  assign n29876 = ~n31019 | ~n30778;
  assign n29871 = ~n29870 & ~n30049;
  assign n29872 = ~n29871 & ~n29897;
  assign n29874 = ~n29872 & ~n30030;
  assign n29873 = ~P3_STATE2_REG_3__SCAN_IN | ~n30750;
  assign n30779 = ~n29874 | ~n29873;
  assign n29875 = ~P3_INSTQUEUE_REG_9__4__SCAN_IN | ~n30779;
  assign n29877 = ~n29876 | ~n29875;
  assign n29879 = ~n29878 & ~n29877;
  assign P3_U2944 = ~n29880 | ~n29879;
  assign n30597 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n41354;
  assign n30877 = ~n41341 & ~n30597;
  assign n30993 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n30877;
  assign n29883 = ~n31018 & ~n30993;
  assign n30994 = ~n29923 & ~n30870;
  assign n30836 = ~n30994;
  assign n30789 = ~n29881 & ~n30870;
  assign n30857 = ~n30789;
  assign n30000 = ~n30836 | ~n30857;
  assign n30786 = ~n41382 | ~n30000;
  assign n29882 = ~n31014 & ~n30786;
  assign n29894 = ~n29883 & ~n29882;
  assign n30707 = ~n41350 & ~n30870;
  assign n30832 = ~n30707;
  assign n29892 = ~n31015 & ~n30832;
  assign n29890 = ~n31019 | ~n30789;
  assign n29912 = ~n41337 & ~n29884;
  assign n29885 = ~n30027 | ~n29912;
  assign n29886 = ~n30836 | ~n29885;
  assign n29887 = ~n29886 | ~n43992;
  assign n29888 = ~n29887 | ~n30857;
  assign n30790 = ~n30874 | ~n29888;
  assign n29889 = ~P3_INSTQUEUE_REG_14__4__SCAN_IN | ~n30790;
  assign n29891 = ~n29890 | ~n29889;
  assign n29893 = ~n29892 & ~n29891;
  assign P3_U2984 = ~n29894 | ~n29893;
  assign n29896 = ~n31018 & ~n30777;
  assign n29898 = ~n43993 & ~n30597;
  assign n30761 = ~n29898 | ~n41382;
  assign n29895 = ~n31014 & ~n30761;
  assign n29908 = ~n29896 & ~n29895;
  assign n30764 = ~n29897 | ~n29997;
  assign n29906 = ~n31015 & ~n30764;
  assign n30990 = ~n29997 | ~n30877;
  assign n30765 = ~n30990;
  assign n29904 = ~n31019 | ~n30765;
  assign n29924 = ~n30777 | ~n30764;
  assign n29899 = ~n30027 | ~n29924;
  assign n29911 = ~n29898;
  assign n29902 = ~n29899 | ~n29911;
  assign n29900 = ~n43992 & ~n30765;
  assign n29901 = ~n29900 & ~n30030;
  assign n30766 = ~n29902 | ~n29901;
  assign n29903 = ~P3_INSTQUEUE_REG_10__4__SCAN_IN | ~n30766;
  assign n29905 = ~n29904 | ~n29903;
  assign n29907 = ~n29906 & ~n29905;
  assign P3_U2952 = ~n29908 | ~n29907;
  assign n29910 = ~n31018 & ~n30750;
  assign n30702 = ~n29912 | ~n41382;
  assign n29909 = ~n31014 & ~n30702;
  assign n29922 = ~n29910 & ~n29909;
  assign n29920 = ~n31015 & ~n30990;
  assign n29918 = ~n31019 | ~n30707;
  assign n29915 = ~n30707 & ~n43992;
  assign n29913 = ~n29911 & ~n30049;
  assign n29914 = ~n29913 & ~n29912;
  assign n29916 = ~n29915 & ~n29914;
  assign n30708 = ~n30874 | ~n29916;
  assign n29917 = ~P3_INSTQUEUE_REG_12__4__SCAN_IN | ~n30708;
  assign n29919 = ~n29918 | ~n29917;
  assign n29921 = ~n29920 & ~n29919;
  assign P3_U2968 = ~n29922 | ~n29921;
  assign n31047 = ~n29923 & ~n30894;
  assign n30740 = ~n31047;
  assign n29926 = ~n31018 & ~n30740;
  assign n30737 = ~n41382 | ~n29924;
  assign n29925 = ~n31014 & ~n30737;
  assign n29937 = ~n29926 & ~n29925;
  assign n29935 = ~n31015 & ~n30773;
  assign n30741 = ~n30764;
  assign n29933 = ~n31019 | ~n30741;
  assign n29928 = ~n30027 | ~n29927;
  assign n29929 = ~n30777 | ~n29928;
  assign n29930 = ~n29929 | ~n43992;
  assign n29931 = ~n29930 | ~n30764;
  assign n30742 = ~n30874 | ~n29931;
  assign n29932 = ~P3_INSTQUEUE_REG_8__4__SCAN_IN | ~n30742;
  assign n29934 = ~n29933 | ~n29932;
  assign n29936 = ~n29935 & ~n29934;
  assign P3_U2936 = ~n29937 | ~n29936;
  assign n31003 = ~BUF2_REG_2__SCAN_IN | ~n30874;
  assign n29939 = ~n31003 & ~n30761;
  assign n31006 = ~BUF2_REG_26__SCAN_IN | ~n41095;
  assign n29938 = ~n31006 & ~n30777;
  assign n29946 = ~n29939 & ~n29938;
  assign n31002 = ~BUF2_REG_18__SCAN_IN | ~n41095;
  assign n29944 = ~n31002 & ~n30764;
  assign n31007 = ~n29940 & ~n30705;
  assign n29942 = ~n31007 | ~n30765;
  assign n29941 = ~P3_INSTQUEUE_REG_10__2__SCAN_IN | ~n30766;
  assign n29943 = ~n29942 | ~n29941;
  assign n29945 = ~n29944 & ~n29943;
  assign P3_U2950 = ~n29946 | ~n29945;
  assign n29948 = ~n31002 & ~n30773;
  assign n29947 = ~n31003 & ~n30737;
  assign n29954 = ~n29948 & ~n29947;
  assign n29952 = ~n31006 & ~n30740;
  assign n29950 = ~n31007 | ~n30741;
  assign n29949 = ~P3_INSTQUEUE_REG_8__2__SCAN_IN | ~n30742;
  assign n29951 = ~n29950 | ~n29949;
  assign n29953 = ~n29952 & ~n29951;
  assign P3_U2934 = ~n29954 | ~n29953;
  assign n29956 = ~n31003 & ~n30797;
  assign n29955 = ~n31006 & ~n31040;
  assign n29962 = ~n29956 & ~n29955;
  assign n29960 = ~n31002 & ~n30800;
  assign n29958 = ~n31007 | ~n30801;
  assign n29957 = ~P3_INSTQUEUE_REG_6__2__SCAN_IN | ~n30802;
  assign n29959 = ~n29958 | ~n29957;
  assign n29961 = ~n29960 & ~n29959;
  assign P3_U2918 = ~n29962 | ~n29961;
  assign n29964 = ~n31002 & ~n30832;
  assign n29963 = ~n31003 & ~n30786;
  assign n29970 = ~n29964 & ~n29963;
  assign n29968 = ~n31006 & ~n30993;
  assign n29966 = ~n31007 | ~n30789;
  assign n29965 = ~P3_INSTQUEUE_REG_14__2__SCAN_IN | ~n30790;
  assign n29967 = ~n29966 | ~n29965;
  assign n29969 = ~n29968 & ~n29967;
  assign P3_U2982 = ~n29970 | ~n29969;
  assign n29974 = ~n30702 & ~n31003;
  assign n29972 = ~P3_INSTQUEUE_REG_12__2__SCAN_IN | ~n30708;
  assign n29971 = ~n31007 | ~n30707;
  assign n29973 = ~n29972 | ~n29971;
  assign n29978 = ~n29974 & ~n29973;
  assign n29976 = ~n31002 & ~n30990;
  assign n29975 = ~n31006 & ~n30750;
  assign n29977 = ~n29976 & ~n29975;
  assign P3_U2966 = ~n29978 | ~n29977;
  assign n29982 = ~n30774 & ~n31003;
  assign n29980 = ~P3_INSTQUEUE_REG_9__2__SCAN_IN | ~n30779;
  assign n29979 = ~n31007 | ~n30778;
  assign n29981 = ~n29980 | ~n29979;
  assign n29986 = ~n29982 & ~n29981;
  assign n29984 = ~n31002 & ~n30777;
  assign n29983 = ~n31006 & ~n30773;
  assign n29985 = ~n29984 & ~n29983;
  assign P3_U2942 = ~n29986 | ~n29985;
  assign n29990 = ~n30809 & ~n31003;
  assign n29988 = ~P3_INSTQUEUE_REG_4__2__SCAN_IN | ~n30814;
  assign n29987 = ~n31007 | ~n30813;
  assign n29989 = ~n29988 | ~n29987;
  assign n29994 = ~n29990 & ~n29989;
  assign n29992 = ~n30812 & ~n31006;
  assign n29991 = ~n31045 & ~n31002;
  assign n29993 = ~n29992 & ~n29991;
  assign P3_U2902 = ~n29994 | ~n29993;
  assign n30213 = ~n41337 & ~n29995;
  assign n30861 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n30213;
  assign n30029 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~n29996;
  assign n30848 = ~n30029 | ~n29997;
  assign n30014 = ~n30861 | ~n30848;
  assign n30821 = ~n41382 | ~n30014;
  assign n29999 = ~n31014 & ~n30821;
  assign n29998 = ~n31015 & ~n30857;
  assign n30010 = ~n29999 & ~n29998;
  assign n30008 = ~n31018 & ~n30836;
  assign n30824 = ~n30848;
  assign n30006 = ~n30824 | ~n31019;
  assign n30001 = ~n30027 | ~n30000;
  assign n30002 = ~n30861 | ~n30001;
  assign n30003 = ~n30002 | ~n43992;
  assign n30004 = ~n30003 | ~n30848;
  assign n30825 = ~n30874 | ~n30004;
  assign n30005 = ~P3_INSTQUEUE_REG_0__4__SCAN_IN | ~n30825;
  assign n30007 = ~n30006 | ~n30005;
  assign n30009 = ~n30008 & ~n30007;
  assign P3_U2872 = ~n30010 | ~n30009;
  assign n30845 = ~n30011 | ~n41382;
  assign n30013 = ~n30845 & ~n31014;
  assign n30012 = ~n30861 & ~n31018;
  assign n30024 = ~n30013 & ~n30012;
  assign n30022 = ~n30848 & ~n31015;
  assign n30849 = ~n31045;
  assign n30020 = ~n30849 | ~n31019;
  assign n30015 = ~n30027 | ~n30014;
  assign n30016 = ~n30812 | ~n30015;
  assign n30017 = ~n30016 | ~n43992;
  assign n30018 = ~n30017 | ~n31045;
  assign n30850 = ~n30874 | ~n30018;
  assign n30019 = ~P3_INSTQUEUE_REG_2__4__SCAN_IN | ~n30850;
  assign n30021 = ~n30020 | ~n30019;
  assign n30023 = ~n30022 & ~n30021;
  assign P3_U2888 = ~n30024 | ~n30023;
  assign n30026 = ~n31018 & ~n30857;
  assign n30858 = ~n30029 | ~n41382;
  assign n30025 = ~n31014 & ~n30858;
  assign n30039 = ~n30026 & ~n30025;
  assign n30037 = ~n30861 & ~n31015;
  assign n30035 = ~n30862 | ~n31019;
  assign n30028 = n30213 & n30027;
  assign n30031 = ~n30029 & ~n30028;
  assign n30033 = ~n30031 & ~n30030;
  assign n30032 = ~P3_STATE2_REG_3__SCAN_IN | ~n30812;
  assign n30863 = ~n30033 | ~n30032;
  assign n30034 = ~P3_INSTQUEUE_REG_1__4__SCAN_IN | ~n30863;
  assign n30036 = ~n30035 | ~n30034;
  assign n30038 = ~n30037 & ~n30036;
  assign P3_U2880 = ~n30039 | ~n30038;
  assign n30041 = ~n31003 & ~n30821;
  assign n30040 = ~n31006 & ~n30836;
  assign n30047 = ~n30041 & ~n30040;
  assign n30045 = ~n31002 & ~n30857;
  assign n30043 = ~n30824 | ~n31007;
  assign n30042 = ~P3_INSTQUEUE_REG_0__2__SCAN_IN | ~n30825;
  assign n30044 = ~n30043 | ~n30042;
  assign n30046 = ~n30045 & ~n30044;
  assign P3_U2870 = ~n30047 | ~n30046;
  assign n30726 = ~n30048 | ~n41382;
  assign n30056 = ~n30726 & ~n31014;
  assign n30050 = ~n41341 | ~n30049;
  assign n30558 = ~n30874 | ~n30050;
  assign n30052 = ~n30558 & ~n30894;
  assign n30051 = ~P3_STATE2_REG_3__SCAN_IN | ~n30777;
  assign n30730 = ~n30052 | ~n30051;
  assign n30054 = ~P3_INSTQUEUE_REG_7__4__SCAN_IN | ~n30730;
  assign n30729 = ~n30777;
  assign n30053 = ~n31019 | ~n30729;
  assign n30055 = ~n30054 | ~n30053;
  assign n30060 = ~n30056 & ~n30055;
  assign n30058 = ~n31018 & ~n30800;
  assign n30057 = ~n31015 & ~n30740;
  assign n30059 = ~n30058 & ~n30057;
  assign P3_U2928 = ~n30060 | ~n30059;
  assign n30064 = ~n30726 & ~n31003;
  assign n30062 = ~P3_INSTQUEUE_REG_7__2__SCAN_IN | ~n30730;
  assign n30061 = ~n31007 | ~n30729;
  assign n30063 = ~n30062 | ~n30061;
  assign n30068 = ~n30064 & ~n30063;
  assign n30066 = ~n31002 & ~n30740;
  assign n30065 = ~n31006 & ~n30800;
  assign n30067 = ~n30066 & ~n30065;
  assign P3_U2926 = ~n30068 | ~n30067;
  assign n30070 = ~n30845 & ~n31003;
  assign n30069 = ~n30848 & ~n31002;
  assign n30076 = ~n30070 & ~n30069;
  assign n30074 = ~n30861 & ~n31006;
  assign n30072 = ~n30849 | ~n31007;
  assign n30071 = ~P3_INSTQUEUE_REG_2__2__SCAN_IN | ~n30850;
  assign n30073 = ~n30072 | ~n30071;
  assign n30075 = ~n30074 & ~n30073;
  assign P3_U2886 = ~n30076 | ~n30075;
  assign n30080 = ~n30858 & ~n31003;
  assign n30078 = ~P3_INSTQUEUE_REG_1__2__SCAN_IN | ~n30863;
  assign n30077 = ~n30862 | ~n31007;
  assign n30079 = ~n30078 | ~n30077;
  assign n30084 = ~n30080 & ~n30079;
  assign n30082 = ~n31006 & ~n30857;
  assign n30081 = ~n30861 & ~n31002;
  assign n30083 = ~n30082 & ~n30081;
  assign P3_U2878 = ~n30084 | ~n30083;
  assign n31026 = ~BUF2_REG_3__SCAN_IN | ~n30874;
  assign n30086 = ~n31026 & ~n30797;
  assign n31030 = ~BUF2_REG_27__SCAN_IN | ~n41095;
  assign n30085 = ~n31030 & ~n31040;
  assign n30092 = ~n30086 & ~n30085;
  assign n31027 = ~BUF2_REG_19__SCAN_IN | ~n41095;
  assign n30090 = ~n31027 & ~n30800;
  assign n31031 = ~n31802 & ~n30705;
  assign n30088 = ~n31031 | ~n30801;
  assign n30087 = ~P3_INSTQUEUE_REG_6__3__SCAN_IN | ~n30802;
  assign n30089 = ~n30088 | ~n30087;
  assign n30091 = ~n30090 & ~n30089;
  assign P3_U2919 = ~n30092 | ~n30091;
  assign n30094 = ~n31026 & ~n30809;
  assign n30093 = ~n31045 & ~n31027;
  assign n30100 = ~n30094 & ~n30093;
  assign n30098 = ~n30812 & ~n31030;
  assign n30096 = ~n31031 | ~n30813;
  assign n30095 = ~P3_INSTQUEUE_REG_4__3__SCAN_IN | ~n30814;
  assign n30097 = ~n30096 | ~n30095;
  assign n30099 = ~n30098 & ~n30097;
  assign P3_U2903 = ~n30100 | ~n30099;
  assign n30102 = ~n31026 & ~n30786;
  assign n30101 = ~n31030 & ~n30993;
  assign n30108 = ~n30102 & ~n30101;
  assign n30106 = ~n31027 & ~n30832;
  assign n30104 = ~n31031 | ~n30789;
  assign n30103 = ~P3_INSTQUEUE_REG_14__3__SCAN_IN | ~n30790;
  assign n30105 = ~n30104 | ~n30103;
  assign n30107 = ~n30106 & ~n30105;
  assign P3_U2983 = ~n30108 | ~n30107;
  assign n30110 = ~n31026 & ~n30761;
  assign n30109 = ~n31030 & ~n30777;
  assign n30116 = ~n30110 & ~n30109;
  assign n30114 = ~n31027 & ~n30764;
  assign n30112 = ~n31031 | ~n30765;
  assign n30111 = ~P3_INSTQUEUE_REG_10__3__SCAN_IN | ~n30766;
  assign n30113 = ~n30112 | ~n30111;
  assign n30115 = ~n30114 & ~n30113;
  assign P3_U2951 = ~n30116 | ~n30115;
  assign n30118 = ~n31026 & ~n30774;
  assign n30117 = ~n31030 & ~n30773;
  assign n30124 = ~n30118 & ~n30117;
  assign n30122 = ~n31027 & ~n30777;
  assign n30120 = ~n31031 | ~n30778;
  assign n30119 = ~P3_INSTQUEUE_REG_9__3__SCAN_IN | ~n30779;
  assign n30121 = ~n30120 | ~n30119;
  assign n30123 = ~n30122 & ~n30121;
  assign P3_U2943 = ~n30124 | ~n30123;
  assign n30126 = ~n31026 & ~n30702;
  assign n30125 = ~n31027 & ~n30990;
  assign n30132 = ~n30126 & ~n30125;
  assign n30130 = ~n31030 & ~n30750;
  assign n30128 = ~n31031 | ~n30707;
  assign n30127 = ~P3_INSTQUEUE_REG_12__3__SCAN_IN | ~n30708;
  assign n30129 = ~n30128 | ~n30127;
  assign n30131 = ~n30130 & ~n30129;
  assign P3_U2967 = ~n30132 | ~n30131;
  assign n30917 = ~BUF2_REG_5__SCAN_IN | ~n30874;
  assign n30134 = ~n30917 & ~n30702;
  assign n30921 = ~BUF2_REG_21__SCAN_IN | ~n41095;
  assign n30133 = ~n30921 & ~n30990;
  assign n30140 = ~n30134 & ~n30133;
  assign n30918 = ~BUF2_REG_29__SCAN_IN | ~n41095;
  assign n30138 = ~n30918 & ~n30750;
  assign n30922 = ~n32475 & ~n30705;
  assign n30136 = ~n30922 | ~n30707;
  assign n30135 = ~P3_INSTQUEUE_REG_12__5__SCAN_IN | ~n30708;
  assign n30137 = ~n30136 | ~n30135;
  assign n30139 = ~n30138 & ~n30137;
  assign P3_U2969 = ~n30140 | ~n30139;
  assign n30142 = ~n30917 & ~n30761;
  assign n30141 = ~n30921 & ~n30764;
  assign n30148 = ~n30142 & ~n30141;
  assign n30146 = ~n30918 & ~n30777;
  assign n30144 = ~n30922 | ~n30765;
  assign n30143 = ~P3_INSTQUEUE_REG_10__5__SCAN_IN | ~n30766;
  assign n30145 = ~n30144 | ~n30143;
  assign n30147 = ~n30146 & ~n30145;
  assign P3_U2953 = ~n30148 | ~n30147;
  assign n30150 = ~n30917 & ~n30797;
  assign n30149 = ~n30918 & ~n31040;
  assign n30156 = ~n30150 & ~n30149;
  assign n30154 = ~n30921 & ~n30800;
  assign n30152 = ~n30922 | ~n30801;
  assign n30151 = ~P3_INSTQUEUE_REG_6__5__SCAN_IN | ~n30802;
  assign n30153 = ~n30152 | ~n30151;
  assign n30155 = ~n30154 & ~n30153;
  assign P3_U2921 = ~n30156 | ~n30155;
  assign n30158 = ~n30917 & ~n30786;
  assign n30157 = ~n30918 & ~n30993;
  assign n30164 = ~n30158 & ~n30157;
  assign n30162 = ~n30921 & ~n30832;
  assign n30160 = ~n30922 | ~n30789;
  assign n30159 = ~P3_INSTQUEUE_REG_14__5__SCAN_IN | ~n30790;
  assign n30161 = ~n30160 | ~n30159;
  assign n30163 = ~n30162 & ~n30161;
  assign P3_U2985 = ~n30164 | ~n30163;
  assign n30168 = ~n30737 & ~n31026;
  assign n30166 = ~P3_INSTQUEUE_REG_8__3__SCAN_IN | ~n30742;
  assign n30165 = ~n31031 | ~n30741;
  assign n30167 = ~n30166 | ~n30165;
  assign n30172 = ~n30168 & ~n30167;
  assign n30170 = ~n31027 & ~n30773;
  assign n30169 = ~n31030 & ~n30740;
  assign n30171 = ~n30170 & ~n30169;
  assign P3_U2935 = ~n30172 | ~n30171;
  assign n30176 = ~n30726 & ~n30917;
  assign n30174 = ~P3_INSTQUEUE_REG_7__5__SCAN_IN | ~n30730;
  assign n30173 = ~n30922 | ~n30729;
  assign n30175 = ~n30174 | ~n30173;
  assign n30180 = ~n30176 & ~n30175;
  assign n30178 = ~n30921 & ~n30740;
  assign n30177 = ~n30918 & ~n30800;
  assign n30179 = ~n30178 & ~n30177;
  assign P3_U2929 = ~n30180 | ~n30179;
  assign n30184 = ~n30809 & ~n30917;
  assign n30182 = ~P3_INSTQUEUE_REG_4__5__SCAN_IN | ~n30814;
  assign n30181 = ~n30922 | ~n30813;
  assign n30183 = ~n30182 | ~n30181;
  assign n30188 = ~n30184 & ~n30183;
  assign n30186 = ~n30812 & ~n30918;
  assign n30185 = ~n31045 & ~n30921;
  assign n30187 = ~n30186 & ~n30185;
  assign P3_U2905 = ~n30188 | ~n30187;
  assign n30192 = ~n30774 & ~n30917;
  assign n30190 = ~P3_INSTQUEUE_REG_9__5__SCAN_IN | ~n30779;
  assign n30189 = ~n30922 | ~n30778;
  assign n30191 = ~n30190 | ~n30189;
  assign n30196 = ~n30192 & ~n30191;
  assign n30194 = ~n30921 & ~n30777;
  assign n30193 = ~n30918 & ~n30773;
  assign n30195 = ~n30194 & ~n30193;
  assign P3_U2945 = ~n30196 | ~n30195;
  assign n30200 = ~n30737 & ~n30917;
  assign n30198 = ~P3_INSTQUEUE_REG_8__5__SCAN_IN | ~n30742;
  assign n30197 = ~n30922 | ~n30741;
  assign n30199 = ~n30198 | ~n30197;
  assign n30204 = ~n30200 & ~n30199;
  assign n30202 = ~n30921 & ~n30773;
  assign n30201 = ~n30918 & ~n30740;
  assign n30203 = ~n30202 & ~n30201;
  assign P3_U2937 = ~n30204 | ~n30203;
  assign n30206 = ~n31026 & ~n30726;
  assign n30205 = ~n31030 & ~n30800;
  assign n30212 = ~n30206 & ~n30205;
  assign n30210 = ~n31027 & ~n30740;
  assign n30208 = ~n31031 | ~n30729;
  assign n30207 = ~P3_INSTQUEUE_REG_7__3__SCAN_IN | ~n30730;
  assign n30209 = ~n30208 | ~n30207;
  assign n30211 = ~n30210 & ~n30209;
  assign P3_U2927 = ~n30212 | ~n30211;
  assign n30833 = ~n30213 | ~n41382;
  assign n30219 = ~n30833 & ~n31014;
  assign n30215 = ~n30870 & ~n30558;
  assign n30214 = ~P3_STATE2_REG_3__SCAN_IN | ~n30861;
  assign n30838 = ~n30215 | ~n30214;
  assign n30217 = ~P3_INSTQUEUE_REG_15__4__SCAN_IN | ~n30838;
  assign n30216 = ~n30837 | ~n31019;
  assign n30218 = ~n30217 | ~n30216;
  assign n30223 = ~n30219 & ~n30218;
  assign n30221 = ~n31018 & ~n30832;
  assign n30220 = ~n31015 & ~n30836;
  assign n30222 = ~n30221 & ~n30220;
  assign P3_U2992 = ~n30223 | ~n30222;
  assign n30929 = ~BUF2_REG_1__SCAN_IN | ~n30874;
  assign n30225 = ~n30929 & ~n30786;
  assign n30930 = ~BUF2_REG_17__SCAN_IN | ~n41095;
  assign n30224 = ~n30930 & ~n30832;
  assign n30231 = ~n30225 & ~n30224;
  assign n30933 = ~BUF2_REG_25__SCAN_IN | ~n41095;
  assign n30229 = ~n30933 & ~n30993;
  assign n30934 = ~n33487 & ~n30705;
  assign n30227 = ~n30934 | ~n30789;
  assign n30226 = ~P3_INSTQUEUE_REG_14__1__SCAN_IN | ~n30790;
  assign n30228 = ~n30227 | ~n30226;
  assign n30230 = ~n30229 & ~n30228;
  assign P3_U2981 = ~n30231 | ~n30230;
  assign n30233 = ~n30929 & ~n30726;
  assign n30232 = ~n30930 & ~n30740;
  assign n30239 = ~n30233 & ~n30232;
  assign n30237 = ~n30933 & ~n30800;
  assign n30235 = ~n30934 | ~n30729;
  assign n30234 = ~P3_INSTQUEUE_REG_7__1__SCAN_IN | ~n30730;
  assign n30236 = ~n30235 | ~n30234;
  assign n30238 = ~n30237 & ~n30236;
  assign P3_U2925 = ~n30239 | ~n30238;
  assign n30241 = ~n30929 & ~n30761;
  assign n30240 = ~n30930 & ~n30764;
  assign n30247 = ~n30241 & ~n30240;
  assign n30245 = ~n30933 & ~n30777;
  assign n30243 = ~n30934 | ~n30765;
  assign n30242 = ~P3_INSTQUEUE_REG_10__1__SCAN_IN | ~n30766;
  assign n30244 = ~n30243 | ~n30242;
  assign n30246 = ~n30245 & ~n30244;
  assign P3_U2949 = ~n30247 | ~n30246;
  assign n30249 = ~n30929 & ~n30737;
  assign n30248 = ~n30933 & ~n30740;
  assign n30255 = ~n30249 & ~n30248;
  assign n30253 = ~n30930 & ~n30773;
  assign n30251 = ~n30934 | ~n30741;
  assign n30250 = ~P3_INSTQUEUE_REG_8__1__SCAN_IN | ~n30742;
  assign n30252 = ~n30251 | ~n30250;
  assign n30254 = ~n30253 & ~n30252;
  assign P3_U2933 = ~n30255 | ~n30254;
  assign n30257 = ~n30929 & ~n30797;
  assign n30256 = ~n30930 & ~n30800;
  assign n30263 = ~n30257 & ~n30256;
  assign n30261 = ~n30933 & ~n31040;
  assign n30259 = ~n30934 | ~n30801;
  assign n30258 = ~P3_INSTQUEUE_REG_6__1__SCAN_IN | ~n30802;
  assign n30260 = ~n30259 | ~n30258;
  assign n30262 = ~n30261 & ~n30260;
  assign P3_U2917 = ~n30263 | ~n30262;
  assign n30267 = ~n30821 & ~n31026;
  assign n30265 = ~P3_INSTQUEUE_REG_0__3__SCAN_IN | ~n30825;
  assign n30264 = ~n30824 | ~n31031;
  assign n30266 = ~n30265 | ~n30264;
  assign n30271 = ~n30267 & ~n30266;
  assign n30269 = ~n31027 & ~n30857;
  assign n30268 = ~n31030 & ~n30836;
  assign n30270 = ~n30269 & ~n30268;
  assign P3_U2871 = ~n30271 | ~n30270;
  assign n30273 = ~n30845 & ~n31026;
  assign n30272 = ~n30848 & ~n31027;
  assign n30279 = ~n30273 & ~n30272;
  assign n30277 = ~n30861 & ~n31030;
  assign n30275 = ~n30849 | ~n31031;
  assign n30274 = ~P3_INSTQUEUE_REG_2__3__SCAN_IN | ~n30850;
  assign n30276 = ~n30275 | ~n30274;
  assign n30278 = ~n30277 & ~n30276;
  assign P3_U2887 = ~n30279 | ~n30278;
  assign n31039 = ~BUF2_REG_7__SCAN_IN | ~n30874;
  assign n30281 = ~n31039 & ~n30737;
  assign n31041 = ~BUF2_REG_23__SCAN_IN | ~n41095;
  assign n30280 = ~n31041 & ~n30773;
  assign n30287 = ~n30281 & ~n30280;
  assign n31044 = ~BUF2_REG_31__SCAN_IN | ~n41095;
  assign n30285 = ~n31044 & ~n30740;
  assign n31046 = ~n32672 & ~n30705;
  assign n30283 = ~n31046 | ~n30741;
  assign n30282 = ~P3_INSTQUEUE_REG_8__7__SCAN_IN | ~n30742;
  assign n30284 = ~n30283 | ~n30282;
  assign n30286 = ~n30285 & ~n30284;
  assign P3_U2939 = ~n30287 | ~n30286;
  assign n30289 = ~n31039 & ~n30797;
  assign n30288 = ~n31041 & ~n30800;
  assign n30295 = ~n30289 & ~n30288;
  assign n30293 = ~n31044 & ~n31040;
  assign n30291 = ~n31046 | ~n30801;
  assign n30290 = ~P3_INSTQUEUE_REG_6__7__SCAN_IN | ~n30802;
  assign n30292 = ~n30291 | ~n30290;
  assign n30294 = ~n30293 & ~n30292;
  assign P3_U2923 = ~n30295 | ~n30294;
  assign n30297 = ~n31039 & ~n30761;
  assign n30296 = ~n31041 & ~n30764;
  assign n30303 = ~n30297 & ~n30296;
  assign n30301 = ~n31044 & ~n30777;
  assign n30299 = ~n31046 | ~n30765;
  assign n30298 = ~P3_INSTQUEUE_REG_10__7__SCAN_IN | ~n30766;
  assign n30300 = ~n30299 | ~n30298;
  assign n30302 = ~n30301 & ~n30300;
  assign P3_U2955 = ~n30303 | ~n30302;
  assign n30305 = ~n31039 & ~n30786;
  assign n30304 = ~n31041 & ~n30832;
  assign n30311 = ~n30305 & ~n30304;
  assign n30309 = ~n31044 & ~n30993;
  assign n30307 = ~n31046 | ~n30789;
  assign n30306 = ~P3_INSTQUEUE_REG_14__7__SCAN_IN | ~n30790;
  assign n30308 = ~n30307 | ~n30306;
  assign n30310 = ~n30309 & ~n30308;
  assign P3_U2987 = ~n30311 | ~n30310;
  assign n30313 = ~n31039 & ~n30726;
  assign n30312 = ~n31041 & ~n30740;
  assign n30319 = ~n30313 & ~n30312;
  assign n30317 = ~n31044 & ~n30800;
  assign n30315 = ~n31046 | ~n30729;
  assign n30314 = ~P3_INSTQUEUE_REG_7__7__SCAN_IN | ~n30730;
  assign n30316 = ~n30315 | ~n30314;
  assign n30318 = ~n30317 & ~n30316;
  assign P3_U2931 = ~n30319 | ~n30318;
  assign n30321 = ~n31039 & ~n30702;
  assign n30320 = ~n31041 & ~n30990;
  assign n30327 = ~n30321 & ~n30320;
  assign n30325 = ~n31044 & ~n30750;
  assign n30323 = ~n31046 | ~n30707;
  assign n30322 = ~P3_INSTQUEUE_REG_12__7__SCAN_IN | ~n30708;
  assign n30324 = ~n30323 | ~n30322;
  assign n30326 = ~n30325 & ~n30324;
  assign P3_U2971 = ~n30327 | ~n30326;
  assign n30329 = ~n30917 & ~n30821;
  assign n30328 = ~n30918 & ~n30836;
  assign n30335 = ~n30329 & ~n30328;
  assign n30333 = ~n30921 & ~n30857;
  assign n30331 = ~n30824 | ~n30922;
  assign n30330 = ~P3_INSTQUEUE_REG_0__5__SCAN_IN | ~n30825;
  assign n30332 = ~n30331 | ~n30330;
  assign n30334 = ~n30333 & ~n30332;
  assign P3_U2873 = ~n30335 | ~n30334;
  assign n30337 = ~n31039 & ~n30809;
  assign n30336 = ~n30812 & ~n31044;
  assign n30343 = ~n30337 & ~n30336;
  assign n30341 = ~n31045 & ~n31041;
  assign n30339 = ~n31046 | ~n30813;
  assign n30338 = ~P3_INSTQUEUE_REG_4__7__SCAN_IN | ~n30814;
  assign n30340 = ~n30339 | ~n30338;
  assign n30342 = ~n30341 & ~n30340;
  assign P3_U2907 = ~n30343 | ~n30342;
  assign n30347 = ~n30809 & ~n30929;
  assign n30345 = ~P3_INSTQUEUE_REG_4__1__SCAN_IN | ~n30814;
  assign n30344 = ~n30934 | ~n30813;
  assign n30346 = ~n30345 | ~n30344;
  assign n30351 = ~n30347 & ~n30346;
  assign n30349 = ~n30812 & ~n30933;
  assign n30348 = ~n31045 & ~n30930;
  assign n30350 = ~n30349 & ~n30348;
  assign P3_U2901 = ~n30351 | ~n30350;
  assign n30355 = ~n30774 & ~n30929;
  assign n30353 = ~P3_INSTQUEUE_REG_9__1__SCAN_IN | ~n30779;
  assign n30352 = ~n30934 | ~n30778;
  assign n30354 = ~n30353 | ~n30352;
  assign n30359 = ~n30355 & ~n30354;
  assign n30357 = ~n30933 & ~n30773;
  assign n30356 = ~n30930 & ~n30777;
  assign n30358 = ~n30357 & ~n30356;
  assign P3_U2941 = ~n30359 | ~n30358;
  assign n30363 = ~n30702 & ~n30929;
  assign n30361 = ~P3_INSTQUEUE_REG_12__1__SCAN_IN | ~n30708;
  assign n30360 = ~n30934 | ~n30707;
  assign n30362 = ~n30361 | ~n30360;
  assign n30367 = ~n30363 & ~n30362;
  assign n30365 = ~n30933 & ~n30750;
  assign n30364 = ~n30930 & ~n30990;
  assign n30366 = ~n30365 & ~n30364;
  assign P3_U2965 = ~n30367 | ~n30366;
  assign n30369 = ~n30845 & ~n30917;
  assign n30368 = ~n30848 & ~n30921;
  assign n30375 = ~n30369 & ~n30368;
  assign n30373 = ~n30861 & ~n30918;
  assign n30371 = ~n30849 | ~n30922;
  assign n30370 = ~P3_INSTQUEUE_REG_2__5__SCAN_IN | ~n30850;
  assign n30372 = ~n30371 | ~n30370;
  assign n30374 = ~n30373 & ~n30372;
  assign P3_U2889 = ~n30375 | ~n30374;
  assign n30379 = ~n30858 & ~n31026;
  assign n30377 = ~P3_INSTQUEUE_REG_1__3__SCAN_IN | ~n30863;
  assign n30376 = ~n30862 | ~n31031;
  assign n30378 = ~n30377 | ~n30376;
  assign n30383 = ~n30379 & ~n30378;
  assign n30381 = ~n31030 & ~n30857;
  assign n30380 = ~n30861 & ~n31027;
  assign n30382 = ~n30381 & ~n30380;
  assign P3_U2879 = ~n30383 | ~n30382;
  assign n30387 = ~n30774 & ~n31039;
  assign n30385 = ~P3_INSTQUEUE_REG_9__7__SCAN_IN | ~n30779;
  assign n30384 = ~n31046 | ~n30778;
  assign n30386 = ~n30385 | ~n30384;
  assign n30391 = ~n30387 & ~n30386;
  assign n30389 = ~n31044 & ~n30773;
  assign n30388 = ~n31041 & ~n30777;
  assign n30390 = ~n30389 & ~n30388;
  assign P3_U2947 = ~n30391 | ~n30390;
  assign n30395 = ~n30858 & ~n30917;
  assign n30393 = ~P3_INSTQUEUE_REG_1__5__SCAN_IN | ~n30863;
  assign n30392 = ~n30862 | ~n30922;
  assign n30394 = ~n30393 | ~n30392;
  assign n30399 = ~n30395 & ~n30394;
  assign n30397 = ~n30918 & ~n30857;
  assign n30396 = ~n30861 & ~n30921;
  assign n30398 = ~n30397 & ~n30396;
  assign P3_U2881 = ~n30399 | ~n30398;
  assign n30401 = ~n31039 & ~n30821;
  assign n30400 = ~n31041 & ~n30857;
  assign n30407 = ~n30401 & ~n30400;
  assign n30405 = ~n31044 & ~n30836;
  assign n30403 = ~n30824 | ~n31046;
  assign n30402 = ~P3_INSTQUEUE_REG_0__7__SCAN_IN | ~n30825;
  assign n30404 = ~n30403 | ~n30402;
  assign n30406 = ~n30405 & ~n30404;
  assign P3_U2875 = ~n30407 | ~n30406;
  assign n30409 = ~n30929 & ~n30821;
  assign n30408 = ~n30933 & ~n30836;
  assign n30415 = ~n30409 & ~n30408;
  assign n30413 = ~n30930 & ~n30857;
  assign n30411 = ~n30824 | ~n30934;
  assign n30410 = ~P3_INSTQUEUE_REG_0__1__SCAN_IN | ~n30825;
  assign n30412 = ~n30411 | ~n30410;
  assign n30414 = ~n30413 & ~n30412;
  assign P3_U2869 = ~n30415 | ~n30414;
  assign n30417 = ~n30845 & ~n31039;
  assign n30416 = ~n30861 & ~n31044;
  assign n30423 = ~n30417 & ~n30416;
  assign n30421 = ~n30848 & ~n31041;
  assign n30419 = ~n30849 | ~n31046;
  assign n30418 = ~P3_INSTQUEUE_REG_2__7__SCAN_IN | ~n30850;
  assign n30420 = ~n30419 | ~n30418;
  assign n30422 = ~n30421 & ~n30420;
  assign P3_U2891 = ~n30423 | ~n30422;
  assign n30425 = ~n30845 & ~n30929;
  assign n30424 = ~n30861 & ~n30933;
  assign n30431 = ~n30425 & ~n30424;
  assign n30429 = ~n30848 & ~n30930;
  assign n30427 = ~n30849 | ~n30934;
  assign n30426 = ~P3_INSTQUEUE_REG_2__1__SCAN_IN | ~n30850;
  assign n30428 = ~n30427 | ~n30426;
  assign n30430 = ~n30429 & ~n30428;
  assign P3_U2885 = ~n30431 | ~n30430;
  assign n30435 = ~n30858 & ~n31039;
  assign n30433 = ~P3_INSTQUEUE_REG_1__7__SCAN_IN | ~n30863;
  assign n30432 = ~n30862 | ~n31046;
  assign n30434 = ~n30433 | ~n30432;
  assign n30439 = ~n30435 & ~n30434;
  assign n30437 = ~n31044 & ~n30857;
  assign n30436 = ~n30861 & ~n31041;
  assign n30438 = ~n30437 & ~n30436;
  assign P3_U2883 = ~n30439 | ~n30438;
  assign n30977 = ~BUF2_REG_0__SCAN_IN | ~n30874;
  assign n30441 = ~n30977 & ~n30774;
  assign n30978 = ~BUF2_REG_16__SCAN_IN | ~n41095;
  assign n30440 = ~n30978 & ~n30777;
  assign n30447 = ~n30441 & ~n30440;
  assign n30981 = ~BUF2_REG_24__SCAN_IN | ~n41095;
  assign n30445 = ~n30981 & ~n30773;
  assign n30982 = ~n33501 & ~n30705;
  assign n30443 = ~n30982 | ~n30778;
  assign n30442 = ~P3_INSTQUEUE_REG_9__0__SCAN_IN | ~n30779;
  assign n30444 = ~n30443 | ~n30442;
  assign n30446 = ~n30445 & ~n30444;
  assign P3_U2940 = ~n30447 | ~n30446;
  assign n30449 = ~n30977 & ~n30786;
  assign n30448 = ~n30978 & ~n30832;
  assign n30455 = ~n30449 & ~n30448;
  assign n30453 = ~n30981 & ~n30993;
  assign n30451 = ~n30982 | ~n30789;
  assign n30450 = ~P3_INSTQUEUE_REG_14__0__SCAN_IN | ~n30790;
  assign n30452 = ~n30451 | ~n30450;
  assign n30454 = ~n30453 & ~n30452;
  assign P3_U2980 = ~n30455 | ~n30454;
  assign n30457 = ~n30977 & ~n30809;
  assign n30456 = ~n31045 & ~n30978;
  assign n30463 = ~n30457 & ~n30456;
  assign n30461 = ~n30981 & ~n30812;
  assign n30459 = ~n30982 | ~n30813;
  assign n30458 = ~P3_INSTQUEUE_REG_4__0__SCAN_IN | ~n30814;
  assign n30460 = ~n30459 | ~n30458;
  assign n30462 = ~n30461 & ~n30460;
  assign P3_U2900 = ~n30463 | ~n30462;
  assign n30465 = ~n30977 & ~n30761;
  assign n30464 = ~n30981 & ~n30777;
  assign n30471 = ~n30465 & ~n30464;
  assign n30469 = ~n30978 & ~n30764;
  assign n30467 = ~n30982 | ~n30765;
  assign n30466 = ~P3_INSTQUEUE_REG_10__0__SCAN_IN | ~n30766;
  assign n30468 = ~n30467 | ~n30466;
  assign n30470 = ~n30469 & ~n30468;
  assign P3_U2948 = ~n30471 | ~n30470;
  assign n30473 = ~n30977 & ~n30737;
  assign n30472 = ~n30981 & ~n30740;
  assign n30479 = ~n30473 & ~n30472;
  assign n30477 = ~n30978 & ~n30773;
  assign n30475 = ~n30982 | ~n30741;
  assign n30474 = ~P3_INSTQUEUE_REG_8__0__SCAN_IN | ~n30742;
  assign n30476 = ~n30475 | ~n30474;
  assign n30478 = ~n30477 & ~n30476;
  assign P3_U2932 = ~n30479 | ~n30478;
  assign n30481 = ~n30977 & ~n30702;
  assign n30480 = ~n30978 & ~n30990;
  assign n30487 = ~n30481 & ~n30480;
  assign n30485 = ~n30981 & ~n30750;
  assign n30483 = ~n30982 | ~n30707;
  assign n30482 = ~P3_INSTQUEUE_REG_12__0__SCAN_IN | ~n30708;
  assign n30484 = ~n30483 | ~n30482;
  assign n30486 = ~n30485 & ~n30484;
  assign P3_U2964 = ~n30487 | ~n30486;
  assign n30489 = ~n30977 & ~n30797;
  assign n30488 = ~n30978 & ~n30800;
  assign n30495 = ~n30489 & ~n30488;
  assign n30493 = ~n30981 & ~n31040;
  assign n30491 = ~n30982 | ~n30801;
  assign n30490 = ~P3_INSTQUEUE_REG_6__0__SCAN_IN | ~n30802;
  assign n30492 = ~n30491 | ~n30490;
  assign n30494 = ~n30493 & ~n30492;
  assign P3_U2916 = ~n30495 | ~n30494;
  assign n30497 = ~n30977 & ~n30726;
  assign n30496 = ~n30978 & ~n30740;
  assign n30503 = ~n30497 & ~n30496;
  assign n30501 = ~n30981 & ~n30800;
  assign n30499 = ~n30982 | ~n30729;
  assign n30498 = ~P3_INSTQUEUE_REG_7__0__SCAN_IN | ~n30730;
  assign n30500 = ~n30499 | ~n30498;
  assign n30502 = ~n30501 & ~n30500;
  assign P3_U2924 = ~n30503 | ~n30502;
  assign n30507 = ~n30858 & ~n30929;
  assign n30505 = ~P3_INSTQUEUE_REG_1__1__SCAN_IN | ~n30863;
  assign n30504 = ~n30862 | ~n30934;
  assign n30506 = ~n30505 | ~n30504;
  assign n30511 = ~n30507 & ~n30506;
  assign n30509 = ~n30933 & ~n30857;
  assign n30508 = ~n30861 & ~n30930;
  assign n30510 = ~n30509 & ~n30508;
  assign P3_U2877 = ~n30511 | ~n30510;
  assign n30513 = ~n31002 & ~n30836;
  assign n30512 = ~n31003 & ~n30833;
  assign n30519 = ~n30513 & ~n30512;
  assign n30517 = ~n31006 & ~n30832;
  assign n30515 = ~n30837 | ~n31007;
  assign n30514 = ~P3_INSTQUEUE_REG_15__2__SCAN_IN | ~n30838;
  assign n30516 = ~n30515 | ~n30514;
  assign n30518 = ~n30517 & ~n30516;
  assign P3_U2990 = ~n30519 | ~n30518;
  assign n30521 = ~n30917 & ~n30833;
  assign n30520 = ~n30921 & ~n30836;
  assign n30527 = ~n30521 & ~n30520;
  assign n30525 = ~n30918 & ~n30832;
  assign n30523 = ~n30837 | ~n30922;
  assign n30522 = ~P3_INSTQUEUE_REG_15__5__SCAN_IN | ~n30838;
  assign n30524 = ~n30523 | ~n30522;
  assign n30526 = ~n30525 & ~n30524;
  assign P3_U2993 = ~n30527 | ~n30526;
  assign n30529 = ~n30929 & ~n30833;
  assign n30528 = ~n30930 & ~n30836;
  assign n30535 = ~n30529 & ~n30528;
  assign n30533 = ~n30933 & ~n30832;
  assign n30531 = ~n30837 | ~n30934;
  assign n30530 = ~P3_INSTQUEUE_REG_15__1__SCAN_IN | ~n30838;
  assign n30532 = ~n30531 | ~n30530;
  assign n30534 = ~n30533 & ~n30532;
  assign P3_U2989 = ~n30535 | ~n30534;
  assign n30537 = ~n31026 & ~n30833;
  assign n30536 = ~n31027 & ~n30836;
  assign n30543 = ~n30537 & ~n30536;
  assign n30541 = ~n31030 & ~n30832;
  assign n30539 = ~n30837 | ~n31031;
  assign n30538 = ~P3_INSTQUEUE_REG_15__3__SCAN_IN | ~n30838;
  assign n30540 = ~n30539 | ~n30538;
  assign n30542 = ~n30541 & ~n30540;
  assign P3_U2991 = ~n30543 | ~n30542;
  assign n30545 = ~n31039 & ~n30833;
  assign n30544 = ~n31044 & ~n30832;
  assign n30551 = ~n30545 & ~n30544;
  assign n30549 = ~n31041 & ~n30836;
  assign n30547 = ~n30837 | ~n31046;
  assign n30546 = ~P3_INSTQUEUE_REG_15__7__SCAN_IN | ~n30838;
  assign n30548 = ~n30547 | ~n30546;
  assign n30550 = ~n30549 & ~n30548;
  assign P3_U2995 = ~n30551 | ~n30550;
  assign n30557 = ~n30848 & ~n30981;
  assign n30715 = ~n30900 | ~n41382;
  assign n30553 = ~n30977 & ~n30715;
  assign n30552 = ~n30812 & ~n30978;
  assign n30555 = ~n30553 & ~n30552;
  assign n30718 = ~n31040;
  assign n30554 = ~n30982 | ~n30718;
  assign n30556 = ~n30555 | ~n30554;
  assign n30562 = ~n30557 & ~n30556;
  assign n30599 = ~n30559 & ~n30558;
  assign n30719 = ~n30560 | ~n30599;
  assign n30561 = ~P3_INSTQUEUE_REG_3__0__SCAN_IN | ~n30719;
  assign P3_U2892 = ~n30562 | ~n30561;
  assign n30566 = ~n30977 & ~n30821;
  assign n30564 = ~n30824 | ~n30982;
  assign n30563 = ~P3_INSTQUEUE_REG_0__0__SCAN_IN | ~n30825;
  assign n30565 = ~n30564 | ~n30563;
  assign n30570 = ~n30566 & ~n30565;
  assign n30568 = ~n30978 & ~n30857;
  assign n30567 = ~n30981 & ~n30836;
  assign n30569 = ~n30568 & ~n30567;
  assign P3_U2868 = ~n30570 | ~n30569;
  assign n30574 = ~n30977 & ~n30833;
  assign n30572 = ~n30837 | ~n30982;
  assign n30571 = ~P3_INSTQUEUE_REG_15__0__SCAN_IN | ~n30838;
  assign n30573 = ~n30572 | ~n30571;
  assign n30578 = ~n30574 & ~n30573;
  assign n30576 = ~n30978 & ~n30836;
  assign n30575 = ~n30981 & ~n30832;
  assign n30577 = ~n30576 & ~n30575;
  assign P3_U2988 = ~n30578 | ~n30577;
  assign n30584 = ~n30981 & ~n30861;
  assign n30580 = ~n30977 & ~n30845;
  assign n30579 = ~n30848 & ~n30978;
  assign n30582 = ~n30580 & ~n30579;
  assign n30581 = ~n30849 | ~n30982;
  assign n30583 = ~n30582 | ~n30581;
  assign n30586 = ~n30584 & ~n30583;
  assign n30585 = ~P3_INSTQUEUE_REG_2__0__SCAN_IN | ~n30850;
  assign P3_U2884 = ~n30586 | ~n30585;
  assign n30588 = ~n30977 & ~n30858;
  assign n30587 = ~n30861 & ~n30978;
  assign n30594 = ~n30588 & ~n30587;
  assign n30592 = ~n30981 & ~n30857;
  assign n30590 = ~n30862 | ~n30982;
  assign n30589 = ~P3_INSTQUEUE_REG_1__0__SCAN_IN | ~n30863;
  assign n30591 = ~n30590 | ~n30589;
  assign n30593 = ~n30592 & ~n30591;
  assign P3_U2876 = ~n30594 | ~n30593;
  assign n30749 = ~n30877 | ~n41382;
  assign n30596 = ~n31003 & ~n30749;
  assign n30595 = ~n31006 & ~n30764;
  assign n30605 = ~n30596 & ~n30595;
  assign n30603 = ~n31002 & ~n30750;
  assign n30753 = ~n30993;
  assign n30601 = ~n31007 | ~n30753;
  assign n30598 = ~n30597;
  assign n30754 = ~n30599 | ~n30598;
  assign n30600 = ~P3_INSTQUEUE_REG_11__2__SCAN_IN | ~n30754;
  assign n30602 = ~n30601 | ~n30600;
  assign n30604 = ~n30603 & ~n30602;
  assign P3_U2958 = ~n30605 | ~n30604;
  assign n30607 = ~n30977 & ~n30749;
  assign n30606 = ~n30981 & ~n30764;
  assign n30613 = ~n30607 & ~n30606;
  assign n30611 = ~n30978 & ~n30750;
  assign n30609 = ~n30982 | ~n30753;
  assign n30608 = ~P3_INSTQUEUE_REG_11__0__SCAN_IN | ~n30754;
  assign n30610 = ~n30609 | ~n30608;
  assign n30612 = ~n30611 & ~n30610;
  assign P3_U2956 = ~n30613 | ~n30612;
  assign n30615 = ~n31026 & ~n30749;
  assign n30614 = ~n31030 & ~n30764;
  assign n30621 = ~n30615 & ~n30614;
  assign n30619 = ~n31027 & ~n30750;
  assign n30617 = ~n31031 | ~n30753;
  assign n30616 = ~P3_INSTQUEUE_REG_11__3__SCAN_IN | ~n30754;
  assign n30618 = ~n30617 | ~n30616;
  assign n30620 = ~n30619 & ~n30618;
  assign P3_U2959 = ~n30621 | ~n30620;
  assign n30623 = ~n30929 & ~n30749;
  assign n30622 = ~n30930 & ~n30750;
  assign n30629 = ~n30623 & ~n30622;
  assign n30627 = ~n30933 & ~n30764;
  assign n30625 = ~n30934 | ~n30753;
  assign n30624 = ~P3_INSTQUEUE_REG_11__1__SCAN_IN | ~n30754;
  assign n30626 = ~n30625 | ~n30624;
  assign n30628 = ~n30627 & ~n30626;
  assign P3_U2957 = ~n30629 | ~n30628;
  assign n30631 = ~n31014 & ~n30749;
  assign n30630 = ~n31015 & ~n30750;
  assign n30637 = ~n30631 & ~n30630;
  assign n30635 = ~n31018 & ~n30764;
  assign n30633 = ~n31019 | ~n30753;
  assign n30632 = ~P3_INSTQUEUE_REG_11__4__SCAN_IN | ~n30754;
  assign n30634 = ~n30633 | ~n30632;
  assign n30636 = ~n30635 & ~n30634;
  assign P3_U2960 = ~n30637 | ~n30636;
  assign n30639 = ~n30917 & ~n30749;
  assign n30638 = ~n30921 & ~n30750;
  assign n30645 = ~n30639 & ~n30638;
  assign n30643 = ~n30918 & ~n30764;
  assign n30641 = ~n30922 | ~n30753;
  assign n30640 = ~P3_INSTQUEUE_REG_11__5__SCAN_IN | ~n30754;
  assign n30642 = ~n30641 | ~n30640;
  assign n30644 = ~n30643 & ~n30642;
  assign P3_U2961 = ~n30645 | ~n30644;
  assign n30647 = ~n31039 & ~n30749;
  assign n30646 = ~n31044 & ~n30764;
  assign n30653 = ~n30647 & ~n30646;
  assign n30651 = ~n31041 & ~n30750;
  assign n30649 = ~n31046 | ~n30753;
  assign n30648 = ~P3_INSTQUEUE_REG_11__7__SCAN_IN | ~n30754;
  assign n30650 = ~n30649 | ~n30648;
  assign n30652 = ~n30651 & ~n30650;
  assign P3_U2963 = ~n30653 | ~n30652;
  assign n30655 = ~n31003 & ~n30715;
  assign n30654 = ~n30848 & ~n31006;
  assign n30661 = ~n30655 & ~n30654;
  assign n30659 = ~n30812 & ~n31002;
  assign n30657 = ~n31007 | ~n30718;
  assign n30656 = ~P3_INSTQUEUE_REG_3__2__SCAN_IN | ~n30719;
  assign n30658 = ~n30657 | ~n30656;
  assign n30660 = ~n30659 & ~n30658;
  assign P3_U2894 = ~n30661 | ~n30660;
  assign n30663 = ~n31039 & ~n30715;
  assign n30662 = ~n30848 & ~n31044;
  assign n30669 = ~n30663 & ~n30662;
  assign n30667 = ~n30812 & ~n31041;
  assign n30665 = ~n31046 | ~n30718;
  assign n30664 = ~P3_INSTQUEUE_REG_3__7__SCAN_IN | ~n30719;
  assign n30666 = ~n30665 | ~n30664;
  assign n30668 = ~n30667 & ~n30666;
  assign P3_U2899 = ~n30669 | ~n30668;
  assign n30671 = ~n31014 & ~n30715;
  assign n30670 = ~n30812 & ~n31015;
  assign n30677 = ~n30671 & ~n30670;
  assign n30675 = ~n30848 & ~n31018;
  assign n30673 = ~n31019 | ~n30718;
  assign n30672 = ~P3_INSTQUEUE_REG_3__4__SCAN_IN | ~n30719;
  assign n30674 = ~n30673 | ~n30672;
  assign n30676 = ~n30675 & ~n30674;
  assign P3_U2896 = ~n30677 | ~n30676;
  assign n30679 = ~n30929 & ~n30715;
  assign n30678 = ~n30812 & ~n30930;
  assign n30685 = ~n30679 & ~n30678;
  assign n30683 = ~n30848 & ~n30933;
  assign n30681 = ~n30934 | ~n30718;
  assign n30680 = ~P3_INSTQUEUE_REG_3__1__SCAN_IN | ~n30719;
  assign n30682 = ~n30681 | ~n30680;
  assign n30684 = ~n30683 & ~n30682;
  assign P3_U2893 = ~n30685 | ~n30684;
  assign n30687 = ~n31026 & ~n30715;
  assign n30686 = ~n30812 & ~n31027;
  assign n30693 = ~n30687 & ~n30686;
  assign n30691 = ~n30848 & ~n31030;
  assign n30689 = ~n31031 | ~n30718;
  assign n30688 = ~P3_INSTQUEUE_REG_3__3__SCAN_IN | ~n30719;
  assign n30690 = ~n30689 | ~n30688;
  assign n30692 = ~n30691 & ~n30690;
  assign P3_U2895 = ~n30693 | ~n30692;
  assign n30695 = ~n30917 & ~n30715;
  assign n30694 = ~n30812 & ~n30921;
  assign n30701 = ~n30695 & ~n30694;
  assign n30699 = ~n30848 & ~n30918;
  assign n30697 = ~n30922 | ~n30718;
  assign n30696 = ~P3_INSTQUEUE_REG_3__5__SCAN_IN | ~n30719;
  assign n30698 = ~n30697 | ~n30696;
  assign n30700 = ~n30699 & ~n30698;
  assign P3_U2897 = ~n30701 | ~n30700;
  assign n30965 = ~BUF2_REG_30__SCAN_IN | ~n41095;
  assign n30704 = ~n30965 & ~n30750;
  assign n30966 = ~BUF2_REG_6__SCAN_IN | ~n30874;
  assign n30703 = ~n30966 & ~n30702;
  assign n30714 = ~n30704 & ~n30703;
  assign n30969 = ~BUF2_REG_22__SCAN_IN | ~n41095;
  assign n30712 = ~n30969 & ~n30990;
  assign n30970 = ~n30706 & ~n30705;
  assign n30710 = ~n30970 | ~n30707;
  assign n30709 = ~P3_INSTQUEUE_REG_12__6__SCAN_IN | ~n30708;
  assign n30711 = ~n30710 | ~n30709;
  assign n30713 = ~n30712 & ~n30711;
  assign P3_U2970 = ~n30714 | ~n30713;
  assign n30717 = ~n30966 & ~n30715;
  assign n30716 = ~n30848 & ~n30965;
  assign n30725 = ~n30717 & ~n30716;
  assign n30723 = ~n30812 & ~n30969;
  assign n30721 = ~n30970 | ~n30718;
  assign n30720 = ~P3_INSTQUEUE_REG_3__6__SCAN_IN | ~n30719;
  assign n30722 = ~n30721 | ~n30720;
  assign n30724 = ~n30723 & ~n30722;
  assign P3_U2898 = ~n30725 | ~n30724;
  assign n30728 = ~n30966 & ~n30726;
  assign n30727 = ~n30969 & ~n30740;
  assign n30736 = ~n30728 & ~n30727;
  assign n30734 = ~n30965 & ~n30800;
  assign n30732 = ~n30970 | ~n30729;
  assign n30731 = ~P3_INSTQUEUE_REG_7__6__SCAN_IN | ~n30730;
  assign n30733 = ~n30732 | ~n30731;
  assign n30735 = ~n30734 & ~n30733;
  assign P3_U2930 = ~n30736 | ~n30735;
  assign n30739 = ~n30966 & ~n30737;
  assign n30738 = ~n30969 & ~n30773;
  assign n30748 = ~n30739 & ~n30738;
  assign n30746 = ~n30965 & ~n30740;
  assign n30744 = ~n30970 | ~n30741;
  assign n30743 = ~P3_INSTQUEUE_REG_8__6__SCAN_IN | ~n30742;
  assign n30745 = ~n30744 | ~n30743;
  assign n30747 = ~n30746 & ~n30745;
  assign P3_U2938 = ~n30748 | ~n30747;
  assign n30752 = ~n30966 & ~n30749;
  assign n30751 = ~n30969 & ~n30750;
  assign n30760 = ~n30752 & ~n30751;
  assign n30758 = ~n30965 & ~n30764;
  assign n30756 = ~n30970 | ~n30753;
  assign n30755 = ~P3_INSTQUEUE_REG_11__6__SCAN_IN | ~n30754;
  assign n30757 = ~n30756 | ~n30755;
  assign n30759 = ~n30758 & ~n30757;
  assign P3_U2962 = ~n30760 | ~n30759;
  assign n30763 = ~n30965 & ~n30777;
  assign n30762 = ~n30966 & ~n30761;
  assign n30772 = ~n30763 & ~n30762;
  assign n30770 = ~n30969 & ~n30764;
  assign n30768 = ~n30970 | ~n30765;
  assign n30767 = ~P3_INSTQUEUE_REG_10__6__SCAN_IN | ~n30766;
  assign n30769 = ~n30768 | ~n30767;
  assign n30771 = ~n30770 & ~n30769;
  assign P3_U2954 = ~n30772 | ~n30771;
  assign n30776 = ~n30965 & ~n30773;
  assign n30775 = ~n30966 & ~n30774;
  assign n30785 = ~n30776 & ~n30775;
  assign n30783 = ~n30969 & ~n30777;
  assign n30781 = ~n30970 | ~n30778;
  assign n30780 = ~P3_INSTQUEUE_REG_9__6__SCAN_IN | ~n30779;
  assign n30782 = ~n30781 | ~n30780;
  assign n30784 = ~n30783 & ~n30782;
  assign P3_U2946 = ~n30785 | ~n30784;
  assign n30788 = ~n30966 & ~n30786;
  assign n30787 = ~n30969 & ~n30832;
  assign n30796 = ~n30788 & ~n30787;
  assign n30794 = ~n30965 & ~n30993;
  assign n30792 = ~n30970 | ~n30789;
  assign n30791 = ~P3_INSTQUEUE_REG_14__6__SCAN_IN | ~n30790;
  assign n30793 = ~n30792 | ~n30791;
  assign n30795 = ~n30794 & ~n30793;
  assign P3_U2986 = ~n30796 | ~n30795;
  assign n30799 = ~n30965 & ~n31040;
  assign n30798 = ~n30966 & ~n30797;
  assign n30808 = ~n30799 & ~n30798;
  assign n30806 = ~n30969 & ~n30800;
  assign n30804 = ~n30970 | ~n30801;
  assign n30803 = ~P3_INSTQUEUE_REG_6__6__SCAN_IN | ~n30802;
  assign n30805 = ~n30804 | ~n30803;
  assign n30807 = ~n30806 & ~n30805;
  assign P3_U2922 = ~n30808 | ~n30807;
  assign n30811 = ~n30966 & ~n30809;
  assign n30810 = ~n31045 & ~n30969;
  assign n30820 = ~n30811 & ~n30810;
  assign n30818 = ~n30812 & ~n30965;
  assign n30816 = ~n30970 | ~n30813;
  assign n30815 = ~P3_INSTQUEUE_REG_4__6__SCAN_IN | ~n30814;
  assign n30817 = ~n30816 | ~n30815;
  assign n30819 = ~n30818 & ~n30817;
  assign P3_U2906 = ~n30820 | ~n30819;
  assign n30823 = ~n30965 & ~n30836;
  assign n30822 = ~n30966 & ~n30821;
  assign n30831 = ~n30823 & ~n30822;
  assign n30829 = ~n30969 & ~n30857;
  assign n30827 = ~n30824 | ~n30970;
  assign n30826 = ~P3_INSTQUEUE_REG_0__6__SCAN_IN | ~n30825;
  assign n30828 = ~n30827 | ~n30826;
  assign n30830 = ~n30829 & ~n30828;
  assign P3_U2874 = ~n30831 | ~n30830;
  assign n30835 = ~n30965 & ~n30832;
  assign n30834 = ~n30966 & ~n30833;
  assign n30844 = ~n30835 & ~n30834;
  assign n30842 = ~n30969 & ~n30836;
  assign n30840 = ~n30837 | ~n30970;
  assign n30839 = ~P3_INSTQUEUE_REG_15__6__SCAN_IN | ~n30838;
  assign n30841 = ~n30840 | ~n30839;
  assign n30843 = ~n30842 & ~n30841;
  assign P3_U2994 = ~n30844 | ~n30843;
  assign n30847 = ~n30845 & ~n30966;
  assign n30846 = ~n30861 & ~n30965;
  assign n30856 = ~n30847 & ~n30846;
  assign n30854 = ~n30848 & ~n30969;
  assign n30852 = ~n30849 | ~n30970;
  assign n30851 = ~P3_INSTQUEUE_REG_2__6__SCAN_IN | ~n30850;
  assign n30853 = ~n30852 | ~n30851;
  assign n30855 = ~n30854 & ~n30853;
  assign P3_U2890 = ~n30856 | ~n30855;
  assign n30860 = ~n30965 & ~n30857;
  assign n30859 = ~n30966 & ~n30858;
  assign n30869 = ~n30860 & ~n30859;
  assign n30867 = ~n30861 & ~n30969;
  assign n30865 = ~n30862 | ~n30970;
  assign n30864 = ~P3_INSTQUEUE_REG_1__6__SCAN_IN | ~n30863;
  assign n30866 = ~n30865 | ~n30864;
  assign n30868 = ~n30867 & ~n30866;
  assign P3_U2882 = ~n30869 | ~n30868;
  assign n30875 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n30870;
  assign n30989 = ~n30875 | ~n41382;
  assign n30872 = ~n30977 & ~n30989;
  assign n30871 = ~n30978 & ~n30993;
  assign n30885 = ~n30872 & ~n30871;
  assign n30883 = ~n30981 & ~n30990;
  assign n30881 = ~n30994 | ~n30982;
  assign n30899 = ~n30874 | ~n30873;
  assign n30876 = ~n30875;
  assign n30879 = ~n30899 & ~n30876;
  assign n30878 = n41095 & n30877;
  assign n30995 = ~n30879 & ~n30878;
  assign n30880 = ~n30995 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n30882 = ~n30881 | ~n30880;
  assign n30884 = ~n30883 & ~n30882;
  assign P3_U2972 = ~n30885 | ~n30884;
  assign n30887 = ~n31002 & ~n30993;
  assign n30886 = ~n31003 & ~n30989;
  assign n30893 = ~n30887 & ~n30886;
  assign n30891 = ~n31006 & ~n30990;
  assign n30889 = ~n30994 | ~n31007;
  assign n30888 = ~n30995 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n30890 = ~n30889 | ~n30888;
  assign n30892 = ~n30891 & ~n30890;
  assign P3_U2974 = ~n30893 | ~n30892;
  assign n30897 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n30894;
  assign n31038 = ~n30897 | ~n41382;
  assign n30896 = ~n30929 & ~n31038;
  assign n30895 = ~n31045 & ~n30933;
  assign n30908 = ~n30896 & ~n30895;
  assign n30906 = ~n30930 & ~n31040;
  assign n30904 = ~n31047 | ~n30934;
  assign n30898 = ~n30897;
  assign n30902 = ~n30899 & ~n30898;
  assign n30901 = n41095 & n30900;
  assign n31048 = ~n30902 & ~n30901;
  assign n30903 = ~n31048 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n30905 = ~n30904 | ~n30903;
  assign n30907 = ~n30906 & ~n30905;
  assign P3_U2909 = ~n30908 | ~n30907;
  assign n30910 = ~n30917 & ~n31038;
  assign n30909 = ~n31045 & ~n30918;
  assign n30916 = ~n30910 & ~n30909;
  assign n30914 = ~n30921 & ~n31040;
  assign n30912 = ~n31047 | ~n30922;
  assign n30911 = ~n31048 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n30913 = ~n30912 | ~n30911;
  assign n30915 = ~n30914 & ~n30913;
  assign P3_U2913 = ~n30916 | ~n30915;
  assign n30920 = ~n30917 & ~n30989;
  assign n30919 = ~n30918 & ~n30990;
  assign n30928 = ~n30920 & ~n30919;
  assign n30926 = ~n30921 & ~n30993;
  assign n30924 = ~n30994 | ~n30922;
  assign n30923 = ~n30995 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n30925 = ~n30924 | ~n30923;
  assign n30927 = ~n30926 & ~n30925;
  assign P3_U2977 = ~n30928 | ~n30927;
  assign n30932 = ~n30929 & ~n30989;
  assign n30931 = ~n30930 & ~n30993;
  assign n30940 = ~n30932 & ~n30931;
  assign n30938 = ~n30933 & ~n30990;
  assign n30936 = ~n30994 | ~n30934;
  assign n30935 = ~n30995 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n30937 = ~n30936 | ~n30935;
  assign n30939 = ~n30938 & ~n30937;
  assign P3_U2973 = ~n30940 | ~n30939;
  assign n30942 = ~n31014 & ~n30989;
  assign n30941 = ~n31015 & ~n30993;
  assign n30948 = ~n30942 & ~n30941;
  assign n30946 = ~n31018 & ~n30990;
  assign n30944 = ~n30994 | ~n31019;
  assign n30943 = ~n30995 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n30945 = ~n30944 | ~n30943;
  assign n30947 = ~n30946 & ~n30945;
  assign P3_U2976 = ~n30948 | ~n30947;
  assign n30950 = ~n31026 & ~n30989;
  assign n30949 = ~n31027 & ~n30993;
  assign n30956 = ~n30950 & ~n30949;
  assign n30954 = ~n31030 & ~n30990;
  assign n30952 = ~n30994 | ~n31031;
  assign n30951 = ~n30995 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n30953 = ~n30952 | ~n30951;
  assign n30955 = ~n30954 & ~n30953;
  assign P3_U2975 = ~n30956 | ~n30955;
  assign n30958 = ~n30966 & ~n31038;
  assign n30957 = ~n31045 & ~n30965;
  assign n30964 = ~n30958 & ~n30957;
  assign n30962 = ~n30969 & ~n31040;
  assign n30960 = ~n31047 | ~n30970;
  assign n30959 = ~n31048 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n30961 = ~n30960 | ~n30959;
  assign n30963 = ~n30962 & ~n30961;
  assign P3_U2914 = ~n30964 | ~n30963;
  assign n30968 = ~n30965 & ~n30990;
  assign n30967 = ~n30966 & ~n30989;
  assign n30976 = ~n30968 & ~n30967;
  assign n30974 = ~n30969 & ~n30993;
  assign n30972 = ~n30994 | ~n30970;
  assign n30971 = ~n30995 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n30973 = ~n30972 | ~n30971;
  assign n30975 = ~n30974 & ~n30973;
  assign P3_U2978 = ~n30976 | ~n30975;
  assign n30980 = ~n30977 & ~n31038;
  assign n30979 = ~n30978 & ~n31040;
  assign n30988 = ~n30980 & ~n30979;
  assign n30986 = ~n30981 & ~n31045;
  assign n30984 = ~n31047 | ~n30982;
  assign n30983 = ~n31048 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n30985 = ~n30984 | ~n30983;
  assign n30987 = ~n30986 & ~n30985;
  assign P3_U2908 = ~n30988 | ~n30987;
  assign n30992 = ~n31039 & ~n30989;
  assign n30991 = ~n31044 & ~n30990;
  assign n31001 = ~n30992 & ~n30991;
  assign n30999 = ~n31041 & ~n30993;
  assign n30997 = ~n30994 | ~n31046;
  assign n30996 = ~n30995 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n30998 = ~n30997 | ~n30996;
  assign n31000 = ~n30999 & ~n30998;
  assign P3_U2979 = ~n31001 | ~n31000;
  assign n31005 = ~n31002 & ~n31040;
  assign n31004 = ~n31003 & ~n31038;
  assign n31013 = ~n31005 & ~n31004;
  assign n31011 = ~n31045 & ~n31006;
  assign n31009 = ~n31047 | ~n31007;
  assign n31008 = ~n31048 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n31010 = ~n31009 | ~n31008;
  assign n31012 = ~n31011 & ~n31010;
  assign P3_U2910 = ~n31013 | ~n31012;
  assign n31017 = ~n31014 & ~n31038;
  assign n31016 = ~n31015 & ~n31040;
  assign n31025 = ~n31017 & ~n31016;
  assign n31023 = ~n31045 & ~n31018;
  assign n31021 = ~n31047 | ~n31019;
  assign n31020 = ~n31048 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n31022 = ~n31021 | ~n31020;
  assign n31024 = ~n31023 & ~n31022;
  assign P3_U2912 = ~n31025 | ~n31024;
  assign n31029 = ~n31026 & ~n31038;
  assign n31028 = ~n31027 & ~n31040;
  assign n31037 = ~n31029 & ~n31028;
  assign n31035 = ~n31045 & ~n31030;
  assign n31033 = ~n31047 | ~n31031;
  assign n31032 = ~n31048 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n31034 = ~n31033 | ~n31032;
  assign n31036 = ~n31035 & ~n31034;
  assign P3_U2911 = ~n31037 | ~n31036;
  assign n31043 = ~n31039 & ~n31038;
  assign n31042 = ~n31041 & ~n31040;
  assign n31054 = ~n31043 & ~n31042;
  assign n31052 = ~n31045 & ~n31044;
  assign n31050 = ~n31047 | ~n31046;
  assign n31049 = ~n31048 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n31051 = ~n31050 | ~n31049;
  assign n31053 = ~n31052 & ~n31051;
  assign P3_U2915 = ~n31054 | ~n31053;
  assign n44002 = n39508 & n31055;
  assign n31200 = ~n31057 | ~n31056;
  assign n31062 = ~n44002 & ~n31196;
  assign n31059 = ~n31058 & ~n32149;
  assign n31060 = ~n31525 | ~n31059;
  assign n31061 = ~P2_MEMORYFETCH_REG_SCAN_IN | ~n31060;
  assign P2_U2814 = ~n31062 | ~n31061;
  assign n31190 = ~n31189 & ~n31063;
  assign n31065 = ~BUF1_REG_7__SCAN_IN | ~n31190;
  assign n31064 = ~P1_DATAO_REG_7__SCAN_IN | ~n31189;
  assign n31067 = n31065 & n31064;
  assign n31066 = ~P2_DATAO_REG_7__SCAN_IN | ~n31193;
  assign U240 = ~n31067 | ~n31066;
  assign n31069 = ~BUF1_REG_24__SCAN_IN | ~n31190;
  assign n31068 = ~P1_DATAO_REG_24__SCAN_IN | ~n31189;
  assign n31071 = n31069 & n31068;
  assign n31070 = ~P2_DATAO_REG_24__SCAN_IN | ~n31193;
  assign U223 = ~n31071 | ~n31070;
  assign n31073 = ~BUF1_REG_0__SCAN_IN | ~n31190;
  assign n31072 = ~P1_DATAO_REG_0__SCAN_IN | ~n31189;
  assign n31075 = n31073 & n31072;
  assign n31074 = ~P2_DATAO_REG_0__SCAN_IN | ~n31193;
  assign U247 = ~n31075 | ~n31074;
  assign n31077 = ~BUF1_REG_18__SCAN_IN | ~n31190;
  assign n31076 = ~P1_DATAO_REG_18__SCAN_IN | ~n31189;
  assign n31079 = n31077 & n31076;
  assign n31078 = ~P2_DATAO_REG_18__SCAN_IN | ~n31193;
  assign U229 = ~n31079 | ~n31078;
  assign n31081 = ~BUF1_REG_3__SCAN_IN | ~n31190;
  assign n31080 = ~P1_DATAO_REG_3__SCAN_IN | ~n31189;
  assign n31083 = n31081 & n31080;
  assign n31082 = ~P2_DATAO_REG_3__SCAN_IN | ~n31193;
  assign U244 = ~n31083 | ~n31082;
  assign n31085 = ~BUF1_REG_6__SCAN_IN | ~n31190;
  assign n31084 = ~P1_DATAO_REG_6__SCAN_IN | ~n31189;
  assign n31087 = n31085 & n31084;
  assign n31086 = ~P2_DATAO_REG_6__SCAN_IN | ~n31193;
  assign U241 = ~n31087 | ~n31086;
  assign n31089 = ~BUF1_REG_20__SCAN_IN | ~n31190;
  assign n31088 = ~P1_DATAO_REG_20__SCAN_IN | ~n31189;
  assign n31091 = n31089 & n31088;
  assign n31090 = ~P2_DATAO_REG_20__SCAN_IN | ~n31193;
  assign U227 = ~n31091 | ~n31090;
  assign n31093 = ~BUF1_REG_29__SCAN_IN | ~n31190;
  assign n31092 = ~P1_DATAO_REG_29__SCAN_IN | ~n31189;
  assign n31095 = n31093 & n31092;
  assign n31094 = ~P2_DATAO_REG_29__SCAN_IN | ~n31193;
  assign U218 = ~n31095 | ~n31094;
  assign n31097 = ~BUF1_REG_27__SCAN_IN | ~n31190;
  assign n31096 = ~P1_DATAO_REG_27__SCAN_IN | ~n31189;
  assign n31099 = n31097 & n31096;
  assign n31098 = ~P2_DATAO_REG_27__SCAN_IN | ~n31193;
  assign U220 = ~n31099 | ~n31098;
  assign n31101 = ~BUF1_REG_4__SCAN_IN | ~n31190;
  assign n31100 = ~P1_DATAO_REG_4__SCAN_IN | ~n31189;
  assign n31103 = n31101 & n31100;
  assign n31102 = ~P2_DATAO_REG_4__SCAN_IN | ~n31193;
  assign U243 = ~n31103 | ~n31102;
  assign n31105 = ~BUF1_REG_16__SCAN_IN | ~n31190;
  assign n31104 = ~P1_DATAO_REG_16__SCAN_IN | ~n31189;
  assign n31107 = n31105 & n31104;
  assign n31106 = ~P2_DATAO_REG_16__SCAN_IN | ~n31193;
  assign U231 = ~n31107 | ~n31106;
  assign n31109 = ~BUF1_REG_15__SCAN_IN | ~n31190;
  assign n31108 = ~P1_DATAO_REG_15__SCAN_IN | ~n31189;
  assign n31111 = n31109 & n31108;
  assign n31110 = ~P2_DATAO_REG_15__SCAN_IN | ~n31193;
  assign U232 = ~n31111 | ~n31110;
  assign n31113 = ~BUF1_REG_25__SCAN_IN | ~n31190;
  assign n31112 = ~P1_DATAO_REG_25__SCAN_IN | ~n31189;
  assign n31115 = n31113 & n31112;
  assign n31114 = ~P2_DATAO_REG_25__SCAN_IN | ~n31193;
  assign U222 = ~n31115 | ~n31114;
  assign n31117 = ~BUF1_REG_13__SCAN_IN | ~n31190;
  assign n31116 = ~P1_DATAO_REG_13__SCAN_IN | ~n31189;
  assign n31119 = n31117 & n31116;
  assign n31118 = ~P2_DATAO_REG_13__SCAN_IN | ~n31193;
  assign U234 = ~n31119 | ~n31118;
  assign n31121 = ~BUF1_REG_9__SCAN_IN | ~n31190;
  assign n31120 = ~P1_DATAO_REG_9__SCAN_IN | ~n31189;
  assign n31123 = n31121 & n31120;
  assign n31122 = ~P2_DATAO_REG_9__SCAN_IN | ~n31193;
  assign U238 = ~n31123 | ~n31122;
  assign n31125 = ~BUF1_REG_22__SCAN_IN | ~n31190;
  assign n31124 = ~P1_DATAO_REG_22__SCAN_IN | ~n31189;
  assign n31127 = n31125 & n31124;
  assign n31126 = ~P2_DATAO_REG_22__SCAN_IN | ~n31193;
  assign U225 = ~n31127 | ~n31126;
  assign n31129 = ~BUF1_REG_8__SCAN_IN | ~n31190;
  assign n31128 = ~P1_DATAO_REG_8__SCAN_IN | ~n31189;
  assign n31131 = n31129 & n31128;
  assign n31130 = ~P2_DATAO_REG_8__SCAN_IN | ~n31193;
  assign U239 = ~n31131 | ~n31130;
  assign n31133 = ~BUF1_REG_2__SCAN_IN | ~n31190;
  assign n31132 = ~P1_DATAO_REG_2__SCAN_IN | ~n31189;
  assign n31135 = n31133 & n31132;
  assign n31134 = ~P2_DATAO_REG_2__SCAN_IN | ~n31193;
  assign U245 = ~n31135 | ~n31134;
  assign n31137 = ~BUF1_REG_17__SCAN_IN | ~n31190;
  assign n31136 = ~P1_DATAO_REG_17__SCAN_IN | ~n31189;
  assign n31139 = n31137 & n31136;
  assign n31138 = ~P2_DATAO_REG_17__SCAN_IN | ~n31193;
  assign U230 = ~n31139 | ~n31138;
  assign n31141 = ~BUF1_REG_30__SCAN_IN | ~n31190;
  assign n31140 = ~P1_DATAO_REG_30__SCAN_IN | ~n31189;
  assign n31143 = n31141 & n31140;
  assign n31142 = ~P2_DATAO_REG_30__SCAN_IN | ~n31193;
  assign U217 = ~n31143 | ~n31142;
  assign n31145 = ~BUF1_REG_28__SCAN_IN | ~n31190;
  assign n31144 = ~P1_DATAO_REG_28__SCAN_IN | ~n31189;
  assign n31147 = n31145 & n31144;
  assign n31146 = ~P2_DATAO_REG_28__SCAN_IN | ~n31193;
  assign U219 = ~n31147 | ~n31146;
  assign n31149 = ~BUF1_REG_1__SCAN_IN | ~n31190;
  assign n31148 = ~P1_DATAO_REG_1__SCAN_IN | ~n31189;
  assign n31151 = n31149 & n31148;
  assign n31150 = ~P2_DATAO_REG_1__SCAN_IN | ~n31193;
  assign U246 = ~n31151 | ~n31150;
  assign n31153 = ~BUF1_REG_14__SCAN_IN | ~n31190;
  assign n31152 = ~P1_DATAO_REG_14__SCAN_IN | ~n31189;
  assign n31155 = n31153 & n31152;
  assign n31154 = ~P2_DATAO_REG_14__SCAN_IN | ~n31193;
  assign U233 = ~n31155 | ~n31154;
  assign n31157 = ~BUF1_REG_21__SCAN_IN | ~n31190;
  assign n31156 = ~P1_DATAO_REG_21__SCAN_IN | ~n31189;
  assign n31159 = n31157 & n31156;
  assign n31158 = ~P2_DATAO_REG_21__SCAN_IN | ~n31193;
  assign U226 = ~n31159 | ~n31158;
  assign n31161 = ~P1_DATAO_REG_11__SCAN_IN | ~n31189;
  assign n31160 = ~BUF1_REG_11__SCAN_IN | ~n31190;
  assign n31163 = n31161 & n31160;
  assign n31162 = ~P2_DATAO_REG_11__SCAN_IN | ~n31193;
  assign U236 = ~n31163 | ~n31162;
  assign n31165 = ~P1_DATAO_REG_23__SCAN_IN | ~n31189;
  assign n31164 = ~BUF1_REG_23__SCAN_IN | ~n31190;
  assign n31167 = n31165 & n31164;
  assign n31166 = ~P2_DATAO_REG_23__SCAN_IN | ~n31193;
  assign U224 = ~n31167 | ~n31166;
  assign n31170 = ~n31168 & ~U212;
  assign n31169 = BUF1_REG_31__SCAN_IN & n31190;
  assign n31172 = ~n31170 & ~n31169;
  assign n31171 = ~P1_DATAO_REG_31__SCAN_IN | ~n31189;
  assign U216 = ~n31172 | ~n31171;
  assign n31174 = ~P1_DATAO_REG_10__SCAN_IN | ~n31189;
  assign n31173 = ~BUF1_REG_10__SCAN_IN | ~n31190;
  assign n31176 = n31174 & n31173;
  assign n31175 = ~P2_DATAO_REG_10__SCAN_IN | ~n31193;
  assign U237 = ~n31176 | ~n31175;
  assign n31178 = ~P1_DATAO_REG_5__SCAN_IN | ~n31189;
  assign n31177 = ~BUF1_REG_5__SCAN_IN | ~n31190;
  assign n31180 = n31178 & n31177;
  assign n31179 = ~P2_DATAO_REG_5__SCAN_IN | ~n31193;
  assign U242 = ~n31180 | ~n31179;
  assign n31182 = ~P1_DATAO_REG_12__SCAN_IN | ~n31189;
  assign n31181 = ~BUF1_REG_12__SCAN_IN | ~n31190;
  assign n31184 = n31182 & n31181;
  assign n31183 = ~P2_DATAO_REG_12__SCAN_IN | ~n31193;
  assign U235 = ~n31184 | ~n31183;
  assign n31186 = ~P1_DATAO_REG_26__SCAN_IN | ~n31189;
  assign n31185 = ~BUF1_REG_26__SCAN_IN | ~n31190;
  assign n31188 = n31186 & n31185;
  assign n31187 = ~P2_DATAO_REG_26__SCAN_IN | ~n31193;
  assign U221 = ~n31188 | ~n31187;
  assign n31192 = ~P1_DATAO_REG_19__SCAN_IN | ~n31189;
  assign n31191 = ~BUF1_REG_19__SCAN_IN | ~n31190;
  assign n31195 = n31192 & n31191;
  assign n31194 = ~P2_DATAO_REG_19__SCAN_IN | ~n31193;
  assign U228 = ~n31195 | ~n31194;
  assign n31197 = ~P2_EAX_REG_29__SCAN_IN;
  assign n31201 = ~n31817 & ~n31197;
  assign n31199 = ~BUF2_REG_13__SCAN_IN | ~n36558;
  assign n31198 = ~BUF1_REG_13__SCAN_IN | ~n36557;
  assign n43634 = n31199 & n31198;
  assign n31224 = ~n43634 & ~n31286;
  assign n31204 = ~n31201 & ~n31224;
  assign n31203 = ~n31353 | ~P2_UWORD_REG_13__SCAN_IN;
  assign P2_U2965 = ~n31204 | ~n31203;
  assign n31207 = n31344 & P2_EAX_REG_12__SCAN_IN;
  assign n31206 = ~BUF2_REG_12__SCAN_IN | ~n36558;
  assign n31205 = ~n36557 | ~BUF1_REG_12__SCAN_IN;
  assign n43111 = n31206 & n31205;
  assign n31253 = ~n43111 & ~n31286;
  assign n31209 = ~n31207 & ~n31253;
  assign n31208 = ~n31353 | ~P2_LWORD_REG_12__SCAN_IN;
  assign P2_U2979 = ~n31209 | ~n31208;
  assign n31211 = ~n31817 & ~n31210;
  assign n31229 = ~n32348 & ~n31286;
  assign n31213 = ~n31211 & ~n31229;
  assign n31212 = ~n31353 | ~P2_LWORD_REG_7__SCAN_IN;
  assign P2_U2974 = ~n31213 | ~n31212;
  assign n31215 = ~n31817 & ~n31214;
  assign n31248 = ~n36001 & ~n31286;
  assign n31217 = ~n31215 & ~n31248;
  assign n31216 = ~n31353 | ~P2_UWORD_REG_3__SCAN_IN;
  assign P2_U2955 = ~n31217 | ~n31216;
  assign n41758 = ~P2_EAX_REG_24__SCAN_IN;
  assign n31220 = ~n31817 & ~n41758;
  assign n31219 = ~BUF2_REG_8__SCAN_IN | ~n36558;
  assign n31218 = ~n36557 | ~BUF1_REG_8__SCAN_IN;
  assign n41757 = n31219 & n31218;
  assign n31233 = ~n41757 & ~n31286;
  assign n31222 = ~n31220 & ~n31233;
  assign n31221 = ~n31353 | ~P2_UWORD_REG_8__SCAN_IN;
  assign P2_U2960 = ~n31222 | ~n31221;
  assign n31225 = ~n31817 & ~n31223;
  assign n31227 = ~n31225 & ~n31224;
  assign n31226 = ~n31353 | ~P2_LWORD_REG_13__SCAN_IN;
  assign P2_U2980 = ~n31227 | ~n31226;
  assign n31230 = ~n31817 & ~n31228;
  assign n31232 = ~n31230 & ~n31229;
  assign n31231 = ~n31353 | ~P2_UWORD_REG_7__SCAN_IN;
  assign P2_U2959 = ~n31232 | ~n31231;
  assign n32260 = ~P2_EAX_REG_8__SCAN_IN;
  assign n31234 = ~n31817 & ~n32260;
  assign n31236 = ~n31234 & ~n31233;
  assign n31235 = ~n31353 | ~P2_LWORD_REG_8__SCAN_IN;
  assign P2_U2975 = ~n31236 | ~n31235;
  assign n31237 = ~P2_EAX_REG_22__SCAN_IN;
  assign n31240 = ~n31817 & ~n31237;
  assign n31239 = ~BUF2_REG_6__SCAN_IN | ~n36558;
  assign n31238 = ~n36557 | ~BUF1_REG_6__SCAN_IN;
  assign n40056 = ~n31239 | ~n31238;
  assign n32225 = ~n40056;
  assign n31262 = ~n32225 & ~n31286;
  assign n31242 = ~n31240 & ~n31262;
  assign n31241 = ~n31353 | ~P2_UWORD_REG_6__SCAN_IN;
  assign P2_U2958 = ~n31242 | ~n31241;
  assign n31245 = n31344 & P2_EAX_REG_14__SCAN_IN;
  assign n31244 = ~BUF2_REG_14__SCAN_IN | ~n36558;
  assign n31243 = ~BUF1_REG_14__SCAN_IN | ~n36557;
  assign n43696 = n31244 & n31243;
  assign n31258 = ~n43696 & ~n31286;
  assign n31247 = ~n31245 & ~n31258;
  assign n31246 = ~n31353 | ~P2_LWORD_REG_14__SCAN_IN;
  assign P2_U2981 = ~n31247 | ~n31246;
  assign n31249 = n31344 & P2_EAX_REG_3__SCAN_IN;
  assign n31251 = ~n31249 & ~n31248;
  assign n31250 = ~n31353 | ~P2_LWORD_REG_3__SCAN_IN;
  assign P2_U2970 = ~n31251 | ~n31250;
  assign n31254 = ~n31817 & ~n31252;
  assign n31256 = ~n31254 & ~n31253;
  assign n31255 = ~n31353 | ~P2_UWORD_REG_12__SCAN_IN;
  assign P2_U2964 = ~n31256 | ~n31255;
  assign n31257 = ~P2_EAX_REG_30__SCAN_IN;
  assign n31259 = ~n31817 & ~n31257;
  assign n31261 = ~n31259 & ~n31258;
  assign n31260 = ~n31353 | ~P2_UWORD_REG_14__SCAN_IN;
  assign P2_U2966 = ~n31261 | ~n31260;
  assign n31263 = ~n31817 & ~n25671;
  assign n31265 = ~n31263 & ~n31262;
  assign n31264 = ~n31353 | ~P2_LWORD_REG_6__SCAN_IN;
  assign P2_U2973 = ~n31265 | ~n31264;
  assign n31267 = ~BUF2_REG_15__SCAN_IN | ~n36558;
  assign n31266 = ~n36557 | ~BUF1_REG_15__SCAN_IN;
  assign n35317 = n31267 & n31266;
  assign n31270 = ~n35317 & ~n31286;
  assign n31269 = ~n31817 & ~n31268;
  assign n31272 = ~n31270 & ~n31269;
  assign n31271 = ~P2_LWORD_REG_15__SCAN_IN | ~n31353;
  assign P2_U2982 = ~n31272 | ~n31271;
  assign n31275 = ~n31717 & ~n31442;
  assign n31274 = ~P1_MEMORYFETCH_REG_SCAN_IN | ~n31273;
  assign P1_U2801 = ~n31275 | ~n31274;
  assign n31278 = ~n31909 | ~n35466;
  assign n31277 = ~n31276 | ~n31898;
  assign n31378 = n31278 & n31277;
  assign n31279 = ~n31378 | ~n44102;
  assign n31281 = ~n31279 | ~P1_CODEFETCH_REG_SCAN_IN;
  assign n31280 = ~n44099 | ~n43722;
  assign P1_U2803 = ~n31281 | ~n31280;
  assign n31283 = ~P2_LWORD_REG_5__SCAN_IN | ~n31353;
  assign n31282 = ~n31344 | ~P2_EAX_REG_5__SCAN_IN;
  assign n31287 = n31283 & n31282;
  assign n31285 = ~BUF2_REG_5__SCAN_IN | ~n36558;
  assign n31284 = ~n36557 | ~BUF1_REG_5__SCAN_IN;
  assign n39675 = ~n31285 | ~n31284;
  assign n31326 = ~n39675 | ~n31322;
  assign P2_U2972 = ~n31287 | ~n31326;
  assign n31289 = ~P2_UWORD_REG_11__SCAN_IN | ~n31353;
  assign n31288 = ~n31344 | ~P2_EAX_REG_27__SCAN_IN;
  assign n31292 = n31289 & n31288;
  assign n31291 = ~BUF2_REG_11__SCAN_IN | ~n36558;
  assign n31290 = ~n36557 | ~BUF1_REG_11__SCAN_IN;
  assign n42803 = ~n31291 | ~n31290;
  assign n31351 = ~n42803 | ~n31322;
  assign P2_U2963 = ~n31292 | ~n31351;
  assign n31294 = ~P2_LWORD_REG_0__SCAN_IN | ~n31353;
  assign n31293 = ~n31344 | ~P2_EAX_REG_0__SCAN_IN;
  assign n31297 = n31294 & n31293;
  assign n31296 = ~BUF2_REG_0__SCAN_IN | ~n36558;
  assign n31295 = ~n36557 | ~BUF1_REG_0__SCAN_IN;
  assign n37112 = ~n31296 | ~n31295;
  assign n31342 = ~n37112 | ~n31322;
  assign P2_U2967 = ~n31297 | ~n31342;
  assign n31299 = ~P2_UWORD_REG_9__SCAN_IN | ~n31353;
  assign n31298 = ~n31344 | ~P2_EAX_REG_25__SCAN_IN;
  assign n31302 = n31299 & n31298;
  assign n31301 = ~BUF2_REG_9__SCAN_IN | ~n36558;
  assign n31300 = ~n36557 | ~BUF1_REG_9__SCAN_IN;
  assign n41659 = ~n31301 | ~n31300;
  assign n31356 = ~n41659 | ~n31322;
  assign P2_U2961 = ~n31302 | ~n31356;
  assign n31304 = ~P2_LWORD_REG_2__SCAN_IN | ~n31353;
  assign n31303 = ~n31344 | ~P2_EAX_REG_2__SCAN_IN;
  assign n31307 = n31304 & n31303;
  assign n31306 = ~BUF2_REG_2__SCAN_IN | ~n36558;
  assign n31305 = ~n36557 | ~BUF1_REG_2__SCAN_IN;
  assign n38018 = ~n31306 | ~n31305;
  assign n31330 = ~n38018 | ~n31322;
  assign P2_U2969 = ~n31307 | ~n31330;
  assign n31309 = ~P2_LWORD_REG_10__SCAN_IN | ~n31353;
  assign n31308 = ~n31344 | ~P2_EAX_REG_10__SCAN_IN;
  assign n31312 = n31309 & n31308;
  assign n31311 = ~BUF2_REG_10__SCAN_IN | ~n36558;
  assign n31310 = ~n36557 | ~BUF1_REG_10__SCAN_IN;
  assign n41831 = ~n31311 | ~n31310;
  assign n31334 = ~n41831 | ~n31322;
  assign P2_U2977 = ~n31312 | ~n31334;
  assign n31314 = ~P2_LWORD_REG_4__SCAN_IN | ~n31353;
  assign n31313 = ~n31344 | ~P2_EAX_REG_4__SCAN_IN;
  assign n31317 = n31314 & n31313;
  assign n31316 = ~BUF2_REG_4__SCAN_IN | ~n36558;
  assign n31315 = ~n36557 | ~BUF1_REG_4__SCAN_IN;
  assign n38972 = ~n31316 | ~n31315;
  assign n31338 = ~n38972 | ~n31322;
  assign P2_U2971 = ~n31317 | ~n31338;
  assign n31319 = ~P2_LWORD_REG_1__SCAN_IN | ~n31353;
  assign n31318 = ~n31344 | ~P2_EAX_REG_1__SCAN_IN;
  assign n31323 = n31319 & n31318;
  assign n31321 = ~BUF2_REG_1__SCAN_IN | ~n36558;
  assign n31320 = ~n36557 | ~BUF1_REG_1__SCAN_IN;
  assign n37434 = ~n31321 | ~n31320;
  assign n31347 = ~n37434 | ~n31322;
  assign P2_U2968 = ~n31323 | ~n31347;
  assign n31325 = ~n31344 | ~P2_EAX_REG_21__SCAN_IN;
  assign n31324 = ~P2_UWORD_REG_5__SCAN_IN | ~n31353;
  assign n31327 = n31325 & n31324;
  assign P2_U2957 = ~n31327 | ~n31326;
  assign n31329 = ~n31344 | ~P2_EAX_REG_18__SCAN_IN;
  assign n31328 = ~P2_UWORD_REG_2__SCAN_IN | ~n31353;
  assign n31331 = n31329 & n31328;
  assign P2_U2954 = ~n31331 | ~n31330;
  assign n31333 = ~n31344 | ~P2_EAX_REG_26__SCAN_IN;
  assign n31332 = ~P2_UWORD_REG_10__SCAN_IN | ~n31353;
  assign n31335 = n31333 & n31332;
  assign P2_U2962 = ~n31335 | ~n31334;
  assign n31337 = ~n31344 | ~P2_EAX_REG_20__SCAN_IN;
  assign n31336 = ~P2_UWORD_REG_4__SCAN_IN | ~n31353;
  assign n31339 = n31337 & n31336;
  assign P2_U2956 = ~n31339 | ~n31338;
  assign n31341 = ~n31344 | ~P2_EAX_REG_16__SCAN_IN;
  assign n31340 = ~P2_UWORD_REG_0__SCAN_IN | ~n31353;
  assign n31343 = n31341 & n31340;
  assign P2_U2952 = ~n31343 | ~n31342;
  assign n31346 = ~n31344 | ~P2_EAX_REG_17__SCAN_IN;
  assign n31345 = ~P2_UWORD_REG_1__SCAN_IN | ~n31353;
  assign n31348 = n31346 & n31345;
  assign P2_U2953 = ~n31348 | ~n31347;
  assign n31350 = ~n31817 & ~n25738;
  assign n31349 = P2_LWORD_REG_11__SCAN_IN & n31353;
  assign n31352 = ~n31350 & ~n31349;
  assign P2_U2978 = ~n31352 | ~n31351;
  assign n31355 = ~n31817 & ~n25724;
  assign n31354 = P2_LWORD_REG_9__SCAN_IN & n31353;
  assign n31357 = ~n31355 & ~n31354;
  assign P2_U2976 = ~n31357 | ~n31356;
  assign n34517 = ~n31358;
  assign n44028 = ~n31361 & ~n31360;
  assign P1_U2905 = n44092 & P1_DATAO_REG_31__SCAN_IN;
  assign n31363 = ~P1_EAX_REG_11__SCAN_IN | ~n44028;
  assign n31362 = ~n44093 | ~P1_LWORD_REG_11__SCAN_IN;
  assign n31365 = n31363 & n31362;
  assign n31364 = ~n44092 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P1_U2925 = ~n31365 | ~n31364;
  assign n31367 = ~n44093 | ~P1_LWORD_REG_13__SCAN_IN;
  assign n31366 = ~P1_EAX_REG_13__SCAN_IN | ~n44028;
  assign n31369 = n31367 & n31366;
  assign n31368 = ~n44092 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P1_U2923 = ~n31369 | ~n31368;
  assign n31373 = n31370 | n41384;
  assign n31826 = ~n31671 & ~n41374;
  assign n31532 = n31371 | n31805;
  assign n32844 = ~n31826 | ~n31670;
  assign n31372 = ~P3_CODEFETCH_REG_SCAN_IN | ~n32844;
  assign P3_U2634 = ~n31373 | ~n31372;
  assign n31375 = ~n31477 | ~n31374;
  assign n31481 = ~n35474 | ~n31374;
  assign n31376 = ~n31375 | ~n31481;
  assign n31377 = n31376 | n44100;
  assign n34496 = ~n31378 | ~n31377;
  assign n31446 = ~n34496 | ~n44102;
  assign n31379 = ~P1_FLUSH_REG_SCAN_IN | ~n31446;
  assign P1_U2806 = ~n43358 | ~n31379;
  assign n31381 = ~n44092 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n31380 = ~n44093 | ~P1_UWORD_REG_0__SCAN_IN;
  assign n31384 = n31381 & n31380;
  assign n31383 = ~n31439 | ~P1_EAX_REG_16__SCAN_IN;
  assign P1_U2920 = ~n31384 | ~n31383;
  assign n31386 = ~n44092 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n31385 = ~n44093 | ~P1_UWORD_REG_7__SCAN_IN;
  assign n31388 = n31386 & n31385;
  assign n31387 = ~n31439 | ~P1_EAX_REG_23__SCAN_IN;
  assign P1_U2913 = ~n31388 | ~n31387;
  assign n31390 = ~n44092 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n31389 = ~n44093 | ~P1_UWORD_REG_10__SCAN_IN;
  assign n31392 = n31390 & n31389;
  assign n31391 = ~n31439 | ~P1_EAX_REG_26__SCAN_IN;
  assign P1_U2910 = ~n31392 | ~n31391;
  assign n31394 = ~n44092 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n31393 = ~n44093 | ~P1_UWORD_REG_2__SCAN_IN;
  assign n31396 = n31394 & n31393;
  assign n31395 = ~n31439 | ~P1_EAX_REG_18__SCAN_IN;
  assign P1_U2918 = ~n31396 | ~n31395;
  assign n31398 = ~n44092 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n31397 = ~n44093 | ~P1_UWORD_REG_12__SCAN_IN;
  assign n31400 = n31398 & n31397;
  assign n31399 = ~n31439 | ~P1_EAX_REG_28__SCAN_IN;
  assign P1_U2908 = ~n31400 | ~n31399;
  assign n31402 = ~n44092 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n31401 = ~n44093 | ~P1_UWORD_REG_8__SCAN_IN;
  assign n31404 = n31402 & n31401;
  assign n31403 = ~n31439 | ~P1_EAX_REG_24__SCAN_IN;
  assign P1_U2912 = ~n31404 | ~n31403;
  assign n31406 = ~n44092 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n31405 = ~n44093 | ~P1_UWORD_REG_11__SCAN_IN;
  assign n31408 = n31406 & n31405;
  assign n31407 = ~n31439 | ~P1_EAX_REG_27__SCAN_IN;
  assign P1_U2909 = ~n31408 | ~n31407;
  assign n31410 = ~n44092 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n31409 = ~n44093 | ~P1_UWORD_REG_9__SCAN_IN;
  assign n31412 = n31410 & n31409;
  assign n31411 = ~n31439 | ~P1_EAX_REG_25__SCAN_IN;
  assign P1_U2911 = ~n31412 | ~n31411;
  assign n31414 = ~n44092 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n31413 = ~n44093 | ~P1_UWORD_REG_1__SCAN_IN;
  assign n31416 = n31414 & n31413;
  assign n31415 = ~n31439 | ~P1_EAX_REG_17__SCAN_IN;
  assign P1_U2919 = ~n31416 | ~n31415;
  assign n31418 = ~n44092 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n31417 = ~n44093 | ~P1_UWORD_REG_14__SCAN_IN;
  assign n31420 = n31418 & n31417;
  assign n31419 = ~n31439 | ~P1_EAX_REG_30__SCAN_IN;
  assign P1_U2906 = ~n31420 | ~n31419;
  assign n31422 = ~n44093 | ~P1_UWORD_REG_6__SCAN_IN;
  assign n31421 = ~n44092 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n31424 = n31422 & n31421;
  assign n31423 = ~n31439 | ~P1_EAX_REG_22__SCAN_IN;
  assign P1_U2914 = ~n31424 | ~n31423;
  assign n31426 = ~n44093 | ~P1_UWORD_REG_13__SCAN_IN;
  assign n31425 = ~n44092 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n31428 = n31426 & n31425;
  assign n31427 = ~n31439 | ~P1_EAX_REG_29__SCAN_IN;
  assign P1_U2907 = ~n31428 | ~n31427;
  assign n31430 = ~n44093 | ~P1_UWORD_REG_4__SCAN_IN;
  assign n31429 = ~n44092 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n31432 = n31430 & n31429;
  assign n31431 = ~n31439 | ~P1_EAX_REG_20__SCAN_IN;
  assign P1_U2916 = ~n31432 | ~n31431;
  assign n31434 = ~n44093 | ~P1_UWORD_REG_3__SCAN_IN;
  assign n31433 = ~n44092 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n31436 = n31434 & n31433;
  assign n31435 = ~n31439 | ~P1_EAX_REG_19__SCAN_IN;
  assign P1_U2917 = ~n31436 | ~n31435;
  assign n31438 = ~n44093 | ~P1_UWORD_REG_5__SCAN_IN;
  assign n31437 = ~n44092 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n31441 = n31438 & n31437;
  assign n31440 = ~n31439 | ~P1_EAX_REG_21__SCAN_IN;
  assign P1_U2915 = ~n31441 | ~n31440;
  assign n32081 = ~n31477 & ~n35474;
  assign n31445 = ~n35473 | ~n32081;
  assign n31443 = n31442 | P1_READREQUEST_REG_SCAN_IN;
  assign n31444 = ~n35465 | ~n31443;
  assign P1_U3487 = ~n31445 | ~n31444;
  assign n31461 = ~P1_MORE_REG_SCAN_IN | ~n31446;
  assign n31459 = ~n31446;
  assign n31457 = ~n31909 & ~n31447;
  assign n34509 = ~n32337;
  assign n31455 = n31448 | n34509;
  assign n31450 = ~n31449;
  assign n31452 = ~n31451 & ~n31450;
  assign n31453 = ~n31452 | ~n32080;
  assign n31454 = ~n31453 | ~n31909;
  assign n31456 = ~n31455 | ~n31454;
  assign n31458 = ~n31457 & ~n31456;
  assign n34499 = ~n31458 & ~n39892;
  assign n31460 = ~n31459 | ~n34499;
  assign P1_U3484 = ~n31461 | ~n31460;
  assign n31465 = ~n32966 | ~n32844;
  assign n31463 = ~n31465 & ~P3_MEMORYFETCH_REG_SCAN_IN;
  assign n31462 = ~n32860 & ~n32844;
  assign P3_U3299 = ~n31463 & ~n31462;
  assign n31464 = ~n31511;
  assign n31467 = ~n32844 & ~n31464;
  assign n31466 = ~n31465 & ~P3_READREQUEST_REG_SCAN_IN;
  assign P3_U3298 = ~n31467 & ~n31466;
  assign n31471 = ~n31468;
  assign n31470 = ~n34518 | ~n31469;
  assign n31472 = ~n31471 | ~n31470;
  assign n31474 = ~n35473 & ~n31472;
  assign n31486 = ~P1_REQUESTPENDING_REG_SCAN_IN | ~n31474;
  assign n31473 = ~n35630;
  assign n31475 = ~n31473 & ~P1_STATE2_REG_0__SCAN_IN;
  assign n31484 = ~n31475 & ~n31474;
  assign n31476 = ~n34515 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n31479 = ~n31477 | ~n31476;
  assign n31480 = ~n31479 | ~n31478;
  assign n31482 = ~n43722 & ~n31480;
  assign n31483 = ~n31482 | ~n31481;
  assign n31485 = ~n31484 | ~n31483;
  assign P1_U3485 = ~n31486 | ~n31485;
  assign n35709 = ~P2_STATE2_REG_0__SCAN_IN & ~n35802;
  assign n31490 = ~n35709 | ~n31487;
  assign n35708 = ~n31488 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n31489 = ~n35708 | ~n39522;
  assign n31491 = ~n31490 | ~n31489;
  assign n31504 = ~n44003 & ~n31491;
  assign n31503 = ~n31504;
  assign n31492 = ~n38321 & ~n31819;
  assign n31497 = ~n31493 & ~n31492;
  assign n31494 = ~n35802 & ~n39511;
  assign n31496 = ~n31495 & ~n31494;
  assign n31501 = ~n31497 & ~n31496;
  assign n31499 = ~n31498 & ~n43061;
  assign n31500 = ~n31499 | ~n31819;
  assign n31502 = ~n31501 | ~n31500;
  assign n31506 = ~n31503 | ~n31502;
  assign n31505 = ~n31504 | ~P2_REQUESTPENDING_REG_SCAN_IN;
  assign P2_U3610 = ~n31506 | ~n31505;
  assign n31510 = ~n35442 & ~n42025;
  assign n31508 = ~n32190 | ~n31667;
  assign n31509 = ~n32844 | ~n31508;
  assign n31519 = ~n31510 & ~n31509;
  assign n31518 = ~n31519;
  assign n31513 = ~P3_STATEBS16_REG_SCAN_IN & ~n32868;
  assign n31512 = ~n32857 | ~n31667;
  assign n31514 = ~n31513 & ~n31512;
  assign n31515 = ~P3_STATE2_REG_2__SCAN_IN | ~n31514;
  assign n31516 = ~P3_STATE2_REG_0__SCAN_IN | ~n31515;
  assign n31517 = ~n42012 | ~n31516;
  assign n31521 = ~n31518 | ~n31517;
  assign n31520 = ~n31519 | ~P3_REQUESTPENDING_REG_SCAN_IN;
  assign P3_U3296 = ~n31521 | ~n31520;
  assign n31531 = ~P2_STATE2_REG_0__SCAN_IN | ~n44002;
  assign n31523 = ~n31522;
  assign n31528 = ~n31524 | ~n31523;
  assign n31526 = ~n31771 | ~n31525;
  assign n31527 = ~n31526 | ~n31766;
  assign n31711 = n31528 & n31527;
  assign n31529 = ~n31711 | ~n35805;
  assign n31530 = ~P2_CODEFETCH_REG_SCAN_IN | ~n31529;
  assign P2_U2816 = ~n31531 | ~n31530;
  assign n35697 = ~P3_EAX_REG_15__SCAN_IN;
  assign n31537 = ~n35697 & ~n31659;
  assign n31535 = ~BUF2_REG_15__SCAN_IN;
  assign n31533 = ~n31667 & ~n33487;
  assign n31621 = n31662 | n33487;
  assign n31536 = ~n31535 & ~n31621;
  assign n31539 = ~n31537 & ~n31536;
  assign n31538 = ~P3_LWORD_REG_15__SCAN_IN | ~n31662;
  assign P3_U2798 = ~n31539 | ~n31538;
  assign n32207 = ~BUF2_REG_4__SCAN_IN;
  assign n31605 = ~n32207 & ~n31621;
  assign n32204 = ~P3_EAX_REG_4__SCAN_IN;
  assign n31540 = ~n32204 & ~n31659;
  assign n31542 = ~n31605 & ~n31540;
  assign n31541 = ~P3_LWORD_REG_4__SCAN_IN | ~n31662;
  assign P3_U2787 = ~n31542 | ~n31541;
  assign n31543 = ~BUF2_REG_2__SCAN_IN;
  assign n31661 = ~n31543 & ~n31621;
  assign n31544 = ~P3_EAX_REG_2__SCAN_IN;
  assign n31545 = ~n31544 & ~n31659;
  assign n31547 = ~n31661 & ~n31545;
  assign n31546 = ~P3_LWORD_REG_2__SCAN_IN | ~n31662;
  assign P3_U2785 = ~n31547 | ~n31546;
  assign n31548 = ~BUF2_REG_6__SCAN_IN;
  assign n31643 = ~n31548 & ~n31621;
  assign n31549 = ~P3_EAX_REG_6__SCAN_IN;
  assign n31550 = ~n31549 & ~n31659;
  assign n31552 = ~n31643 & ~n31550;
  assign n31551 = ~P3_LWORD_REG_6__SCAN_IN | ~n31662;
  assign P3_U2789 = ~n31552 | ~n31551;
  assign n31553 = ~BUF2_REG_13__SCAN_IN;
  assign n31592 = ~n31553 & ~n31621;
  assign n31554 = ~P3_EAX_REG_13__SCAN_IN;
  assign n31555 = ~n31554 & ~n31659;
  assign n31557 = ~n31592 & ~n31555;
  assign n31556 = ~P3_LWORD_REG_13__SCAN_IN | ~n31662;
  assign P3_U2796 = ~n31557 | ~n31556;
  assign n31558 = ~BUF2_REG_0__SCAN_IN;
  assign n31635 = ~n31558 & ~n31621;
  assign n32280 = ~P3_EAX_REG_0__SCAN_IN;
  assign n31559 = ~n32280 & ~n31659;
  assign n31561 = ~n31635 & ~n31559;
  assign n31560 = ~P3_LWORD_REG_0__SCAN_IN | ~n31662;
  assign P3_U2783 = ~n31561 | ~n31560;
  assign n34351 = ~BUF2_REG_11__SCAN_IN;
  assign n31601 = ~n34351 & ~n31621;
  assign n34356 = ~P3_EAX_REG_11__SCAN_IN;
  assign n31562 = ~n34356 & ~n31659;
  assign n31564 = ~n31601 & ~n31562;
  assign n31563 = ~P3_LWORD_REG_11__SCAN_IN | ~n31662;
  assign P3_U2794 = ~n31564 | ~n31563;
  assign n33222 = ~BUF2_REG_10__SCAN_IN;
  assign n31614 = ~n33222 & ~n31621;
  assign n31565 = ~P3_EAX_REG_10__SCAN_IN;
  assign n31566 = ~n31565 & ~n31659;
  assign n31568 = ~n31614 & ~n31566;
  assign n31567 = ~P3_LWORD_REG_10__SCAN_IN | ~n31662;
  assign P3_U2793 = ~n31568 | ~n31567;
  assign n32283 = ~BUF2_REG_1__SCAN_IN;
  assign n31651 = ~n32283 & ~n31621;
  assign n32279 = ~P3_EAX_REG_1__SCAN_IN;
  assign n31569 = ~n32279 & ~n31659;
  assign n31571 = ~n31651 & ~n31569;
  assign n31570 = ~P3_LWORD_REG_1__SCAN_IN | ~n31662;
  assign P3_U2784 = ~n31571 | ~n31570;
  assign n32323 = ~BUF2_REG_8__SCAN_IN;
  assign n31584 = ~n32323 & ~n31621;
  assign n43952 = ~P3_EAX_REG_24__SCAN_IN;
  assign n31572 = ~n43952 & ~n31659;
  assign n31574 = ~n31584 & ~n31572;
  assign n31573 = ~P3_UWORD_REG_8__SCAN_IN | ~n31662;
  assign P3_U2776 = ~n31574 | ~n31573;
  assign n31575 = ~BUF2_REG_14__SCAN_IN;
  assign n31626 = ~n31575 & ~n31621;
  assign n36280 = ~P3_EAX_REG_30__SCAN_IN;
  assign n31576 = ~n36280 & ~n31659;
  assign n31578 = ~n31626 & ~n31576;
  assign n31577 = ~P3_UWORD_REG_14__SCAN_IN | ~n31662;
  assign P3_U2782 = ~n31578 | ~n31577;
  assign n32834 = ~BUF2_REG_9__SCAN_IN;
  assign n31630 = ~n32834 & ~n31621;
  assign n32839 = ~P3_EAX_REG_9__SCAN_IN;
  assign n31579 = ~n32839 & ~n31659;
  assign n31581 = ~n31630 & ~n31579;
  assign n31580 = ~P3_LWORD_REG_9__SCAN_IN | ~n31662;
  assign P3_U2792 = ~n31581 | ~n31580;
  assign n31582 = ~P3_EAX_REG_8__SCAN_IN;
  assign n31583 = ~n31582 & ~n31659;
  assign n31586 = ~n31584 & ~n31583;
  assign n31585 = ~P3_LWORD_REG_8__SCAN_IN | ~n31662;
  assign P3_U2791 = ~n31586 | ~n31585;
  assign n31597 = ~n34844 & ~n31621;
  assign n31587 = ~P3_EAX_REG_12__SCAN_IN;
  assign n31588 = ~n31587 & ~n31659;
  assign n31590 = ~n31597 & ~n31588;
  assign n31589 = ~P3_LWORD_REG_12__SCAN_IN | ~n31662;
  assign P3_U2795 = ~n31590 | ~n31589;
  assign n43937 = ~P3_EAX_REG_29__SCAN_IN;
  assign n31591 = ~n43937 & ~n31659;
  assign n31594 = ~n31592 & ~n31591;
  assign n31593 = ~P3_UWORD_REG_13__SCAN_IN | ~n31662;
  assign P3_U2781 = ~n31594 | ~n31593;
  assign n31595 = ~P3_EAX_REG_28__SCAN_IN;
  assign n31596 = ~n31595 & ~n31659;
  assign n31599 = ~n31597 & ~n31596;
  assign n31598 = ~P3_UWORD_REG_12__SCAN_IN | ~n31662;
  assign P3_U2780 = ~n31599 | ~n31598;
  assign n43942 = ~P3_EAX_REG_27__SCAN_IN;
  assign n31600 = ~n43942 & ~n31659;
  assign n31603 = ~n31601 & ~n31600;
  assign n31602 = ~P3_UWORD_REG_11__SCAN_IN | ~n31662;
  assign P3_U2779 = ~n31603 | ~n31602;
  assign n43972 = ~P3_EAX_REG_20__SCAN_IN;
  assign n31604 = ~n43972 & ~n31659;
  assign n31607 = ~n31605 & ~n31604;
  assign n31606 = ~P3_UWORD_REG_4__SCAN_IN | ~n31662;
  assign P3_U2772 = ~n31607 | ~n31606;
  assign n31608 = ~BUF2_REG_5__SCAN_IN;
  assign n31647 = ~n31608 & ~n31621;
  assign n31609 = ~n32499 & ~n31659;
  assign n31611 = ~n31647 & ~n31609;
  assign n31610 = ~P3_LWORD_REG_5__SCAN_IN | ~n31662;
  assign P3_U2788 = ~n31611 | ~n31610;
  assign n31612 = ~P3_EAX_REG_26__SCAN_IN;
  assign n31613 = ~n31612 & ~n31659;
  assign n31616 = ~n31614 & ~n31613;
  assign n31615 = ~P3_UWORD_REG_10__SCAN_IN | ~n31662;
  assign P3_U2778 = ~n31616 | ~n31615;
  assign n31617 = ~BUF2_REG_3__SCAN_IN;
  assign n31656 = ~n31617 & ~n31621;
  assign n32815 = ~P3_EAX_REG_3__SCAN_IN;
  assign n31618 = ~n32815 & ~n31659;
  assign n31620 = ~n31656 & ~n31618;
  assign n31619 = ~P3_LWORD_REG_3__SCAN_IN | ~n31662;
  assign P3_U2786 = ~n31620 | ~n31619;
  assign n32353 = ~BUF2_REG_7__SCAN_IN;
  assign n31639 = ~n32353 & ~n31621;
  assign n32328 = ~P3_EAX_REG_7__SCAN_IN;
  assign n31622 = ~n32328 & ~n31659;
  assign n31624 = ~n31639 & ~n31622;
  assign n31623 = ~P3_LWORD_REG_7__SCAN_IN | ~n31662;
  assign P3_U2790 = ~n31624 | ~n31623;
  assign n34969 = ~P3_EAX_REG_14__SCAN_IN;
  assign n31625 = ~n34969 & ~n31659;
  assign n31628 = ~n31626 & ~n31625;
  assign n31627 = ~P3_LWORD_REG_14__SCAN_IN | ~n31662;
  assign P3_U2797 = ~n31628 | ~n31627;
  assign n43947 = ~P3_EAX_REG_25__SCAN_IN;
  assign n31629 = ~n43947 & ~n31659;
  assign n31632 = ~n31630 & ~n31629;
  assign n31631 = ~P3_UWORD_REG_9__SCAN_IN | ~n31662;
  assign P3_U2777 = ~n31632 | ~n31631;
  assign n31634 = ~n31633 & ~n31659;
  assign n31637 = ~n31635 & ~n31634;
  assign n31636 = ~P3_UWORD_REG_0__SCAN_IN | ~n31662;
  assign P3_U2768 = ~n31637 | ~n31636;
  assign n43957 = ~P3_EAX_REG_23__SCAN_IN;
  assign n31638 = ~n43957 & ~n31659;
  assign n31641 = ~n31639 & ~n31638;
  assign n31640 = ~P3_UWORD_REG_7__SCAN_IN | ~n31662;
  assign P3_U2775 = ~n31641 | ~n31640;
  assign n43962 = ~P3_EAX_REG_22__SCAN_IN;
  assign n31642 = ~n43962 & ~n31659;
  assign n31645 = ~n31643 & ~n31642;
  assign n31644 = ~P3_UWORD_REG_6__SCAN_IN | ~n31662;
  assign P3_U2774 = ~n31645 | ~n31644;
  assign n31646 = ~n43967 & ~n31659;
  assign n31649 = ~n31647 & ~n31646;
  assign n31648 = ~P3_UWORD_REG_5__SCAN_IN | ~n31662;
  assign P3_U2773 = ~n31649 | ~n31648;
  assign n43983 = ~P3_EAX_REG_17__SCAN_IN;
  assign n31650 = ~n43983 & ~n31659;
  assign n31653 = ~n31651 & ~n31650;
  assign n31652 = ~P3_UWORD_REG_1__SCAN_IN | ~n31662;
  assign P3_U2769 = ~n31653 | ~n31652;
  assign n31654 = ~P3_EAX_REG_19__SCAN_IN;
  assign n31655 = ~n31654 & ~n31659;
  assign n31658 = ~n31656 & ~n31655;
  assign n31657 = ~P3_UWORD_REG_3__SCAN_IN | ~n31662;
  assign P3_U2771 = ~n31658 | ~n31657;
  assign n43977 = ~P3_EAX_REG_18__SCAN_IN;
  assign n31660 = ~n43977 & ~n31659;
  assign n31664 = ~n31661 & ~n31660;
  assign n31663 = ~P3_UWORD_REG_2__SCAN_IN | ~n31662;
  assign P3_U2770 = ~n31664 | ~n31663;
  assign n31668 = ~n31667 | ~n31666;
  assign n41359 = ~n32200 | ~n31668;
  assign n31791 = ~n42025 | ~n41359;
  assign n31678 = ~P3_MORE_REG_SCAN_IN | ~n31791;
  assign n31676 = ~n31791;
  assign n31669 = ~n40442 | ~n41235;
  assign n31675 = ~n31669 | ~n31808;
  assign n31672 = ~n31671 | ~n31670;
  assign n31673 = ~n31672 | ~n40202;
  assign n31674 = ~n31673 | ~n31788;
  assign n31677 = ~n31676 | ~n41365;
  assign P3_U3295 = ~n31678 | ~n31677;
  assign n31680 = ~n31679 | ~n40693;
  assign n31693 = ~n31680 | ~P1_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n31683 = ~n31681;
  assign n31685 = ~n31683 & ~n31682;
  assign n35468 = ~n31685 & ~n31684;
  assign n31691 = ~n35468 & ~n43729;
  assign n31695 = ~n43033 & ~n31686;
  assign n31689 = ~n31695;
  assign n31702 = ~n31687 ^ n32552;
  assign n31688 = ~n43707 | ~n31702;
  assign n31690 = ~n31689 | ~n31688;
  assign n31692 = ~n31691 & ~n31690;
  assign P1_U2999 = ~n31693 | ~n31692;
  assign n34285 = n32532 & n42922;
  assign n31701 = ~n34285 & ~n32552;
  assign n31694 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN & ~n42927;
  assign n31699 = ~n31695 & ~n31694;
  assign n31696 = ~n40080 & ~P1_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n35470 = ~n31697 & ~n31696;
  assign n31698 = ~n35470 | ~n43344;
  assign n31700 = ~n31699 | ~n31698;
  assign n31704 = ~n31701 & ~n31700;
  assign n31703 = ~n36906 | ~n31702;
  assign P1_U3031 = ~n31704 | ~n31703;
  assign n31707 = ~n35468 & ~n44019;
  assign n31706 = ~n31705 & ~n43300;
  assign n31709 = ~n31707 & ~n31706;
  assign n31708 = ~n44021 | ~n35470;
  assign P1_U2872 = ~n31709 | ~n31708;
  assign n31710 = ~n44000 | ~n31819;
  assign n31712 = ~n31710 | ~n36364;
  assign n35738 = ~n31712 | ~n31711;
  assign n31784 = ~n35738 | ~n35805;
  assign n31713 = ~P2_FLUSH_REG_SCAN_IN | ~n31784;
  assign P2_U2819 = ~n31714 | ~n31713;
  assign n31720 = ~n31960 | ~P1_EAX_REG_11__SCAN_IN;
  assign n31719 = ~P1_LWORD_REG_11__SCAN_IN | ~n32110;
  assign n31725 = n31720 & n31719;
  assign n31724 = ~DATAI_11_ | ~n39896;
  assign n31723 = ~n39901 | ~BUF1_REG_11__SCAN_IN;
  assign n42736 = ~n31724 | ~n31723;
  assign P1_U2963 = ~n31725 | ~n31748;
  assign n31727 = ~n31960 | ~P1_EAX_REG_30__SCAN_IN;
  assign n31726 = ~P1_UWORD_REG_14__SCAN_IN | ~n32110;
  assign n31730 = n31727 & n31726;
  assign n31729 = ~DATAI_14_ | ~n39896;
  assign n31728 = ~n39901 | ~BUF1_REG_14__SCAN_IN;
  assign n43305 = ~n31729 | ~n31728;
  assign n31981 = ~n32107 | ~n43305;
  assign P1_U2951 = ~n31730 | ~n31981;
  assign n31732 = ~P1_LWORD_REG_13__SCAN_IN | ~n32110;
  assign n31731 = ~n31960 | ~P1_EAX_REG_13__SCAN_IN;
  assign n31735 = n31732 & n31731;
  assign n31734 = ~DATAI_13_ | ~n39896;
  assign n31733 = ~n39901 | ~BUF1_REG_13__SCAN_IN;
  assign n43121 = ~n31734 | ~n31733;
  assign P1_U2965 = ~n31735 | ~n31757;
  assign n31737 = ~P1_UWORD_REG_8__SCAN_IN | ~n32110;
  assign n31736 = ~n31960 | ~P1_EAX_REG_24__SCAN_IN;
  assign n31740 = n31737 & n31736;
  assign n31739 = ~DATAI_8_ | ~n39896;
  assign n31738 = ~n39901 | ~BUF1_REG_8__SCAN_IN;
  assign n42043 = ~n31739 | ~n31738;
  assign n32055 = ~n32107 | ~n42043;
  assign P1_U2945 = ~n31740 | ~n32055;
  assign n31742 = ~P1_UWORD_REG_12__SCAN_IN | ~n32110;
  assign n31741 = ~n31960 | ~P1_EAX_REG_28__SCAN_IN;
  assign n31745 = n31742 & n31741;
  assign n31744 = ~DATAI_12_ | ~n39896;
  assign n31743 = ~n39901 | ~BUF1_REG_12__SCAN_IN;
  assign n42942 = ~n31744 | ~n31743;
  assign n32059 = ~n32107 | ~n42942;
  assign P1_U2949 = ~n31745 | ~n32059;
  assign n31747 = ~P1_UWORD_REG_11__SCAN_IN | ~n32110;
  assign n31746 = ~n31960 | ~P1_EAX_REG_27__SCAN_IN;
  assign n31749 = n31747 & n31746;
  assign P1_U2948 = ~n31749 | ~n31748;
  assign n31751 = ~P1_UWORD_REG_10__SCAN_IN | ~n32110;
  assign n31750 = ~n31960 | ~P1_EAX_REG_26__SCAN_IN;
  assign n31754 = n31751 & n31750;
  assign n31753 = ~DATAI_10_ | ~n39896;
  assign n31752 = ~n39901 | ~BUF1_REG_10__SCAN_IN;
  assign n42688 = ~n31753 | ~n31752;
  assign n32047 = ~n32107 | ~n42688;
  assign P1_U2947 = ~n31754 | ~n32047;
  assign n31756 = ~P1_UWORD_REG_13__SCAN_IN | ~n32110;
  assign n31755 = ~n31960 | ~P1_EAX_REG_29__SCAN_IN;
  assign n31758 = n31756 & n31755;
  assign P1_U2950 = ~n31758 | ~n31757;
  assign n31760 = ~P1_UWORD_REG_9__SCAN_IN | ~n32110;
  assign n31759 = ~n31960 | ~P1_EAX_REG_25__SCAN_IN;
  assign n31763 = n31760 & n31759;
  assign n31762 = ~DATAI_9_ | ~n39896;
  assign n31761 = ~n39901 | ~BUF1_REG_9__SCAN_IN;
  assign n42029 = ~n31762 | ~n31761;
  assign n32051 = ~n32107 | ~n42029;
  assign P1_U2946 = ~n31763 | ~n32051;
  assign n31786 = ~P2_MORE_REG_SCAN_IN | ~n31784;
  assign n31783 = ~n31765 & ~n31764;
  assign n31767 = ~n31766;
  assign n31769 = ~n31768 & ~n31767;
  assign n31776 = ~n31779 & ~n31769;
  assign n31774 = ~n31771 | ~n31770;
  assign n31773 = ~n35801 | ~n31772;
  assign n31775 = ~n31774 | ~n31773;
  assign n31781 = ~n31776 & ~n31775;
  assign n31778 = ~n31777;
  assign n31780 = ~n31779 | ~n31778;
  assign n31782 = ~n31781 | ~n31780;
  assign n35742 = ~n31783 & ~n31782;
  assign n31785 = n35742 | n31784;
  assign P2_U3609 = ~n31786 | ~n31785;
  assign n31789 = n40202 | n31788;
  assign n33488 = ~n42025 | ~n41362;
  assign n31792 = ~P3_FLUSH_REG_SCAN_IN | ~n31791;
  assign P3_U2637 = ~n33488 | ~n31792;
  assign n35485 = n31794 ^ n31793;
  assign n31798 = ~n35485 & ~n43298;
  assign n35484 = ~n31796 ^ n31795;
  assign n31797 = ~n35484 & ~n44019;
  assign n31800 = ~n31798 & ~n31797;
  assign n31799 = ~P1_EBX_REG_1__SCAN_IN | ~n44023;
  assign P1_U2871 = ~n31800 | ~n31799;
  assign n32526 = ~n32848 | ~n32196;
  assign n42052 = ~n32489 & ~n32526;
  assign n31811 = ~n32253;
  assign n35917 = ~P3_EBX_REG_0__SCAN_IN & ~P3_EBX_REG_1__SCAN_IN;
  assign n33507 = ~n31811 & ~n35917;
  assign n31813 = ~n42052 | ~n33507;
  assign n31812 = ~P3_EBX_REG_1__SCAN_IN | ~n32526;
  assign n31815 = n31813 & n31812;
  assign n31814 = ~P3_INSTQUEUE_REG_0__1__SCAN_IN | ~n42135;
  assign P3_U2702 = ~n31815 | ~n31814;
  assign n31822 = ~n31816 | ~P2_STATE2_REG_1__SCAN_IN;
  assign P2_U2920 = n33545 & P2_DATAO_REG_31__SCAN_IN;
  assign n32156 = n31826 & n32366;
  assign P3_U2736 = n43984 & P3_DATAO_REG_31__SCAN_IN;
  assign n31828 = ~P3_EAX_REG_8__SCAN_IN | ~n32156;
  assign n31827 = ~n32190 | ~P3_LWORD_REG_8__SCAN_IN;
  assign n31830 = n31828 & n31827;
  assign n31829 = ~n43984 | ~P3_DATAO_REG_8__SCAN_IN;
  assign P3_U2759 = ~n31830 | ~n31829;
  assign n31832 = ~P3_EAX_REG_10__SCAN_IN | ~n32156;
  assign n31831 = ~n32190 | ~P3_LWORD_REG_10__SCAN_IN;
  assign n31834 = n31832 & n31831;
  assign n31833 = ~n43984 | ~P3_DATAO_REG_10__SCAN_IN;
  assign P3_U2757 = ~n31834 | ~n31833;
  assign n31836 = ~P3_EAX_REG_9__SCAN_IN | ~n32156;
  assign n31835 = ~n32190 | ~P3_LWORD_REG_9__SCAN_IN;
  assign n31838 = n31836 & n31835;
  assign n31837 = ~n43984 | ~P3_DATAO_REG_9__SCAN_IN;
  assign P3_U2758 = ~n31838 | ~n31837;
  assign n31840 = ~P3_EAX_REG_5__SCAN_IN | ~n32156;
  assign n31839 = ~n32190 | ~P3_LWORD_REG_5__SCAN_IN;
  assign n31842 = n31840 & n31839;
  assign n31841 = ~n43984 | ~P3_DATAO_REG_5__SCAN_IN;
  assign P3_U2762 = ~n31842 | ~n31841;
  assign n31844 = ~P3_EAX_REG_2__SCAN_IN | ~n32156;
  assign n31843 = ~n32190 | ~P3_LWORD_REG_2__SCAN_IN;
  assign n31846 = n31844 & n31843;
  assign n31845 = ~n43984 | ~P3_DATAO_REG_2__SCAN_IN;
  assign P3_U2765 = ~n31846 | ~n31845;
  assign n31848 = ~n32190 | ~P3_LWORD_REG_7__SCAN_IN;
  assign n31847 = ~P3_EAX_REG_7__SCAN_IN | ~n32156;
  assign n31850 = n31848 & n31847;
  assign n31849 = ~n43984 | ~P3_DATAO_REG_7__SCAN_IN;
  assign P3_U2760 = ~n31850 | ~n31849;
  assign n31852 = ~P3_EAX_REG_3__SCAN_IN | ~n32156;
  assign n31851 = ~n32190 | ~P3_LWORD_REG_3__SCAN_IN;
  assign n31854 = n31852 & n31851;
  assign n31853 = ~n43984 | ~P3_DATAO_REG_3__SCAN_IN;
  assign P3_U2764 = ~n31854 | ~n31853;
  assign n31856 = ~P3_EAX_REG_1__SCAN_IN | ~n32156;
  assign n31855 = ~n32190 | ~P3_LWORD_REG_1__SCAN_IN;
  assign n31858 = n31856 & n31855;
  assign n31857 = ~n43984 | ~P3_DATAO_REG_1__SCAN_IN;
  assign P3_U2766 = ~n31858 | ~n31857;
  assign n31860 = ~P3_EAX_REG_4__SCAN_IN | ~n32156;
  assign n31859 = ~n32190 | ~P3_LWORD_REG_4__SCAN_IN;
  assign n31862 = n31860 & n31859;
  assign n31861 = ~n43984 | ~P3_DATAO_REG_4__SCAN_IN;
  assign P3_U2763 = ~n31862 | ~n31861;
  assign n31864 = ~n32190 | ~P3_LWORD_REG_0__SCAN_IN;
  assign n31863 = ~P3_EAX_REG_0__SCAN_IN | ~n32156;
  assign n31866 = n31864 & n31863;
  assign n31865 = ~n43984 | ~P3_DATAO_REG_0__SCAN_IN;
  assign P3_U2767 = ~n31866 | ~n31865;
  assign n31868 = ~P3_EAX_REG_6__SCAN_IN | ~n32156;
  assign n31867 = ~n32190 | ~P3_LWORD_REG_6__SCAN_IN;
  assign n31870 = n31868 & n31867;
  assign n31869 = ~n43984 | ~P3_DATAO_REG_6__SCAN_IN;
  assign P3_U2761 = ~n31870 | ~n31869;
  assign n31872 = ~P3_EAX_REG_14__SCAN_IN | ~n32156;
  assign n31871 = ~n32190 | ~P3_LWORD_REG_14__SCAN_IN;
  assign n31874 = n31872 & n31871;
  assign n31873 = ~n43984 | ~P3_DATAO_REG_14__SCAN_IN;
  assign P3_U2753 = ~n31874 | ~n31873;
  assign n31876 = ~P3_EAX_REG_15__SCAN_IN | ~n32156;
  assign n31875 = ~n32190 | ~P3_LWORD_REG_15__SCAN_IN;
  assign n31878 = n31876 & n31875;
  assign n31877 = ~n43984 | ~P3_DATAO_REG_15__SCAN_IN;
  assign P3_U2752 = ~n31878 | ~n31877;
  assign n31880 = ~P3_EAX_REG_13__SCAN_IN | ~n32156;
  assign n31879 = ~n32190 | ~P3_LWORD_REG_13__SCAN_IN;
  assign n31882 = n31880 & n31879;
  assign n31881 = ~n43984 | ~P3_DATAO_REG_13__SCAN_IN;
  assign P3_U2754 = ~n31882 | ~n31881;
  assign n31884 = ~P3_EAX_REG_12__SCAN_IN | ~n32156;
  assign n31883 = ~n32190 | ~P3_LWORD_REG_12__SCAN_IN;
  assign n31886 = n31884 & n31883;
  assign n31885 = ~n43984 | ~P3_DATAO_REG_12__SCAN_IN;
  assign P3_U2755 = ~n31886 | ~n31885;
  assign n31888 = ~P3_EAX_REG_11__SCAN_IN | ~n32156;
  assign n31887 = ~n32190 | ~P3_LWORD_REG_11__SCAN_IN;
  assign n31890 = n31888 & n31887;
  assign n31889 = ~n43984 | ~P3_DATAO_REG_11__SCAN_IN;
  assign P3_U2756 = ~n31890 | ~n31889;
  assign n39307 = ~P1_STATE2_REG_3__SCAN_IN;
  assign n34071 = ~P1_STATE2_REG_0__SCAN_IN & ~n39307;
  assign n31893 = ~n31892 & ~n31891;
  assign n31906 = n31894 | n31893;
  assign n31897 = ~n32131 | ~n31895;
  assign n31902 = ~n31897 | ~n31896;
  assign n31899 = ~n31898;
  assign n31900 = ~n31899 & ~n34515;
  assign n31901 = ~n31909 & ~n31900;
  assign n32234 = ~n31912 & ~n31911;
  assign n31915 = ~n34495 | ~n44102;
  assign n34523 = ~n34550 & ~n33710;
  assign n31914 = ~P1_FLUSH_REG_SCAN_IN | ~n34523;
  assign n32101 = ~n32341;
  assign n31917 = ~n32232;
  assign n31918 = ~n31917 | ~n31916;
  assign n31919 = ~n32337 & ~n31918;
  assign n31926 = ~n34552 | ~n32116;
  assign n31924 = ~n32080 | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n31940 = ~n31921;
  assign n31923 = ~n31940 | ~n31922;
  assign n31925 = ~n31924 | ~n31923;
  assign n34478 = ~n31926 | ~n31925;
  assign n31931 = ~n34478 | ~n32336;
  assign n31929 = ~n33714 & ~P1_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n35631 = ~n31927 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n31928 = ~n35631 & ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n31930 = ~n31929 & ~n31928;
  assign n31932 = ~n31931 | ~n31930;
  assign n31934 = ~n32101 | ~n31932;
  assign n31933 = ~n32341 | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign P1_U3474 = ~n31934 | ~n31933;
  assign n31935 = ~n35631;
  assign n32076 = ~n31935 | ~n32084;
  assign n31949 = ~n32076 & ~n33727;
  assign n31944 = ~n39301 | ~n32116;
  assign n31942 = ~n32080 & ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n31939 = ~n31938 & ~n31937;
  assign n31941 = ~n31940 & ~n31939;
  assign n31943 = ~n31942 & ~n31941;
  assign n34477 = ~n31944 | ~n31943;
  assign n31947 = ~n34477 | ~n32336;
  assign n32097 = ~P1_INSTADDRPOINTER_REG_31__SCAN_IN ^ n32556;
  assign n31945 = ~n32552 & ~n32097;
  assign n31946 = ~P1_STATE2_REG_1__SCAN_IN | ~n31945;
  assign n31948 = ~n31947 | ~n31946;
  assign n31950 = n31949 | n31948;
  assign n31952 = ~n32101 | ~n31950;
  assign n31951 = ~n32341 | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign P1_U3473 = ~n31952 | ~n31951;
  assign n35916 = ~P3_EBX_REG_2__SCAN_IN;
  assign n33163 = ~P3_EBX_REG_3__SCAN_IN;
  assign n33139 = ~n35916 & ~n33163;
  assign n32255 = ~P3_EBX_REG_4__SCAN_IN | ~n33139;
  assign n31955 = ~n32255 & ~n32253;
  assign n31957 = ~n42135 & ~n32671;
  assign n31956 = ~n33527 | ~n32251;
  assign n31959 = ~n31957 | ~n31956;
  assign n31958 = ~P3_INSTQUEUE_REG_0__7__SCAN_IN | ~n42135;
  assign P3_U2696 = ~n31959 | ~n31958;
  assign n31961 = ~P1_EAX_REG_18__SCAN_IN;
  assign n31964 = ~n31718 & ~n31961;
  assign n31963 = ~DATAI_2_ | ~n39896;
  assign n31962 = ~n39901 | ~BUF1_REG_2__SCAN_IN;
  assign n41049 = ~n31963 | ~n31962;
  assign n34228 = ~n41049;
  assign n32015 = ~n32237 & ~n34228;
  assign n31966 = ~n31964 & ~n32015;
  assign n31965 = ~P1_UWORD_REG_2__SCAN_IN | ~n32110;
  assign P1_U2939 = ~n31966 | ~n31965;
  assign n31967 = ~P1_EAX_REG_20__SCAN_IN;
  assign n31970 = ~n31718 & ~n31967;
  assign n31969 = ~DATAI_4_ | ~n39896;
  assign n31968 = ~n39901 | ~BUF1_REG_4__SCAN_IN;
  assign n41462 = ~n31969 | ~n31968;
  assign n34136 = ~n41462;
  assign n32023 = ~n32237 & ~n34136;
  assign n31972 = ~n31970 & ~n32023;
  assign n31971 = ~P1_UWORD_REG_4__SCAN_IN | ~n32110;
  assign P1_U2941 = ~n31972 | ~n31971;
  assign n31976 = ~n31718 & ~n31973;
  assign n31975 = ~DATAI_3_ | ~n39896;
  assign n31974 = ~n39901 | ~BUF1_REG_3__SCAN_IN;
  assign n41040 = ~n31975 | ~n31974;
  assign n34166 = ~n41040;
  assign n32011 = ~n32237 & ~n34166;
  assign n31978 = ~n31976 & ~n32011;
  assign n31977 = ~P1_UWORD_REG_3__SCAN_IN | ~n32110;
  assign P1_U2940 = ~n31978 | ~n31977;
  assign n31980 = ~n31718 & ~n44034;
  assign n31979 = P1_LWORD_REG_14__SCAN_IN & n32110;
  assign n31982 = ~n31980 & ~n31979;
  assign P1_U2966 = ~n31982 | ~n31981;
  assign n31986 = ~n31718 & ~n31983;
  assign n31985 = ~DATAI_1_ | ~n39896;
  assign n31984 = ~n39901 | ~BUF1_REG_1__SCAN_IN;
  assign n40550 = ~n31985 | ~n31984;
  assign n34189 = ~n40550;
  assign n32033 = ~n32237 & ~n34189;
  assign n31988 = ~n31986 & ~n32033;
  assign n31987 = ~P1_UWORD_REG_1__SCAN_IN | ~n32110;
  assign P1_U2938 = ~n31988 | ~n31987;
  assign n31992 = ~n31718 & ~n31989;
  assign n31991 = ~DATAI_0_ | ~n39896;
  assign n31990 = ~n39901 | ~BUF1_REG_0__SCAN_IN;
  assign n39894 = ~n31991 | ~n31990;
  assign n32007 = ~n32237 & ~n34243;
  assign n31994 = ~n31992 & ~n32007;
  assign n31993 = ~P1_UWORD_REG_0__SCAN_IN | ~n32110;
  assign P1_U2937 = ~n31994 | ~n31993;
  assign n31998 = ~n31718 & ~n31995;
  assign n31997 = ~DATAI_5_ | ~n39896;
  assign n31996 = ~n39901 | ~BUF1_REG_5__SCAN_IN;
  assign n41426 = ~n31997 | ~n31996;
  assign n34606 = ~n41426;
  assign n32019 = ~n32237 & ~n34606;
  assign n32000 = ~n31998 & ~n32019;
  assign n31999 = ~P1_UWORD_REG_5__SCAN_IN | ~n32110;
  assign P1_U2942 = ~n32000 | ~n31999;
  assign n32004 = ~n31718 & ~n32001;
  assign n32003 = ~DATAI_7_ | ~n39896;
  assign n32002 = ~n39901 | ~BUF1_REG_7__SCAN_IN;
  assign n41688 = ~n32003 | ~n32002;
  assign n34074 = ~n41688;
  assign n32037 = ~n32237 & ~n34074;
  assign n32006 = ~n32004 & ~n32037;
  assign n32005 = ~P1_UWORD_REG_7__SCAN_IN | ~n32110;
  assign P1_U2944 = ~n32006 | ~n32005;
  assign n32008 = ~n31718 & ~n24804;
  assign n32010 = ~n32008 & ~n32007;
  assign n32009 = ~P1_LWORD_REG_0__SCAN_IN | ~n32110;
  assign P1_U2952 = ~n32010 | ~n32009;
  assign n32012 = ~n31718 & ~n24818;
  assign n32014 = ~n32012 & ~n32011;
  assign n32013 = ~P1_LWORD_REG_3__SCAN_IN | ~n32110;
  assign P1_U2955 = ~n32014 | ~n32013;
  assign n32016 = ~n31718 & ~n24788;
  assign n32018 = ~n32016 & ~n32015;
  assign n32017 = ~P1_LWORD_REG_2__SCAN_IN | ~n32110;
  assign P1_U2954 = ~n32018 | ~n32017;
  assign n44068 = ~P1_EAX_REG_5__SCAN_IN;
  assign n32020 = ~n31718 & ~n44068;
  assign n32022 = ~n32020 & ~n32019;
  assign n32021 = ~P1_LWORD_REG_5__SCAN_IN | ~n32110;
  assign P1_U2957 = ~n32022 | ~n32021;
  assign n44073 = ~P1_EAX_REG_4__SCAN_IN;
  assign n32024 = ~n31718 & ~n44073;
  assign n32026 = ~n32024 & ~n32023;
  assign n32025 = ~P1_LWORD_REG_4__SCAN_IN | ~n32110;
  assign P1_U2956 = ~n32026 | ~n32025;
  assign n32027 = ~P1_EAX_REG_22__SCAN_IN;
  assign n32030 = ~n31718 & ~n32027;
  assign n32029 = ~DATAI_6_ | ~n39896;
  assign n32028 = ~n39901 | ~BUF1_REG_6__SCAN_IN;
  assign n41773 = ~n32029 | ~n32028;
  assign n34151 = ~n41773;
  assign n32041 = ~n32237 & ~n34151;
  assign n32032 = ~n32030 & ~n32041;
  assign n32031 = ~P1_UWORD_REG_6__SCAN_IN | ~n32110;
  assign P1_U2943 = ~n32032 | ~n32031;
  assign n44086 = ~P1_EAX_REG_1__SCAN_IN;
  assign n32034 = ~n31718 & ~n44086;
  assign n32036 = ~n32034 & ~n32033;
  assign n32035 = ~P1_LWORD_REG_1__SCAN_IN | ~n32110;
  assign P1_U2953 = ~n32036 | ~n32035;
  assign n32038 = ~n31718 & ~n24862;
  assign n32040 = ~n32038 & ~n32037;
  assign n32039 = ~P1_LWORD_REG_7__SCAN_IN | ~n32110;
  assign P1_U2959 = ~n32040 | ~n32039;
  assign n44063 = ~P1_EAX_REG_6__SCAN_IN;
  assign n32042 = ~n31718 & ~n44063;
  assign n32044 = ~n32042 & ~n32041;
  assign n32043 = ~P1_LWORD_REG_6__SCAN_IN | ~n32110;
  assign P1_U2958 = ~n32044 | ~n32043;
  assign n44044 = ~P1_EAX_REG_10__SCAN_IN;
  assign n32046 = ~n31718 & ~n44044;
  assign n32045 = P1_LWORD_REG_10__SCAN_IN & n32110;
  assign n32048 = ~n32046 & ~n32045;
  assign P1_U2962 = ~n32048 | ~n32047;
  assign n44049 = ~P1_EAX_REG_9__SCAN_IN;
  assign n32050 = ~n31718 & ~n44049;
  assign n32049 = P1_LWORD_REG_9__SCAN_IN & n32110;
  assign n32052 = ~n32050 & ~n32049;
  assign P1_U2961 = ~n32052 | ~n32051;
  assign n44054 = ~P1_EAX_REG_8__SCAN_IN;
  assign n32054 = ~n31718 & ~n44054;
  assign n32053 = P1_LWORD_REG_8__SCAN_IN & n32110;
  assign n32056 = ~n32054 & ~n32053;
  assign P1_U2960 = ~n32056 | ~n32055;
  assign n44039 = ~P1_EAX_REG_12__SCAN_IN;
  assign n32058 = ~n31718 & ~n44039;
  assign n32057 = P1_LWORD_REG_12__SCAN_IN & n32110;
  assign n32060 = ~n32058 & ~n32057;
  assign P1_U2964 = ~n32060 | ~n32059;
  assign n32064 = ~n32061;
  assign n32063 = ~n32062 | ~n32556;
  assign n32529 = ~n32064 | ~n32063;
  assign n32068 = ~n43358 & ~n32529;
  assign n32534 = ~n43033 & ~n35494;
  assign n32066 = ~n32534;
  assign n32065 = ~n43709 | ~P1_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n32067 = ~n32066 | ~n32065;
  assign n32072 = ~n32068 & ~n32067;
  assign n32070 = ~n43713 & ~P1_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n32069 = ~n35484 & ~n43729;
  assign n32071 = ~n32070 & ~n32069;
  assign P1_U2998 = ~n32072 | ~n32071;
  assign n32073 = ~P2_FLUSH_REG_SCAN_IN & ~n35801;
  assign n32074 = ~n35800 & ~n32073;
  assign P2_U3047 = ~n34913 & ~n32075;
  assign n32077 = ~n32101 | ~n32076;
  assign n32104 = ~n32077 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n32078 = ~n32118 | ~n32083;
  assign n32096 = ~n35631 & ~n32078;
  assign n34580 = ~n36136;
  assign n32090 = ~n34580 | ~n32116;
  assign n32079 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n32088 = ~n32080 & ~n32079;
  assign n32114 = ~n32082 | ~n32081;
  assign n32113 = ~n32084 | ~n32083;
  assign n32086 = ~n32113;
  assign n32085 = ~n32084 & ~n32083;
  assign n32091 = ~n32086 & ~n32085;
  assign n32087 = ~n32114 & ~n32091;
  assign n32089 = ~n32088 & ~n32087;
  assign n32094 = ~n32090 | ~n32089;
  assign n32092 = ~n32091;
  assign n32093 = ~n32123 & ~n32092;
  assign n33711 = ~n32094 & ~n32093;
  assign n32095 = ~n33711 & ~n32136;
  assign n32100 = ~n32096 & ~n32095;
  assign n32098 = P1_INSTADDRPOINTER_REG_0__SCAN_IN & n32097;
  assign n32099 = ~P1_STATE2_REG_1__SCAN_IN | ~n32098;
  assign n32102 = ~n32100 | ~n32099;
  assign n32103 = ~n32102 | ~n32101;
  assign P1_U3472 = ~n32104 | ~n32103;
  assign n32106 = ~DATAI_15_ | ~n39896;
  assign n32105 = ~n39901 | ~BUF1_REG_15__SCAN_IN;
  assign n39931 = ~n32106 | ~n32105;
  assign n32109 = n32107 & n39931;
  assign n44029 = ~P1_EAX_REG_15__SCAN_IN;
  assign n32108 = ~n31718 & ~n44029;
  assign n32112 = ~n32109 & ~n32108;
  assign n32111 = ~P1_LWORD_REG_15__SCAN_IN | ~n32110;
  assign P1_U2967 = ~n32112 | ~n32111;
  assign n32115 = n32113 ^ n33721;
  assign n32135 = ~n32115 & ~n32114;
  assign n35870 = ~n34569;
  assign n32117 = ~n32116;
  assign n32125 = ~n35870 & ~n32117;
  assign n32120 = ~n32118 & ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n32122 = ~n32120 & ~n32119;
  assign n32137 = ~n32122 | ~n32121;
  assign n32124 = ~n32123 & ~n32137;
  assign n32133 = ~n32125 & ~n32124;
  assign n32126 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n32129 = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n32126;
  assign n32128 = ~n32127;
  assign n32130 = ~n32129 | ~n32128;
  assign n32132 = ~n32131 | ~n32130;
  assign n32134 = ~n32133 | ~n32132;
  assign n32139 = ~n33718 & ~n32136;
  assign n32138 = ~n35631 & ~n32137;
  assign n32140 = ~n32139 & ~n32138;
  assign n32142 = n32341 | n32140;
  assign n32141 = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n32341;
  assign P1_U3469 = ~n32142 | ~n32141;
  assign n32146 = ~n37637 | ~n23415;
  assign n32151 = ~n32146 | ~n37302;
  assign n32150 = ~n32148 & ~n32147;
  assign n32153 = ~n32151 | ~n43525;
  assign n32152 = ~P2_EBX_REG_1__SCAN_IN | ~n35967;
  assign P2_U2886 = ~n32153 | ~n32152;
  assign n32155 = ~n43984 | ~P3_DATAO_REG_26__SCAN_IN;
  assign n32154 = ~n32190 | ~P3_UWORD_REG_10__SCAN_IN;
  assign n32158 = n32155 & n32154;
  assign n43982 = ~n32156 | ~n32860;
  assign n32157 = ~P3_EAX_REG_26__SCAN_IN | ~n32193;
  assign P3_U2741 = ~n32158 | ~n32157;
  assign n32160 = ~n43984 | ~P3_DATAO_REG_16__SCAN_IN;
  assign n32159 = ~n32190 | ~P3_UWORD_REG_0__SCAN_IN;
  assign n32162 = n32160 & n32159;
  assign n32161 = ~P3_EAX_REG_16__SCAN_IN | ~n32193;
  assign P3_U2751 = ~n32162 | ~n32161;
  assign n32164 = ~n43984 | ~P3_DATAO_REG_28__SCAN_IN;
  assign n32163 = ~n32190 | ~P3_UWORD_REG_12__SCAN_IN;
  assign n32166 = n32164 & n32163;
  assign n32165 = ~P3_EAX_REG_28__SCAN_IN | ~n32193;
  assign P3_U2739 = ~n32166 | ~n32165;
  assign n39510 = ~P2_STATEBS16_REG_SCAN_IN & ~n39524;
  assign n34901 = ~n36365 & ~n39510;
  assign n32170 = ~n37945 & ~n34901;
  assign n37303 = ~n32168 ^ n32167;
  assign n32169 = ~n32271 & ~n39522;
  assign n32171 = ~n32170 & ~n32169;
  assign n32900 = ~n37945 | ~n34909;
  assign n32172 = ~n32171 | ~n32900;
  assign n32174 = ~n34913 | ~n32172;
  assign n32173 = ~n34914 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign P2_U3604 = ~n32174 | ~n32173;
  assign n32179 = ~n32175 & ~n39522;
  assign n32178 = ~n32177 & ~n32176;
  assign n32182 = ~n32179 & ~n32178;
  assign n32181 = n38279 | n32180;
  assign n32183 = ~n32182 | ~n32181;
  assign n32185 = ~n34913 | ~n32183;
  assign n32184 = ~n34914 | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign P2_U3605 = ~n32185 | ~n32184;
  assign n32187 = ~n36280 & ~n43982;
  assign n32186 = n43984 & P3_DATAO_REG_30__SCAN_IN;
  assign n32189 = ~n32187 & ~n32186;
  assign n32188 = ~n32190 | ~P3_UWORD_REG_14__SCAN_IN;
  assign P3_U2737 = ~n32189 | ~n32188;
  assign n32192 = ~n32190 | ~P3_UWORD_REG_3__SCAN_IN;
  assign n32191 = ~n43984 | ~P3_DATAO_REG_19__SCAN_IN;
  assign n32195 = n32192 & n32191;
  assign n32194 = ~P3_EAX_REG_19__SCAN_IN | ~n32193;
  assign P3_U2748 = ~n32195 | ~n32194;
  assign n32824 = ~n32279 & ~n32280;
  assign n32816 = ~P3_EAX_REG_2__SCAN_IN | ~n32824;
  assign n32814 = ~n32815 & ~n32816;
  assign n33090 = ~n32202 & ~n32201;
  assign n32203 = ~n32814 | ~n32807;
  assign n32205 = ~n32204 | ~n32203;
  assign n34968 = ~n32672 & ~n33090;
  assign n32498 = ~n32204 & ~n32203;
  assign n32497 = ~n34968 & ~n32498;
  assign n32212 = ~n32205 | ~n32497;
  assign n32210 = ~n34843 & ~n32207;
  assign n35459 = ~n32807 | ~n35267;
  assign n32209 = ~n35459 & ~n32208;
  assign n32211 = ~n32210 & ~n32209;
  assign P3_U2731 = ~n32212 | ~n32211;
  assign n37280 = n32214 ^ n32213;
  assign n32216 = ~n37947 & ~n37280;
  assign n32273 = ~n37947 | ~n37280;
  assign n32215 = ~n43693 | ~n32273;
  assign n32222 = ~n32216 & ~n32215;
  assign n32220 = ~n41756 | ~n37280;
  assign n32218 = ~n32217;
  assign n32219 = ~n36955 | ~n37112;
  assign n32221 = ~n32220 | ~n32219;
  assign n32224 = ~n32222 & ~n32221;
  assign n32223 = ~P2_EAX_REG_0__SCAN_IN | ~n43698;
  assign P2_U2919 = ~n32224 | ~n32223;
  assign n32227 = ~n36002 & ~n32225;
  assign n32226 = ~n25671 & ~n41759;
  assign n32229 = ~n32227 & ~n32226;
  assign n32228 = n39737 | n33786;
  assign P2_U2913 = ~n32229 | ~n32228;
  assign n32230 = ~n34134 | ~n39892;
  assign n32231 = ~n32230 & ~n34149;
  assign n32241 = ~n32239 | ~n32238;
  assign n32240 = ~n32241;
  assign n34898 = ~n43734 | ~n32240;
  assign n32244 = ~n34898 & ~n34243;
  assign n32242 = n43734 & n32241;
  assign n32243 = ~n39934 & ~n35468;
  assign n32246 = ~n32244 & ~n32243;
  assign n32245 = ~P1_EAX_REG_0__SCAN_IN | ~n43732;
  assign P1_U2904 = ~n32246 | ~n32245;
  assign n32248 = ~n34898 & ~n34189;
  assign n32247 = ~n39934 & ~n35484;
  assign n32250 = ~n32248 & ~n32247;
  assign n32249 = ~P1_EAX_REG_1__SCAN_IN | ~n43732;
  assign P1_U2903 = ~n32250 | ~n32249;
  assign n32252 = ~P3_EBX_REG_6__SCAN_IN | ~n32251;
  assign n32257 = ~n32252 & ~n42135;
  assign n43932 = ~n32253 & ~n41059;
  assign n32254 = ~n43932;
  assign n33480 = ~n32255 & ~n32254;
  assign n33481 = ~P3_EBX_REG_5__SCAN_IN | ~n33480;
  assign n32256 = ~n33481 & ~P3_EBX_REG_6__SCAN_IN;
  assign n32259 = ~n32257 & ~n32256;
  assign n32258 = ~P3_INSTQUEUE_REG_0__6__SCAN_IN | ~n42135;
  assign P3_U2697 = ~n32259 | ~n32258;
  assign n32262 = ~n36002 & ~n41757;
  assign n32261 = ~n32260 & ~n41759;
  assign n32266 = ~n32262 & ~n32261;
  assign n41081 = ~n32264 ^ n32263;
  assign n32265 = ~n41081 | ~n35381;
  assign P2_U2911 = ~n32266 | ~n32265;
  assign n32270 = ~n43695 & ~n32271;
  assign n32268 = ~P2_EAX_REG_1__SCAN_IN | ~n43698;
  assign n32267 = ~n36955 | ~n37434;
  assign n32269 = ~n32268 | ~n32267;
  assign n32278 = ~n32270 & ~n32269;
  assign n32272 = ~n37637 & ~n37303;
  assign n33217 = ~n37945 & ~n32271;
  assign n32274 = n32272 | n33217;
  assign n33216 = ~n32274 & ~n32273;
  assign n32276 = ~n33216 & ~n41754;
  assign n32275 = ~n32274 | ~n32273;
  assign n32277 = ~n32276 | ~n32275;
  assign P2_U2918 = ~n32278 | ~n32277;
  assign n32813 = ~n36242;
  assign n33094 = ~P3_EAX_REG_0__SCAN_IN & ~n32813;
  assign n32822 = ~n33090 & ~n33094;
  assign n32282 = ~n32279 & ~n32822;
  assign n32821 = ~n36242 | ~n32279;
  assign n32281 = ~n32280 & ~n32821;
  assign n32288 = ~n32282 & ~n32281;
  assign n32286 = ~n34843 & ~n32283;
  assign n32285 = ~n35459 & ~n32284;
  assign n32287 = ~n32286 & ~n32285;
  assign P3_U2734 = ~n32288 | ~n32287;
  assign n32289 = ~n37947 | ~n23415;
  assign n32290 = ~n32289 | ~n37279;
  assign n32292 = ~n32290 | ~n43525;
  assign n32291 = ~P2_EBX_REG_0__SCAN_IN | ~n35967;
  assign P2_U2887 = ~n32292 | ~n32291;
  assign n32294 = ~n22917 | ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n32293 = ~n36311 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n32298 = ~n32294 | ~n32293;
  assign n32296 = ~n22913 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n32295 = ~n36307 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n32297 = ~n32296 | ~n32295;
  assign n32306 = ~n32298 & ~n32297;
  assign n32300 = ~n22903 | ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n32299 = ~n36317 | ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n32304 = ~n32300 | ~n32299;
  assign n32302 = ~n22910 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n32301 = ~n22914 | ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n32303 = ~n32302 | ~n32301;
  assign n32305 = ~n32304 & ~n32303;
  assign n32322 = ~n32306 | ~n32305;
  assign n32308 = ~n22902 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n32307 = ~n22912 | ~P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n32312 = ~n32308 | ~n32307;
  assign n32310 = ~n36298 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n32309 = ~n22923 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n32311 = ~n32310 | ~n32309;
  assign n32320 = ~n32312 & ~n32311;
  assign n32314 = ~n22919 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n32313 = ~n35392 | ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n32318 = ~n32314 | ~n32313;
  assign n32316 = ~n36294 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n32315 = ~n36320 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n32317 = ~n32316 | ~n32315;
  assign n32319 = ~n32318 & ~n32317;
  assign n32321 = ~n32320 | ~n32319;
  assign n32677 = ~n32322 & ~n32321;
  assign n32325 = ~n35459 & ~n32677;
  assign n32324 = ~n32323 & ~n34843;
  assign n32333 = ~n32325 & ~n32324;
  assign n32329 = ~P3_EAX_REG_8__SCAN_IN | ~n36243;
  assign n32327 = ~P3_EAX_REG_4__SCAN_IN | ~n32814;
  assign n32326 = ~P3_EAX_REG_6__SCAN_IN | ~P3_EAX_REG_5__SCAN_IN;
  assign n32485 = ~n32327 & ~n32326;
  assign n32357 = ~n32330;
  assign n32331 = ~n32329 | ~n32357;
  assign n32332 = ~n32331 | ~n32838;
  assign P3_U2727 = ~n32333 | ~n32332;
  assign n32335 = ~n32334 & ~n34258;
  assign n35500 = n32335 ^ n24830;
  assign n32338 = ~n32337 | ~n32336;
  assign n32339 = ~n35500 & ~n32338;
  assign n32343 = ~n32340 | ~n32339;
  assign n32342 = ~n32341 | ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign P1_U3468 = ~n32343 | ~n32342;
  assign n32346 = ~n32345 & ~n32344;
  assign n40775 = ~n32347 & ~n32346;
  assign n32350 = n40775 & n35381;
  assign n32349 = ~n36002 & ~n32348;
  assign n32352 = ~n32350 & ~n32349;
  assign n32351 = ~P2_EAX_REG_7__SCAN_IN | ~n43698;
  assign P2_U2912 = ~n32352 | ~n32351;
  assign n32355 = n36333 & n39615;
  assign n32354 = ~n34843 & ~n32353;
  assign n32360 = ~n32355 & ~n32354;
  assign n32356 = ~P3_EAX_REG_7__SCAN_IN | ~n36243;
  assign n32358 = ~n32356 | ~n32566;
  assign n32359 = ~n32358 | ~n32357;
  assign P3_U2728 = ~n32360 | ~n32359;
  assign n35670 = ~n36057;
  assign n32365 = ~n33486 & ~n32361;
  assign n32363 = ~n36052 | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n32364 = ~n32363 | ~n32362;
  assign n41363 = ~n32365 | ~n32364;
  assign n32378 = ~n35670 & ~n41363;
  assign n32375 = ~n41371 & ~n41374;
  assign n32377 = ~n32375 & ~n32374;
  assign n32376 = ~P3_FLUSH_REG_SCAN_IN | ~n41672;
  assign n32380 = ~n32378 | ~n36061;
  assign n32379 = ~n36063 | ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign P3_U3284 = ~n32380 | ~n32379;
  assign n32382 = ~n36294 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n32381 = ~n36311 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n32386 = ~n32382 | ~n32381;
  assign n32384 = ~n35392 | ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n32383 = ~n36320 | ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n32385 = ~n32384 | ~n32383;
  assign n32394 = ~n32386 & ~n32385;
  assign n32388 = ~n22903 | ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n32387 = ~n36317 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n32392 = ~n32388 | ~n32387;
  assign n32390 = ~n22919 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n32389 = ~n36307 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n32391 = ~n32390 | ~n32389;
  assign n32393 = ~n32392 & ~n32391;
  assign n32410 = ~n32394 | ~n32393;
  assign n32396 = ~n22902 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n32395 = ~n22920 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n32400 = ~n32396 | ~n32395;
  assign n32398 = ~n36310 | ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n32397 = ~n22913 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n32399 = ~n32398 | ~n32397;
  assign n32408 = ~n32400 & ~n32399;
  assign n32402 = ~n36298 | ~P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n32401 = ~n22923 | ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n32406 = ~n32402 | ~n32401;
  assign n32404 = ~n22914 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n32403 = ~n22917 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n32405 = ~n32404 | ~n32403;
  assign n32407 = ~n32406 & ~n32405;
  assign n32409 = ~n32408 | ~n32407;
  assign n32613 = ~n32410 & ~n32409;
  assign n32412 = ~n36298 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n32411 = ~n36307 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n32416 = ~n32412 | ~n32411;
  assign n32414 = ~n35392 | ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n32413 = ~n22923 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n32415 = ~n32414 | ~n32413;
  assign n32424 = ~n32416 & ~n32415;
  assign n32418 = ~n22903 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n32417 = ~n36317 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n32422 = ~n32418 | ~n32417;
  assign n32420 = ~n36310 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n32419 = ~n22914 | ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n32421 = ~n32420 | ~n32419;
  assign n32423 = ~n32422 & ~n32421;
  assign n32440 = ~n32424 | ~n32423;
  assign n32426 = ~n36320 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n32425 = ~n36311 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n32430 = ~n32426 | ~n32425;
  assign n32428 = ~n36294 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n32427 = ~n22913 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n32429 = ~n32428 | ~n32427;
  assign n32438 = ~n32430 & ~n32429;
  assign n32432 = ~n22919 | ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n32431 = ~n22902 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n32436 = ~n32432 | ~n32431;
  assign n32434 = ~n22917 | ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n32433 = ~n22920 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n32435 = ~n32434 | ~n32433;
  assign n32437 = ~n32436 & ~n32435;
  assign n32439 = ~n32438 | ~n32437;
  assign n32612 = ~n32440 & ~n32439;
  assign n32787 = ~n32613 & ~n32612;
  assign n32442 = ~n22902 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n32441 = ~n36311 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n32445 = ~n32442 | ~n32441;
  assign n34768 = ~n22923;
  assign n32443 = ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n32444 = ~n34768 & ~n32443;
  assign n32447 = ~n32445 & ~n32444;
  assign n32446 = ~n36294 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n32451 = ~n32447 | ~n32446;
  assign n32449 = ~n36310 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n32448 = ~n22914 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n32450 = ~n32449 | ~n32448;
  assign n32471 = ~n32451 & ~n32450;
  assign n32453 = ~n36317 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n32452 = ~n36307 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n32457 = ~n32453 | ~n32452;
  assign n32455 = ~n22913 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n32454 = ~n22920 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n32456 = ~n32455 | ~n32454;
  assign n32465 = ~n32457 & ~n32456;
  assign n32459 = ~n22903 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n32458 = ~n35392 | ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n32463 = ~n32459 | ~n32458;
  assign n32461 = ~n22917 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n32460 = ~n36320 | ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n32462 = ~n32461 | ~n32460;
  assign n32464 = ~n32463 & ~n32462;
  assign n32469 = ~n32465 | ~n32464;
  assign n32467 = ~n22919 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n32466 = ~n36298 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n32468 = ~n32467 | ~n32466;
  assign n32470 = ~n32469 & ~n32468;
  assign n32786 = ~n32471 | ~n32470;
  assign n40542 = n32787 ^ n32786;
  assign n32474 = ~n36333 | ~n40542;
  assign n32473 = ~n36282 | ~BUF2_REG_24__SCAN_IN;
  assign n32493 = ~n32474 | ~n32473;
  assign n32491 = ~BUF2_REG_8__SCAN_IN | ~n36338;
  assign n32476 = ~P3_EAX_REG_19__SCAN_IN | ~P3_EAX_REG_17__SCAN_IN;
  assign n32986 = ~n43977 & ~n32476;
  assign n32477 = ~P3_EAX_REG_21__SCAN_IN | ~P3_EAX_REG_20__SCAN_IN;
  assign n32478 = ~n43962 & ~n32477;
  assign n32487 = ~n32986 | ~n32478;
  assign n35694 = ~P3_EAX_REG_15__SCAN_IN | ~P3_EAX_REG_14__SCAN_IN;
  assign n32480 = ~P3_EAX_REG_11__SCAN_IN | ~P3_EAX_REG_10__SCAN_IN;
  assign n32479 = ~P3_EAX_REG_13__SCAN_IN | ~P3_EAX_REG_12__SCAN_IN;
  assign n34967 = ~n32480 & ~n32479;
  assign n32482 = ~P3_EAX_REG_9__SCAN_IN | ~P3_EAX_REG_8__SCAN_IN;
  assign n32481 = ~P3_EAX_REG_7__SCAN_IN | ~P3_EAX_REG_16__SCAN_IN;
  assign n32483 = ~n32482 & ~n32481;
  assign n32484 = ~n34967 | ~n32483;
  assign n32565 = ~n35694 & ~n32484;
  assign n32486 = ~n32485 | ~n32565;
  assign n32607 = ~n32487 & ~n32486;
  assign n32488 = ~n32607 & ~n32489;
  assign n32490 = ~n32792 | ~n43952;
  assign n32492 = ~n32491 | ~n32490;
  assign n32496 = ~n32493 & ~n32492;
  assign n32495 = ~P3_EAX_REG_24__SCAN_IN | ~n32494;
  assign P3_U2711 = ~n32496 | ~n32495;
  assign n32513 = ~n32497 & ~n32499;
  assign n32516 = ~n32672 | ~n32498;
  assign n32500 = n32499 & n32516;
  assign n32503 = ~n32513 & ~n32500;
  assign n32502 = n36333 & n32501;
  assign n32505 = ~n32503 & ~n32502;
  assign n32504 = ~BUF2_REG_5__SCAN_IN | ~n35462;
  assign P3_U2730 = ~n32505 | ~n32504;
  assign n32510 = ~n36543 & ~n36532;
  assign n32507 = ~n32506 & ~n35715;
  assign n32508 = ~n32507 & ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n35740 = ~n32509 & ~n32508;
  assign n32512 = ~n32510 | ~n35740;
  assign n32511 = ~n36543 | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign P2_U3595 = ~n32512 | ~n32511;
  assign n32514 = ~n34968 & ~n32513;
  assign n32523 = ~n32514 | ~P3_EAX_REG_6__SCAN_IN;
  assign n32521 = ~n35459 & ~n32515;
  assign n32517 = ~P3_EAX_REG_6__SCAN_IN & ~n32516;
  assign n32519 = ~n32517 | ~P3_EAX_REG_5__SCAN_IN;
  assign n32518 = ~n35462 | ~BUF2_REG_6__SCAN_IN;
  assign n32520 = ~n32519 | ~n32518;
  assign n32522 = ~n32521 & ~n32520;
  assign P3_U2729 = ~n32523 | ~n32522;
  assign n32525 = ~n41059 & ~P3_EBX_REG_0__SCAN_IN;
  assign n35407 = ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n43930 = ~n42135;
  assign n32524 = ~n35407 & ~n43930;
  assign n32528 = ~n32525 & ~n32524;
  assign n32527 = ~P3_EBX_REG_0__SCAN_IN | ~n32526;
  assign P3_U2703 = ~n32528 | ~n32527;
  assign n32538 = ~n43341 & ~n32529;
  assign n32531 = ~n42922 & ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n32530 = ~n35485 & ~n43441;
  assign n32536 = ~n32531 & ~n32530;
  assign n32533 = ~n32556 & ~n32532;
  assign n32535 = ~n32534 & ~n32533;
  assign n32537 = ~n32536 | ~n32535;
  assign n32543 = ~n32538 & ~n32537;
  assign n32539 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN & ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n32541 = ~n32539 & ~n42927;
  assign n32542 = ~n32541 | ~n32540;
  assign P1_U3030 = ~n32543 | ~n32542;
  assign n32544 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN & ~n34279;
  assign n32564 = ~n32544 | ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n32548 = n32546 | n32545;
  assign n32624 = ~n32548 | ~n32547;
  assign n32562 = ~n43341 & ~n32624;
  assign n32626 = ~P1_REIP_REG_2__SCAN_IN | ~n43469;
  assign n44022 = n32550 ^ n32549;
  assign n32551 = ~n44022 | ~n43344;
  assign n32555 = ~n32626 | ~n32551;
  assign n34286 = ~n32552 & ~n34283;
  assign n32553 = ~n34286 & ~n34290;
  assign n32554 = ~n41976 & ~n32553;
  assign n32560 = ~n32555 & ~n32554;
  assign n32557 = ~n32556 | ~n41979;
  assign n32558 = ~n32557 | ~n36893;
  assign n32559 = ~n32558 | ~P1_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n32561 = ~n32560 | ~n32559;
  assign n32563 = ~n32562 & ~n32561;
  assign P1_U3029 = ~n32564 | ~n32563;
  assign n32567 = ~n32565;
  assign n32985 = ~n32567 & ~n32566;
  assign n33268 = P3_EAX_REG_17__SCAN_IN & n32985;
  assign n32568 = ~n43983 & ~n34968;
  assign n32569 = ~n32985 & ~n32568;
  assign n32573 = ~n33268 & ~n32569;
  assign n32571 = ~n36282 | ~BUF2_REG_17__SCAN_IN;
  assign n32570 = ~n36338 | ~BUF2_REG_1__SCAN_IN;
  assign n32572 = ~n32571 | ~n32570;
  assign n32605 = ~n32573 & ~n32572;
  assign n32575 = ~n36320 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n32574 = ~n36311 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n32579 = ~n32575 | ~n32574;
  assign n32577 = ~n22913 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n32576 = ~n35392 | ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n32578 = ~n32577 | ~n32576;
  assign n32603 = ~n32579 & ~n32578;
  assign n32581 = ~n36294 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n32580 = ~n22910 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n32585 = ~n32581 | ~n32580;
  assign n32583 = ~n36298 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n32582 = ~n22917 | ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n32584 = ~n32583 | ~n32582;
  assign n32593 = ~n32585 & ~n32584;
  assign n32587 = ~n22903 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n32586 = ~n36317 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n32591 = ~n32587 | ~n32586;
  assign n32589 = ~n22902 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n32588 = ~n36307 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n32590 = ~n32589 | ~n32588;
  assign n32592 = ~n32591 & ~n32590;
  assign n32601 = ~n32593 | ~n32592;
  assign n32595 = ~n22919 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n32594 = ~n22914 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n32599 = ~n32595 | ~n32594;
  assign n32597 = ~n22923 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n32596 = ~n22912 | ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n32598 = ~n32597 | ~n32596;
  assign n32600 = n32599 | n32598;
  assign n32602 = ~n32601 & ~n32600;
  assign n35550 = ~n32603 | ~n32602;
  assign n32604 = ~n36333 | ~n35550;
  assign P3_U2718 = ~n32605 | ~n32604;
  assign n32617 = ~n32606 & ~n43957;
  assign n32609 = ~n32607;
  assign n32611 = ~n32609 & ~n32608;
  assign n32610 = BUF2_REG_23__SCAN_IN & n36282;
  assign n32615 = ~n32611 & ~n32610;
  assign n39740 = n32613 ^ n32612;
  assign n32614 = ~n39740 | ~n36333;
  assign n32616 = ~n32615 | ~n32614;
  assign n32619 = ~n32617 & ~n32616;
  assign n32618 = ~BUF2_REG_7__SCAN_IN | ~n36338;
  assign P3_U2712 = ~n32619 | ~n32618;
  assign n32621 = ~P2_EAX_REG_10__SCAN_IN | ~n43698;
  assign n32620 = ~n36955 | ~n41831;
  assign n32623 = n32621 & n32620;
  assign n32622 = n40298 | n33786;
  assign P2_U2909 = ~n32623 | ~n32622;
  assign n32628 = ~n43358 & ~n32624;
  assign n32625 = ~n43709 | ~P1_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n32627 = ~n32626 | ~n32625;
  assign n32636 = ~n32628 & ~n32627;
  assign n32634 = ~n36144 & ~n43713;
  assign n32632 = n32630 | n32629;
  assign n32633 = ~n44020 & ~n43729;
  assign n32635 = ~n32634 & ~n32633;
  assign P1_U2997 = ~n32636 | ~n32635;
  assign n32638 = ~n34898 & ~n34228;
  assign n32637 = ~n39934 & ~n44020;
  assign n32640 = ~n32638 & ~n32637;
  assign n32639 = ~P1_EAX_REG_2__SCAN_IN | ~n43732;
  assign P1_U2902 = ~n32640 | ~n32639;
  assign n32642 = ~n22919 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n32641 = ~n36317 | ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n32646 = ~n32642 | ~n32641;
  assign n32644 = ~n22914 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n32643 = ~n22917 | ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n32645 = ~n32644 | ~n32643;
  assign n32654 = ~n32646 & ~n32645;
  assign n32648 = ~n22903 | ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n32647 = ~n36310 | ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n32652 = ~n32648 | ~n32647;
  assign n32650 = ~n36298 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n32649 = ~n35392 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n32651 = ~n32650 | ~n32649;
  assign n32653 = ~n32652 & ~n32651;
  assign n32670 = ~n32654 | ~n32653;
  assign n32656 = ~n22902 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n32655 = ~n22920 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n32660 = ~n32656 | ~n32655;
  assign n32658 = ~n36294 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n32657 = ~n36320 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n32659 = ~n32658 | ~n32657;
  assign n32668 = ~n32660 & ~n32659;
  assign n32662 = ~n22913 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n32661 = ~n36311 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n32666 = ~n32662 | ~n32661;
  assign n32664 = ~n36307 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n32663 = ~n22923 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n32665 = ~n32664 | ~n32663;
  assign n32667 = ~n32666 & ~n32665;
  assign n32669 = ~n32668 | ~n32667;
  assign n33221 = ~n32670 & ~n32669;
  assign n32676 = n33221 | n43930;
  assign n32673 = ~P3_EBX_REG_10__SCAN_IN | ~n43930;
  assign n32674 = ~n32673 | ~n32716;
  assign n33066 = ~P3_EBX_REG_10__SCAN_IN;
  assign n32750 = ~n32752;
  assign n32675 = ~n32674 | ~n32750;
  assign P3_U2693 = ~n32676 | ~n32675;
  assign n32683 = n32677 | n43930;
  assign n32679 = ~P3_EBX_REG_8__SCAN_IN | ~n43930;
  assign n32681 = ~n32679 | ~n32678;
  assign n32714 = ~n32680;
  assign n32682 = ~n32681 | ~n32714;
  assign P3_U2695 = ~n32683 | ~n32682;
  assign n32685 = ~n22903 | ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n32684 = ~n22913 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n32689 = ~n32685 | ~n32684;
  assign n32687 = ~n22917 | ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n32686 = ~n36320 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n32688 = ~n32687 | ~n32686;
  assign n32697 = ~n32689 & ~n32688;
  assign n32691 = ~n22919 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n32690 = ~n36317 | ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n32695 = ~n32691 | ~n32690;
  assign n32693 = ~n22909 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n32692 = ~n35392 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n32694 = ~n32693 | ~n32692;
  assign n32696 = ~n32695 & ~n32694;
  assign n32713 = ~n32697 | ~n32696;
  assign n32699 = ~n22910 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n32698 = ~n22912 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n32703 = ~n32699 | ~n32698;
  assign n32701 = ~n36294 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n32700 = ~n36307 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n32702 = ~n32701 | ~n32700;
  assign n32711 = ~n32703 & ~n32702;
  assign n32705 = ~n22902 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n32704 = ~n22914 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n32709 = ~n32705 | ~n32704;
  assign n32707 = ~n22923 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n32706 = ~n36311 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n32708 = ~n32707 | ~n32706;
  assign n32710 = ~n32709 & ~n32708;
  assign n32712 = ~n32711 | ~n32710;
  assign n32833 = ~n32713 & ~n32712;
  assign n32719 = n32833 | n43930;
  assign n32715 = ~P3_EBX_REG_9__SCAN_IN | ~n43930;
  assign n32717 = ~n32715 | ~n32714;
  assign n32718 = ~n32717 | ~n32716;
  assign P3_U2694 = ~n32719 | ~n32718;
  assign n32721 = ~n22919 | ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n32720 = ~n22903 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n32725 = ~n32721 | ~n32720;
  assign n32723 = ~n22914 | ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n32722 = ~n22917 | ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n32724 = ~n32723 | ~n32722;
  assign n32733 = ~n32725 & ~n32724;
  assign n32727 = ~n36317 | ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n32726 = ~n22923 | ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n32731 = ~n32727 | ~n32726;
  assign n32729 = ~n36298 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n32728 = ~n35392 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n32730 = ~n32729 | ~n32728;
  assign n32732 = ~n32731 & ~n32730;
  assign n32749 = ~n32733 | ~n32732;
  assign n32735 = ~n36320 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n32734 = ~n22920 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n32739 = ~n32735 | ~n32734;
  assign n32737 = ~n36310 | ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n32736 = ~n36311 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n32738 = ~n32737 | ~n32736;
  assign n32747 = ~n32739 & ~n32738;
  assign n32741 = ~n36294 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n32740 = ~n22902 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n32745 = ~n32741 | ~n32740;
  assign n32743 = ~n22913 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n32742 = ~n36307 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n32744 = ~n32743 | ~n32742;
  assign n32746 = ~n32745 & ~n32744;
  assign n32748 = ~n32747 | ~n32746;
  assign n34350 = ~n32749 & ~n32748;
  assign n32755 = n34350 | n43930;
  assign n32751 = ~P3_EBX_REG_11__SCAN_IN | ~n43930;
  assign n32753 = ~n32751 | ~n32750;
  assign n32754 = ~n32753 | ~n32938;
  assign P3_U2692 = ~n32755 | ~n32754;
  assign n32791 = BUF2_REG_25__SCAN_IN & n36282;
  assign n32757 = ~n22902 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n32756 = ~n36311 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n32761 = ~n32757 | ~n32756;
  assign n32759 = ~n35392 | ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n32758 = ~n36320 | ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n32760 = ~n32759 | ~n32758;
  assign n32769 = ~n32761 & ~n32760;
  assign n32763 = ~n22903 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n32762 = ~n36317 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n32767 = ~n32763 | ~n32762;
  assign n32765 = ~n36298 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n32764 = ~n22913 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n32766 = ~n32765 | ~n32764;
  assign n32768 = ~n32767 & ~n32766;
  assign n32785 = ~n32769 | ~n32768;
  assign n32771 = ~n22917 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n32770 = ~n36307 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n32775 = ~n32771 | ~n32770;
  assign n32773 = ~n22919 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n32772 = ~n36310 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n32774 = ~n32773 | ~n32772;
  assign n32783 = ~n32775 & ~n32774;
  assign n32777 = ~n22914 | ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n32776 = ~n22920 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n32781 = ~n32777 | ~n32776;
  assign n32779 = ~n36294 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n32778 = ~n22923 | ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n32780 = ~n32779 | ~n32778;
  assign n32782 = ~n32781 & ~n32780;
  assign n32784 = ~n32783 | ~n32782;
  assign n33169 = ~n32785 & ~n32784;
  assign n33168 = ~n32787 | ~n32786;
  assign n40809 = n33169 ^ n33168;
  assign n32789 = ~n36333 | ~n40809;
  assign n32788 = ~n36338 | ~BUF2_REG_9__SCAN_IN;
  assign n32790 = ~n32789 | ~n32788;
  assign n32797 = ~n32791 & ~n32790;
  assign n32793 = ~P3_EAX_REG_25__SCAN_IN | ~n36243;
  assign n32795 = ~n32793 | ~n32794;
  assign n33206 = ~n33208;
  assign n32796 = ~n32795 | ~n33206;
  assign P3_U2710 = ~n32797 | ~n32796;
  assign n32802 = ~n32798;
  assign n32801 = ~n32800 | ~n32799;
  assign n32804 = ~n41703 & ~n33786;
  assign n32803 = ~n25724 & ~n41759;
  assign n32806 = ~n32804 & ~n32803;
  assign n32805 = ~n36955 | ~n41659;
  assign P2_U2910 = ~n32806 | ~n32805;
  assign n32812 = ~n32807 & ~n32815;
  assign n32810 = ~n35462 | ~BUF2_REG_3__SCAN_IN;
  assign n32809 = ~n32808 | ~n36333;
  assign n32811 = ~n32810 | ~n32809;
  assign n32820 = ~n32812 & ~n32811;
  assign n32818 = ~n32814 & ~n32813;
  assign n32817 = ~n32816 | ~n32815;
  assign n32819 = ~n32818 | ~n32817;
  assign P3_U2732 = ~n32820 | ~n32819;
  assign n32823 = ~n32822 | ~n32821;
  assign n32832 = ~n32823 | ~P3_EAX_REG_2__SCAN_IN;
  assign n32825 = ~n32824 | ~n36242;
  assign n32830 = ~n32825 & ~P3_EAX_REG_2__SCAN_IN;
  assign n32828 = ~n35462 | ~BUF2_REG_2__SCAN_IN;
  assign n32827 = ~n32826 | ~n36333;
  assign n32829 = ~n32828 | ~n32827;
  assign n32831 = ~n32830 & ~n32829;
  assign P3_U2733 = ~n32832 | ~n32831;
  assign n32836 = ~n35459 & ~n32833;
  assign n32835 = ~n32834 & ~n34843;
  assign n32842 = ~n32836 & ~n32835;
  assign n32837 = ~P3_EAX_REG_9__SCAN_IN | ~n36243;
  assign n32840 = ~n32837 | ~n32838;
  assign n33225 = ~n34966;
  assign n32841 = ~n32840 | ~n33225;
  assign P3_U2726 = ~n32842 | ~n32841;
  assign n35918 = ~n35917 | ~n35916;
  assign n33925 = ~P3_EBX_REG_3__SCAN_IN & ~n35918;
  assign n33872 = ~P3_EBX_REG_4__SCAN_IN;
  assign n33873 = ~n33925 | ~n33872;
  assign n33765 = ~P3_EBX_REG_5__SCAN_IN & ~n33873;
  assign n33764 = ~P3_EBX_REG_6__SCAN_IN;
  assign n33766 = ~n33765 | ~n33764;
  assign n33621 = ~P3_EBX_REG_7__SCAN_IN & ~n33766;
  assign n33739 = ~P3_EBX_REG_12__SCAN_IN;
  assign n36176 = ~P3_EBX_REG_18__SCAN_IN;
  assign n37324 = ~P3_EBX_REG_20__SCAN_IN;
  assign n40544 = ~P3_EBX_REG_24__SCAN_IN;
  assign n32851 = ~n33801 & ~n40544;
  assign n32866 = ~n41375 & ~P3_STATEBS16_REG_SCAN_IN;
  assign n32847 = ~n35452 & ~n32843;
  assign n34626 = ~n32847 & ~n32846;
  assign n35642 = ~P3_EBX_REG_31__SCAN_IN | ~n34611;
  assign n32850 = ~n35944 | ~n33906;
  assign n32879 = ~n32851 & ~n32850;
  assign n32852 = ~n35979 & ~n35904;
  assign n33870 = ~P3_REIP_REG_3__SCAN_IN | ~n32852;
  assign n33106 = ~n36966 & ~n33870;
  assign n33770 = ~P3_REIP_REG_5__SCAN_IN | ~n33106;
  assign n33516 = ~n33757 & ~n33770;
  assign n32967 = ~P3_REIP_REG_7__SCAN_IN | ~n33516;
  assign n32960 = ~n32969 & ~n32968;
  assign n33116 = ~P3_REIP_REG_10__SCAN_IN | ~n32960;
  assign n33705 = ~P3_REIP_REG_12__SCAN_IN | ~P3_REIP_REG_11__SCAN_IN;
  assign n33647 = ~n37088 & ~n33705;
  assign n33661 = ~P3_REIP_REG_14__SCAN_IN | ~n33647;
  assign n33856 = ~n33662 & ~n33661;
  assign n34546 = ~P3_REIP_REG_16__SCAN_IN | ~n33856;
  assign n32854 = ~n32853 & ~n34546;
  assign n33970 = ~P3_REIP_REG_17__SCAN_IN | ~n32854;
  assign n32855 = ~n33116 & ~n33970;
  assign n32856 = ~P3_REIP_REG_19__SCAN_IN | ~n32855;
  assign n33155 = ~n32967 & ~n32856;
  assign n33819 = ~P3_REIP_REG_20__SCAN_IN | ~n33155;
  assign n33594 = ~n33821 & ~n33819;
  assign n34625 = ~P3_REIP_REG_22__SCAN_IN | ~n33594;
  assign n32872 = ~n37757 & ~n34625;
  assign n32862 = ~n32872;
  assign n33923 = ~n32861 | ~n32860;
  assign n33891 = ~n33772 | ~n33900;
  assign n32864 = ~n32862 & ~n33891;
  assign n39426 = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n32863 = ~n39426 & ~n35947;
  assign n32877 = ~n32864 & ~n32863;
  assign n41325 = n32867 & n32866;
  assign n32869 = ~n32868;
  assign n35945 = ~n32871 & ~n36153;
  assign n32875 = ~n40544 & ~n35945;
  assign n32873 = ~n32872 & ~n33923;
  assign n33892 = ~n32873 & ~n34626;
  assign n32874 = ~n33900 & ~n33892;
  assign n32876 = ~n32875 & ~n32874;
  assign n32878 = ~n32877 | ~n32876;
  assign n32888 = ~n32879 & ~n32878;
  assign n37758 = ~P3_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n33945 = ~P3_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n32975 = ~n36963 & ~n36918;
  assign n35995 = ~n36659 | ~n32975;
  assign n35997 = P3_PHYADDRPOINTER_REG_6__SCAN_IN & P3_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n32976 = ~n35997 | ~P3_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n35842 = ~n36439 & ~n36433;
  assign n32882 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN | ~P3_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n37578 = ~n37575 | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n33835 = ~n37577 & ~n37578;
  assign n33602 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN | ~n33835;
  assign n33601 = ~P3_PHYADDRPOINTER_REG_0__SCAN_IN & ~n33602;
  assign n33814 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN | ~n33601;
  assign n32884 = ~n37758 & ~n33814;
  assign n41092 = ~P3_PHYADDRPOINTER_REG_27__SCAN_IN | ~P3_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n38910 = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN | ~P3_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n35939 = n41518 | n41402;
  assign n41401 = ~P3_PHYADDRPOINTER_REG_31__SCAN_IN ^ n35939;
  assign n32885 = ~n32884 & ~n34979;
  assign n33894 = n38909 | n36220;
  assign n39425 = ~n39426 ^ n33894;
  assign n32886 = ~n32885 ^ n39425;
  assign n35942 = ~P3_STATE2_REG_1__SCAN_IN | ~n33496;
  assign n32887 = ~n32886 | ~n35930;
  assign P3_U2647 = ~n32888 | ~n32887;
  assign n40311 = n32890 ^ n32889;
  assign n32899 = ~n40311 & ~n39522;
  assign n32897 = ~n37637 | ~n34909;
  assign n32898 = ~n40325 & ~n32897;
  assign n32903 = ~n32899 & ~n32898;
  assign n32901 = ~n32900 | ~n34901;
  assign n32902 = ~n40325 | ~n32901;
  assign n32904 = ~n32903 | ~n32902;
  assign n32906 = ~n34913 | ~n32904;
  assign n32905 = ~n34914 | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign P2_U3603 = ~n32906 | ~n32905;
  assign n32908 = ~n36298 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n32907 = ~n36307 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n32912 = ~n32908 | ~n32907;
  assign n32910 = ~n22919 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n32909 = ~n36320 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n32911 = ~n32910 | ~n32909;
  assign n32920 = ~n32912 & ~n32911;
  assign n32914 = ~n22903 | ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n32913 = ~n36317 | ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n32918 = ~n32914 | ~n32913;
  assign n32916 = ~n22914 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n32915 = ~n36311 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n32917 = ~n32916 | ~n32915;
  assign n32919 = ~n32918 & ~n32917;
  assign n32936 = ~n32920 | ~n32919;
  assign n32922 = ~n22902 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n32921 = ~n22917 | ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n32926 = ~n32922 | ~n32921;
  assign n32924 = ~n22910 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n32923 = ~n35392 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n32925 = ~n32924 | ~n32923;
  assign n32934 = ~n32926 & ~n32925;
  assign n32928 = ~n36294 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n32927 = ~n22913 | ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n32932 = ~n32928 | ~n32927;
  assign n32930 = ~n22923 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n32929 = ~n22920 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n32931 = ~n32930 | ~n32929;
  assign n32933 = ~n32932 & ~n32931;
  assign n32935 = ~n32934 | ~n32933;
  assign n34842 = ~n32936 & ~n32935;
  assign n32941 = n34842 | n43930;
  assign n32937 = ~P3_EBX_REG_12__SCAN_IN | ~n43930;
  assign n32939 = ~n32937 | ~n32938;
  assign n33260 = ~n33262;
  assign n32940 = ~n32939 | ~n33260;
  assign P3_U2691 = ~n32941 | ~n32940;
  assign n34869 = n32943 ^ n32942;
  assign n32947 = ~n43913 | ~n34869;
  assign n34853 = n32945 ^ n32944;
  assign n32946 = ~n43809 | ~n34853;
  assign n32951 = ~n32947 | ~n32946;
  assign n32949 = ~n40320 | ~n43896;
  assign n32948 = ~n43917 | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n32950 = ~n32949 | ~n32948;
  assign n32955 = ~n32951 & ~n32950;
  assign n35720 = ~n40306;
  assign n32953 = ~n43915 & ~n35720;
  assign n32952 = P2_REIP_REG_2__SCAN_IN & n43880;
  assign n32954 = ~n32953 & ~n32952;
  assign P2_U3012 = ~n32955 | ~n32954;
  assign n32956 = ~n23700 | ~n23415;
  assign n32957 = ~n32956 | ~n38820;
  assign n32959 = ~n32957 | ~n43525;
  assign n32958 = ~P2_EBX_REG_3__SCAN_IN | ~n35967;
  assign P2_U2884 = ~n32959 | ~n32958;
  assign n32961 = ~n32969 & ~n35951;
  assign n33073 = ~n32960 | ~n33630;
  assign n32965 = ~n32961 | ~n33073;
  assign n32963 = ~n33067 & ~n35642;
  assign n32962 = ~P3_EBX_REG_9__SCAN_IN | ~n33622;
  assign n32964 = ~n32963 | ~n32962;
  assign n32982 = ~n32965 | ~n32964;
  assign n34990 = ~n34626 & ~n32966;
  assign n32972 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN | ~n36154;
  assign n33619 = n33923 | n32967;
  assign n32970 = ~n32968 & ~n33619;
  assign n32971 = ~n32970 | ~n32969;
  assign n32973 = ~n32972 | ~n32971;
  assign n32980 = ~n34990 & ~n32973;
  assign n33944 = ~P3_PHYADDRPOINTER_REG_2__SCAN_IN | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n32974 = ~n33945 & ~n33944;
  assign n33866 = ~P3_PHYADDRPOINTER_REG_4__SCAN_IN | ~n32974;
  assign n33758 = ~n36918 & ~n33866;
  assign n33529 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN | ~n33758;
  assign n33759 = ~n33529;
  assign n33615 = P3_PHYADDRPOINTER_REG_7__SCAN_IN & n33759;
  assign n33077 = ~P3_PHYADDRPOINTER_REG_8__SCAN_IN | ~n33615;
  assign n36411 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN ^ n33077;
  assign n33947 = ~n32974;
  assign n33867 = ~P3_PHYADDRPOINTER_REG_0__SCAN_IN & ~n33947;
  assign n33761 = ~n32975 | ~n33867;
  assign n32977 = ~n32976 & ~n33761;
  assign n33080 = ~n32977 & ~n34979;
  assign n32978 = n36411 ^ n33080;
  assign n32979 = ~n35930 | ~n32978;
  assign n32981 = ~n32980 | ~n32979;
  assign n32984 = ~n32982 & ~n32981;
  assign n32983 = ~P3_EBX_REG_9__SCAN_IN | ~n35935;
  assign P3_U2662 = ~n32984 | ~n32983;
  assign n34013 = ~n43972 & ~n33062;
  assign n32988 = ~n33062;
  assign n32987 = ~n43972 & ~n34968;
  assign n32989 = ~n32988 & ~n32987;
  assign n33023 = ~n34013 & ~n32989;
  assign n33021 = ~BUF2_REG_20__SCAN_IN | ~n36282;
  assign n33141 = ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n32991 = n22921 | n33141;
  assign n32990 = ~n22902 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n32995 = ~n32991 | ~n32990;
  assign n32993 = ~n22914 | ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n32992 = ~n35392 | ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n32994 = ~n32993 | ~n32992;
  assign n32999 = n32995 | n32994;
  assign n32997 = ~n22919 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n32996 = ~n22923 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n32998 = ~n32997 | ~n32996;
  assign n33019 = ~n32999 & ~n32998;
  assign n33001 = ~n36317 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n33000 = ~n36307 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n33005 = ~n33001 | ~n33000;
  assign n33003 = ~n36310 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n33002 = ~n36311 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n33004 = ~n33003 | ~n33002;
  assign n33013 = ~n33005 & ~n33004;
  assign n33007 = ~n22903 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n33006 = ~n22909 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n33011 = ~n33007 | ~n33006;
  assign n33009 = ~n22917 | ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n33008 = ~n36320 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n33010 = ~n33009 | ~n33008;
  assign n33012 = ~n33011 & ~n33010;
  assign n33017 = ~n33013 | ~n33012;
  assign n33015 = ~n36294 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n33014 = ~n22913 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n33016 = ~n33015 | ~n33014;
  assign n33018 = ~n33017 & ~n33016;
  assign n37322 = ~n33019 | ~n33018;
  assign n33020 = ~n36333 | ~n37322;
  assign n33022 = ~n33021 | ~n33020;
  assign n33025 = ~n33023 & ~n33022;
  assign n33024 = ~n36338 | ~BUF2_REG_4__SCAN_IN;
  assign P3_U2715 = ~n33025 | ~n33024;
  assign n33060 = BUF2_REG_19__SCAN_IN & n36282;
  assign n33058 = ~BUF2_REG_3__SCAN_IN | ~n36338;
  assign n33027 = ~n22920 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n33026 = ~n36311 | ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n33030 = ~n33027 | ~n33026;
  assign n33028 = ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n33029 = ~n34042 & ~n33028;
  assign n33032 = ~n33030 & ~n33029;
  assign n33031 = ~n36294 | ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n33036 = ~n33032 | ~n33031;
  assign n33034 = ~n22913 | ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n33033 = ~n36307 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n33035 = ~n33034 | ~n33033;
  assign n33056 = ~n33036 & ~n33035;
  assign n33038 = ~n22919 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n33037 = ~n22903 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n33042 = ~n33038 | ~n33037;
  assign n33040 = ~n36310 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n33039 = ~n22923 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n33041 = ~n33040 | ~n33039;
  assign n33050 = ~n33042 & ~n33041;
  assign n33044 = ~n22902 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n33043 = ~n36317 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n33048 = ~n33044 | ~n33043;
  assign n33046 = ~n22914 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n33045 = ~n22917 | ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n33047 = ~n33046 | ~n33045;
  assign n33049 = ~n33048 & ~n33047;
  assign n33054 = ~n33050 | ~n33049;
  assign n33052 = ~n35392 | ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n33051 = ~n36320 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n33053 = ~n33052 | ~n33051;
  assign n33055 = ~n33054 & ~n33053;
  assign n36400 = ~n33056 | ~n33055;
  assign n33057 = ~n36333 | ~n36400;
  assign n33059 = ~n33058 | ~n33057;
  assign n33065 = ~n33060 & ~n33059;
  assign n33061 = ~P3_EAX_REG_19__SCAN_IN | ~n36243;
  assign n33266 = ~P3_EAX_REG_18__SCAN_IN | ~n33268;
  assign n33063 = ~n33061 | ~n33266;
  assign n33064 = ~n33063 | ~n33062;
  assign P3_U2716 = ~n33065 | ~n33064;
  assign n33069 = ~n33067 & ~n33066;
  assign n33068 = ~n35944 | ~n33124;
  assign n33070 = ~n33069 & ~n33068;
  assign n33072 = ~n33070 & ~n34990;
  assign n33071 = ~n36154 | ~P3_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n33087 = ~n33072 | ~n33071;
  assign n33076 = ~n33074 | ~n33073;
  assign n33075 = ~n33116;
  assign n33672 = ~n34536;
  assign n33131 = ~n35951 & ~n33672;
  assign n33085 = ~n33076 | ~n33131;
  assign n36412 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n33078 = ~n36412 & ~n33077;
  assign n33079 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN & ~n33078;
  assign n33119 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN | ~n33078;
  assign n33117 = ~n33119;
  assign n36460 = ~n33079 & ~n33117;
  assign n33081 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN & ~n34979;
  assign n33082 = ~n33081 & ~n33080;
  assign n33083 = ~n36460 ^ n33082;
  assign n33084 = ~n33083 | ~n35930;
  assign n33086 = ~n33085 | ~n33084;
  assign n33089 = ~n33087 & ~n33086;
  assign n33088 = ~P3_EBX_REG_10__SCAN_IN | ~n35935;
  assign P3_U2661 = ~n33089 | ~n33088;
  assign n33092 = ~P3_EAX_REG_0__SCAN_IN | ~n33090;
  assign n33091 = ~n35462 | ~BUF2_REG_0__SCAN_IN;
  assign n33093 = ~n33092 | ~n33091;
  assign n33097 = ~n33094 & ~n33093;
  assign n33096 = ~n33095 | ~n36333;
  assign P3_U2735 = ~n33097 | ~n33096;
  assign n33098 = ~n33923 & ~P3_REIP_REG_5__SCAN_IN;
  assign n33102 = ~n33098 | ~n33106;
  assign n33100 = ~n33765 & ~n35642;
  assign n33099 = ~P3_EBX_REG_5__SCAN_IN | ~n33873;
  assign n33101 = ~n33100 | ~n33099;
  assign n33103 = ~n33102 | ~n33101;
  assign n33105 = ~n34990 & ~n33103;
  assign n33104 = ~n36154 | ~P3_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n33110 = ~n33105 | ~n33104;
  assign n33108 = ~P3_EBX_REG_5__SCAN_IN | ~n35935;
  assign n33871 = n33106 | n33923;
  assign n33888 = ~n33496 | ~n33871;
  assign n33107 = ~P3_REIP_REG_5__SCAN_IN | ~n33888;
  assign n33109 = ~n33108 | ~n33107;
  assign n33115 = ~n33110 & ~n33109;
  assign n33111 = ~n33866 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n33112 = ~n33111 & ~n34979;
  assign n36915 = ~n36918 ^ n33866;
  assign n33113 = ~n33112 ^ n36915;
  assign n33114 = ~n35930 | ~n33113;
  assign P3_U2666 = ~n33115 | ~n33114;
  assign n33135 = ~P3_REIP_REG_11__SCAN_IN & ~n34545;
  assign n33118 = ~P3_PHYADDRPOINTER_REG_11__SCAN_IN & ~n33117;
  assign n35849 = ~n36439 & ~n33119;
  assign n36436 = ~n33118 & ~n35849;
  assign n33120 = ~n33119 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n33121 = ~n33120 & ~n34979;
  assign n33122 = ~n36436 ^ n33121;
  assign n33130 = ~n33122 & ~n35942;
  assign n33123 = ~n35947 & ~n36439;
  assign n33128 = ~n33123 & ~n34990;
  assign n33126 = ~n33738 & ~n35642;
  assign n33125 = ~P3_EBX_REG_11__SCAN_IN | ~n33124;
  assign n33127 = ~n33126 | ~n33125;
  assign n33129 = ~n33128 | ~n33127;
  assign n33133 = ~n33130 & ~n33129;
  assign n33132 = ~P3_REIP_REG_11__SCAN_IN | ~n33131;
  assign n33134 = ~n33133 | ~n33132;
  assign n33137 = ~n33135 & ~n33134;
  assign n33136 = ~P3_EBX_REG_11__SCAN_IN | ~n35935;
  assign P3_U2660 = ~n33137 | ~n33136;
  assign n33138 = ~n33872 & ~n42135;
  assign n33162 = ~P3_EBX_REG_2__SCAN_IN | ~n43932;
  assign n33164 = ~P3_EBX_REG_3__SCAN_IN | ~n43933;
  assign n33145 = ~n33138 | ~n33164;
  assign n33140 = ~n33139 | ~n43932;
  assign n33143 = ~n33140 & ~P3_EBX_REG_4__SCAN_IN;
  assign n33142 = ~n33141 & ~n43930;
  assign n33144 = ~n33143 & ~n33142;
  assign P3_U2699 = ~n33145 | ~n33144;
  assign n37584 = ~P3_PHYADDRPOINTER_REG_20__SCAN_IN ^ n37578;
  assign n33836 = ~P3_PHYADDRPOINTER_REG_0__SCAN_IN & ~n37578;
  assign n33146 = ~n33836 & ~n34979;
  assign n33147 = ~n37584 ^ n33146;
  assign n33151 = ~n35942 & ~n33147;
  assign n33149 = ~P3_PHYADDRPOINTER_REG_20__SCAN_IN | ~n36154;
  assign n33148 = ~P3_EBX_REG_20__SCAN_IN | ~n35935;
  assign n33150 = ~n33149 | ~n33148;
  assign n33161 = ~n33151 & ~n33150;
  assign n33153 = ~n33953 & ~n37324;
  assign n33152 = ~n35944 | ~n33824;
  assign n33159 = ~n33153 & ~n33152;
  assign n33154 = n33819 & n33772;
  assign n33822 = ~n33154 & ~n34626;
  assign n33156 = n33772 & n33155;
  assign n33157 = ~P3_REIP_REG_20__SCAN_IN & ~n33156;
  assign n33158 = ~n33822 & ~n33157;
  assign n33160 = ~n33159 & ~n33158;
  assign P3_U2651 = ~n33161 | ~n33160;
  assign n33167 = ~P3_INSTQUEUE_REG_0__3__SCAN_IN | ~n42135;
  assign n33165 = ~n33163 | ~n33162;
  assign n33166 = ~n33165 | ~n33164;
  assign P3_U2700 = ~n33167 | ~n33166;
  assign n33205 = BUF2_REG_26__SCAN_IN & n36282;
  assign n34329 = ~n33169 & ~n33168;
  assign n33171 = ~n22919 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n33170 = ~n22913 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n33175 = ~n33171 | ~n33170;
  assign n33173 = ~n36298 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n33172 = ~n22914 | ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n33174 = ~n33173 | ~n33172;
  assign n33201 = ~n33175 & ~n33174;
  assign n33177 = ~n36310 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n33176 = ~n22917 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n33181 = ~n33177 | ~n33176;
  assign n33179 = ~n36320 | ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n33178 = ~n36311 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n33180 = ~n33179 | ~n33178;
  assign n33189 = ~n33181 & ~n33180;
  assign n33183 = ~n22903 | ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n33182 = ~n36317 | ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n33187 = ~n33183 | ~n33182;
  assign n33185 = ~n22902 | ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n33184 = ~n36307 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n33186 = ~n33185 | ~n33184;
  assign n33188 = ~n33187 & ~n33186;
  assign n33199 = ~n33189 | ~n33188;
  assign n33190 = ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n33195 = ~n33191 & ~n33190;
  assign n33193 = ~n22923 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n33192 = ~n22920 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n33194 = ~n33193 | ~n33192;
  assign n33197 = ~n33195 & ~n33194;
  assign n33196 = ~n36294 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n33198 = ~n33197 | ~n33196;
  assign n33200 = ~n33199 & ~n33198;
  assign n34328 = ~n33201 | ~n33200;
  assign n41065 = n34329 ^ n34328;
  assign n33203 = ~n36333 | ~n41065;
  assign n33202 = ~n36338 | ~BUF2_REG_10__SCAN_IN;
  assign n33204 = ~n33203 | ~n33202;
  assign n33211 = ~n33205 & ~n33204;
  assign n33207 = ~P3_EAX_REG_26__SCAN_IN | ~n36243;
  assign n33209 = ~n33207 | ~n33206;
  assign n33210 = ~n33209 | ~n34335;
  assign P3_U2709 = ~n33211 | ~n33210;
  assign n33215 = ~n43695 & ~n40311;
  assign n33213 = ~P2_EAX_REG_2__SCAN_IN | ~n43698;
  assign n33212 = ~n36955 | ~n38018;
  assign n33214 = ~n33213 | ~n33212;
  assign n33220 = ~n33215 & ~n33214;
  assign n36003 = n37638 ^ n40311;
  assign n36004 = ~n33217 & ~n33216;
  assign n33218 = ~n36003 ^ n36004;
  assign n33219 = ~n33218 | ~n43693;
  assign P2_U2917 = ~n33220 | ~n33219;
  assign n33224 = ~n35459 & ~n33221;
  assign n33223 = ~n33222 & ~n34843;
  assign n33229 = ~n33224 & ~n33223;
  assign n33226 = ~P3_EAX_REG_10__SCAN_IN | ~n36243;
  assign n33227 = ~n33226 | ~n33225;
  assign n33228 = ~n33227 | ~n34355;
  assign P3_U2725 = ~n33229 | ~n33228;
  assign n33231 = ~n22909 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n33230 = ~n36310 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n33235 = ~n33231 | ~n33230;
  assign n33233 = ~n22919 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n33232 = ~n22912 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n33234 = ~n33233 | ~n33232;
  assign n33243 = ~n33235 & ~n33234;
  assign n33237 = ~n22903 | ~P3_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n33236 = ~n36317 | ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n33241 = ~n33237 | ~n33236;
  assign n33239 = ~n22923 | ~P3_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n33238 = ~n36311 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n33240 = ~n33239 | ~n33238;
  assign n33242 = ~n33241 & ~n33240;
  assign n33259 = ~n33243 | ~n33242;
  assign n33245 = ~n22913 | ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n33244 = ~n35392 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n33249 = ~n33245 | ~n33244;
  assign n33247 = ~n22902 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n33246 = ~n22914 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n33248 = ~n33247 | ~n33246;
  assign n33257 = ~n33249 & ~n33248;
  assign n33251 = ~n22917 | ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n33250 = ~n36307 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n33255 = ~n33251 | ~n33250;
  assign n33253 = ~n36294 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n33252 = ~n36320 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n33254 = ~n33253 | ~n33252;
  assign n33256 = ~n33255 & ~n33254;
  assign n33258 = ~n33257 | ~n33256;
  assign n35458 = ~n33259 & ~n33258;
  assign n33265 = n35458 | n43930;
  assign n33261 = ~P3_EBX_REG_13__SCAN_IN | ~n43930;
  assign n33263 = ~n33261 | ~n33260;
  assign n34401 = ~n33262 | ~P3_EBX_REG_13__SCAN_IN;
  assign n33264 = ~n33263 | ~n34401;
  assign P3_U2690 = ~n33265 | ~n33264;
  assign n33270 = ~n33266;
  assign n33267 = ~n43977 & ~n34968;
  assign n33269 = ~n33268 & ~n33267;
  assign n33274 = ~n33270 & ~n33269;
  assign n33272 = ~n36282 | ~BUF2_REG_18__SCAN_IN;
  assign n33271 = ~n36338 | ~BUF2_REG_2__SCAN_IN;
  assign n33273 = ~n33272 | ~n33271;
  assign n33308 = ~n33274 & ~n33273;
  assign n33276 = ~n36307 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n33275 = ~n35392 | ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n33280 = ~n33276 | ~n33275;
  assign n33278 = ~n22919 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n33277 = ~n22923 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n33279 = ~n33278 | ~n33277;
  assign n33306 = ~n33280 & ~n33279;
  assign n33282 = ~n22917 | ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n33281 = ~n36311 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n33286 = ~n33282 | ~n33281;
  assign n33284 = ~n22909 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n33283 = ~n22914 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n33285 = ~n33284 | ~n33283;
  assign n33294 = ~n33286 & ~n33285;
  assign n33288 = ~n22903 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n33287 = ~n36317 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n33292 = ~n33288 | ~n33287;
  assign n33290 = ~n36310 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n33289 = ~n36320 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n33291 = ~n33290 | ~n33289;
  assign n33293 = ~n33292 & ~n33291;
  assign n33304 = ~n33294 | ~n33293;
  assign n33296 = n22901 | n43931;
  assign n33295 = ~n22902 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n33300 = ~n33296 | ~n33295;
  assign n33297 = ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n33299 = ~n33298 & ~n33297;
  assign n33302 = ~n33300 & ~n33299;
  assign n33301 = ~n36294 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n33303 = ~n33302 | ~n33301;
  assign n33305 = ~n33304 & ~n33303;
  assign n36174 = ~n33306 | ~n33305;
  assign n33307 = ~n36333 | ~n36174;
  assign P3_U2717 = ~n33308 | ~n33307;
  assign n33312 = ~n33792;
  assign n33311 = ~n33310 | ~n33309;
  assign n35869 = ~n33312 | ~n33311;
  assign n33319 = ~n35869 & ~n43298;
  assign n33316 = ~n33313;
  assign n33315 = ~n33314;
  assign n33317 = ~n33316 | ~n33315;
  assign n33318 = ~n34063 & ~n44019;
  assign n33321 = ~n33319 & ~n33318;
  assign n33320 = ~P1_EBX_REG_3__SCAN_IN | ~n44023;
  assign P1_U2869 = ~n33321 | ~n33320;
  assign n33322 = ~n34400 & ~n42135;
  assign n33356 = ~n33322 | ~n34401;
  assign n33354 = ~n34401 & ~P3_EBX_REG_14__SCAN_IN;
  assign n33324 = ~n36294 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n33323 = ~n36311 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n33328 = ~n33324 | ~n33323;
  assign n33326 = ~n22914 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n33325 = ~n36307 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n33327 = ~n33326 | ~n33325;
  assign n33336 = ~n33328 & ~n33327;
  assign n33330 = ~n22903 | ~P3_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n33329 = ~n36317 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n33334 = ~n33330 | ~n33329;
  assign n33332 = ~n36310 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n33331 = ~n22913 | ~P3_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n33333 = ~n33332 | ~n33331;
  assign n33335 = ~n33334 & ~n33333;
  assign n33352 = ~n33336 | ~n33335;
  assign n33338 = ~n22919 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n33337 = ~n35392 | ~P3_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n33342 = ~n33338 | ~n33337;
  assign n33340 = ~n22909 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n33339 = ~n22920 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n33341 = ~n33340 | ~n33339;
  assign n33350 = ~n33342 & ~n33341;
  assign n33344 = ~n22902 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n33343 = ~n22917 | ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n33348 = ~n33344 | ~n33343;
  assign n33346 = ~n36320 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n33345 = ~n22923 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n33347 = ~n33346 | ~n33345;
  assign n33349 = ~n33348 & ~n33347;
  assign n33351 = ~n33350 | ~n33349;
  assign n34965 = ~n33352 & ~n33351;
  assign n33353 = ~n43930 & ~n34965;
  assign n33355 = ~n33354 & ~n33353;
  assign P3_U2689 = ~n33356 | ~n33355;
  assign n33544 = ~n33357 & ~n33545;
  assign n33359 = ~n33544 | ~P2_EAX_REG_29__SCAN_IN;
  assign n33358 = ~n33545 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n33361 = n33359 & n33358;
  assign n33360 = ~n33548 | ~P2_UWORD_REG_13__SCAN_IN;
  assign P2_U2922 = ~n33361 | ~n33360;
  assign n33363 = ~n33544 | ~P2_EAX_REG_28__SCAN_IN;
  assign n33362 = ~n33545 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n33365 = n33363 & n33362;
  assign n33364 = ~n33548 | ~P2_UWORD_REG_12__SCAN_IN;
  assign P2_U2923 = ~n33365 | ~n33364;
  assign n33367 = ~n33544 | ~P2_EAX_REG_27__SCAN_IN;
  assign n33366 = ~n33545 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n33369 = n33367 & n33366;
  assign n33368 = ~n33548 | ~P2_UWORD_REG_11__SCAN_IN;
  assign P2_U2924 = ~n33369 | ~n33368;
  assign n33371 = ~n33544 | ~P2_EAX_REG_26__SCAN_IN;
  assign n33370 = ~n33545 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n33373 = n33371 & n33370;
  assign n33372 = ~n33548 | ~P2_UWORD_REG_10__SCAN_IN;
  assign P2_U2925 = ~n33373 | ~n33372;
  assign n33375 = ~n33544 | ~P2_EAX_REG_25__SCAN_IN;
  assign n33374 = ~n33545 | ~P2_DATAO_REG_25__SCAN_IN;
  assign n33377 = n33375 & n33374;
  assign n33376 = ~n33548 | ~P2_UWORD_REG_9__SCAN_IN;
  assign P2_U2926 = ~n33377 | ~n33376;
  assign n33379 = ~n33545 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n33378 = ~n33544 | ~P2_EAX_REG_24__SCAN_IN;
  assign n33381 = n33379 & n33378;
  assign n33380 = ~n33548 | ~P2_UWORD_REG_8__SCAN_IN;
  assign P2_U2927 = ~n33381 | ~n33380;
  assign n33383 = ~n33544 | ~P2_EAX_REG_23__SCAN_IN;
  assign n33382 = ~n33545 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n33385 = n33383 & n33382;
  assign n33384 = ~n33548 | ~P2_UWORD_REG_7__SCAN_IN;
  assign P2_U2928 = ~n33385 | ~n33384;
  assign n33387 = ~n33544 | ~P2_EAX_REG_22__SCAN_IN;
  assign n33386 = ~n33545 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n33389 = n33387 & n33386;
  assign n33388 = ~n33548 | ~P2_UWORD_REG_6__SCAN_IN;
  assign P2_U2929 = ~n33389 | ~n33388;
  assign n33391 = ~n33544 | ~P2_EAX_REG_21__SCAN_IN;
  assign n33390 = ~n33545 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n33393 = n33391 & n33390;
  assign n33392 = ~n33548 | ~P2_UWORD_REG_5__SCAN_IN;
  assign P2_U2930 = ~n33393 | ~n33392;
  assign n33395 = ~n33544 | ~P2_EAX_REG_20__SCAN_IN;
  assign n33394 = ~n33545 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n33397 = n33395 & n33394;
  assign n33396 = ~n33548 | ~P2_UWORD_REG_4__SCAN_IN;
  assign P2_U2931 = ~n33397 | ~n33396;
  assign n33399 = ~n33545 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n33398 = ~n33544 | ~P2_EAX_REG_19__SCAN_IN;
  assign n33401 = n33399 & n33398;
  assign n33400 = ~n33548 | ~P2_UWORD_REG_3__SCAN_IN;
  assign P2_U2932 = ~n33401 | ~n33400;
  assign n33403 = ~n33544 | ~P2_EAX_REG_18__SCAN_IN;
  assign n33402 = ~n33545 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n33405 = n33403 & n33402;
  assign n33404 = ~n33548 | ~P2_UWORD_REG_2__SCAN_IN;
  assign P2_U2933 = ~n33405 | ~n33404;
  assign n33407 = ~n33544 | ~P2_EAX_REG_17__SCAN_IN;
  assign n33406 = ~n33545 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n33409 = n33407 & n33406;
  assign n33408 = ~n33548 | ~P2_UWORD_REG_1__SCAN_IN;
  assign P2_U2934 = ~n33409 | ~n33408;
  assign n33411 = ~n33544 | ~P2_EAX_REG_16__SCAN_IN;
  assign n33410 = ~n33545 | ~P2_DATAO_REG_16__SCAN_IN;
  assign n33413 = n33411 & n33410;
  assign n33412 = ~n33548 | ~P2_UWORD_REG_0__SCAN_IN;
  assign P2_U2935 = ~n33413 | ~n33412;
  assign n33415 = ~P2_EAX_REG_15__SCAN_IN | ~n33474;
  assign n33414 = ~n33545 | ~P2_DATAO_REG_15__SCAN_IN;
  assign n33417 = n33415 & n33414;
  assign n33416 = ~n33548 | ~P2_LWORD_REG_15__SCAN_IN;
  assign P2_U2936 = ~n33417 | ~n33416;
  assign n33419 = ~P2_EAX_REG_14__SCAN_IN | ~n33474;
  assign n33418 = ~n33545 | ~P2_DATAO_REG_14__SCAN_IN;
  assign n33421 = n33419 & n33418;
  assign n33420 = ~n33548 | ~P2_LWORD_REG_14__SCAN_IN;
  assign P2_U2937 = ~n33421 | ~n33420;
  assign n33423 = ~n33545 | ~P2_DATAO_REG_13__SCAN_IN;
  assign n33422 = ~P2_EAX_REG_13__SCAN_IN | ~n33474;
  assign n33425 = n33423 & n33422;
  assign P2_U2938 = ~n33425 | ~n33424;
  assign n33427 = ~P2_EAX_REG_12__SCAN_IN | ~n33474;
  assign n33426 = ~n33545 | ~P2_DATAO_REG_12__SCAN_IN;
  assign n33429 = n33427 & n33426;
  assign P2_U2939 = ~n33429 | ~n33428;
  assign n33431 = ~n33545 | ~P2_DATAO_REG_11__SCAN_IN;
  assign n33430 = ~P2_EAX_REG_11__SCAN_IN | ~n33474;
  assign n33433 = n33431 & n33430;
  assign P2_U2940 = ~n33433 | ~n33432;
  assign n33435 = ~n33545 | ~P2_DATAO_REG_10__SCAN_IN;
  assign n33434 = ~P2_EAX_REG_10__SCAN_IN | ~n33474;
  assign n33437 = n33435 & n33434;
  assign P2_U2941 = ~n33437 | ~n33436;
  assign n33439 = ~n33545 | ~P2_DATAO_REG_9__SCAN_IN;
  assign n33438 = ~P2_EAX_REG_9__SCAN_IN | ~n33474;
  assign n33441 = n33439 & n33438;
  assign P2_U2942 = ~n33441 | ~n33440;
  assign n33443 = ~n33545 | ~P2_DATAO_REG_8__SCAN_IN;
  assign n33442 = ~P2_EAX_REG_8__SCAN_IN | ~n33474;
  assign n33445 = n33443 & n33442;
  assign P2_U2943 = ~n33445 | ~n33444;
  assign n33447 = ~P2_EAX_REG_7__SCAN_IN | ~n33474;
  assign n33446 = ~n33545 | ~P2_DATAO_REG_7__SCAN_IN;
  assign n33449 = n33447 & n33446;
  assign P2_U2944 = ~n33449 | ~n33448;
  assign n33451 = ~n33545 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n33450 = ~P2_EAX_REG_6__SCAN_IN | ~n33474;
  assign n33453 = n33451 & n33450;
  assign P2_U2945 = ~n33453 | ~n33452;
  assign n33455 = ~P2_EAX_REG_5__SCAN_IN | ~n33474;
  assign n33454 = ~n33545 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n33457 = n33455 & n33454;
  assign P2_U2946 = ~n33457 | ~n33456;
  assign n33459 = ~n33545 | ~P2_DATAO_REG_4__SCAN_IN;
  assign n33458 = ~P2_EAX_REG_4__SCAN_IN | ~n33474;
  assign n33461 = n33459 & n33458;
  assign P2_U2947 = ~n33461 | ~n33460;
  assign n33463 = ~n33545 | ~P2_DATAO_REG_2__SCAN_IN;
  assign n33462 = ~P2_EAX_REG_2__SCAN_IN | ~n33474;
  assign n33465 = n33463 & n33462;
  assign P2_U2949 = ~n33465 | ~n33464;
  assign n33467 = ~n33545 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n33466 = ~P2_EAX_REG_1__SCAN_IN | ~n33474;
  assign n33469 = n33467 & n33466;
  assign P2_U2950 = ~n33469 | ~n33468;
  assign n33471 = ~n33545 | ~P2_DATAO_REG_0__SCAN_IN;
  assign n33470 = ~P2_EAX_REG_0__SCAN_IN | ~n33474;
  assign n33473 = n33471 & n33470;
  assign P2_U2951 = ~n33473 | ~n33472;
  assign n33476 = ~P2_EAX_REG_3__SCAN_IN | ~n33474;
  assign n33475 = ~n33545 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n33478 = n33476 & n33475;
  assign P2_U2948 = ~n33478 | ~n33477;
  assign n33484 = ~P3_INSTQUEUE_REG_0__5__SCAN_IN | ~n42135;
  assign n33479 = n43930 & P3_EBX_REG_5__SCAN_IN;
  assign n33482 = n33480 | n33479;
  assign n33483 = ~n33482 | ~n33481;
  assign P3_U2698 = ~n33484 | ~n33483;
  assign n33485 = ~n35443 & ~n41145;
  assign n33493 = ~n33485 | ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n40743 = ~n33488 & ~n33486;
  assign n35893 = ~n35974 & ~n35975;
  assign n33491 = ~n41397 & ~n35893;
  assign n35902 = ~n41145 | ~P3_REIP_REG_0__SCAN_IN;
  assign n36914 = n33488 | n33487;
  assign n36975 = ~n36914;
  assign n33489 = ~n36975 | ~n35893;
  assign n33490 = ~n35902 | ~n33489;
  assign n33492 = ~n33491 & ~n33490;
  assign P3_U2830 = ~n33493 | ~n33492;
  assign n33495 = ~n35942 & ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n33494 = ~n41401 | ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n33499 = ~n33495 | ~n33494;
  assign n33497 = ~n35979 & ~n33496;
  assign n33930 = ~P3_REIP_REG_1__SCAN_IN & ~n33923;
  assign n33498 = ~n33497 & ~n33930;
  assign n33511 = ~n33499 | ~n33498;
  assign n34615 = ~n33501 | ~n33500;
  assign n35613 = ~n33502 | ~n36049;
  assign n33506 = ~n34615 & ~n35613;
  assign n35924 = ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n33503 = ~n36164 & ~n35924;
  assign n33504 = ~n36154 & ~n33503;
  assign n33505 = ~n36220 & ~n33504;
  assign n33509 = ~n33506 & ~n33505;
  assign n33508 = ~n35944 | ~n33507;
  assign n33510 = ~n33509 | ~n33508;
  assign n33513 = ~n33511 & ~n33510;
  assign n33512 = ~P3_EBX_REG_1__SCAN_IN | ~n35935;
  assign P3_U2670 = ~n33513 | ~n33512;
  assign n33526 = ~n33515 & ~n33756;
  assign n33517 = ~n33923 & ~P3_REIP_REG_7__SCAN_IN;
  assign n33521 = ~n33517 | ~n33516;
  assign n33519 = ~n33621 & ~n35642;
  assign n33518 = ~P3_EBX_REG_7__SCAN_IN | ~n33766;
  assign n33520 = ~n33519 | ~n33518;
  assign n33522 = ~n33521 | ~n33520;
  assign n33524 = ~n34990 & ~n33522;
  assign n33523 = ~n36154 | ~P3_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n33525 = ~n33524 | ~n33523;
  assign n33536 = ~n33526 & ~n33525;
  assign n33534 = ~n33527 & ~n35945;
  assign n33528 = ~P3_PHYADDRPOINTER_REG_7__SCAN_IN & ~n33759;
  assign n35986 = ~n33528 & ~n33615;
  assign n33530 = ~n33529 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n33531 = ~n33530 & ~n34979;
  assign n33532 = ~n35986 ^ n33531;
  assign n33533 = ~n35942 & ~n33532;
  assign n33535 = ~n33534 & ~n33533;
  assign P3_U2664 = ~n33536 | ~n33535;
  assign n33541 = ~n43525 & ~n33537;
  assign n33539 = P2_INSTQUEUE_REG_0__6__SCAN_IN ^ n36253;
  assign n33538 = ~n43525 | ~n23415;
  assign n33540 = ~n33539 & ~n33538;
  assign n33543 = ~n33541 & ~n33540;
  assign n33542 = ~n40154 | ~n43525;
  assign P2_U2881 = ~n33543 | ~n33542;
  assign n33547 = ~n33544 | ~P2_EAX_REG_30__SCAN_IN;
  assign n33546 = ~n33545 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n33550 = n33547 & n33546;
  assign n33549 = ~P2_UWORD_REG_14__SCAN_IN | ~n33548;
  assign P2_U2921 = ~n33550 | ~n33549;
  assign n33552 = ~n34898 & ~n34166;
  assign n33551 = ~n39934 & ~n34063;
  assign n33554 = ~n33552 & ~n33551;
  assign n33553 = ~P1_EAX_REG_3__SCAN_IN | ~n43732;
  assign P1_U2901 = ~n33554 | ~n33553;
  assign n33558 = ~n33784;
  assign n33557 = ~n33556 | ~n33555;
  assign n33560 = ~n42568 & ~n33786;
  assign n33559 = ~n25738 & ~n41759;
  assign n33562 = ~n33560 & ~n33559;
  assign n33561 = ~n36955 | ~n42803;
  assign P2_U2908 = ~n33562 | ~n33561;
  assign n33565 = n33563 | P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n35784 = ~n33565 | ~n33564;
  assign n33574 = ~n43924 & ~n35784;
  assign n33568 = ~P2_PHYADDRPOINTER_REG_1__SCAN_IN & ~n43911;
  assign n33566 = ~n43813 | ~n35790;
  assign n35782 = ~P2_REIP_REG_1__SCAN_IN | ~n43880;
  assign n33567 = ~n33566 | ~n35782;
  assign n33572 = ~n33568 & ~n33567;
  assign n33570 = ~n33569 ^ P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n35785 = n33570 ^ n34880;
  assign n33571 = ~n43913 | ~n35785;
  assign n33573 = ~n33572 | ~n33571;
  assign n33576 = ~n33574 & ~n33573;
  assign n33575 = ~n43917 | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign P2_U3013 = ~n33576 | ~n33575;
  assign n33578 = ~n33577 & ~n43917;
  assign n33592 = ~n33578 & ~n37286;
  assign n33584 = ~n43915 & ~n37279;
  assign n33581 = ~n34880;
  assign n33580 = ~n37290 | ~n33579;
  assign n33582 = ~n33581 | ~n33580;
  assign n33583 = ~n43811 & ~n33582;
  assign n33590 = ~n33584 & ~n33583;
  assign n33587 = ~n33585;
  assign n33586 = ~n34885 | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n33588 = ~n33587 | ~n33586;
  assign n33589 = ~n43809 | ~n33588;
  assign n33591 = ~n33590 | ~n33589;
  assign n33593 = ~n33592 & ~n33591;
  assign n34877 = ~n43880 | ~P2_REIP_REG_0__SCAN_IN;
  assign P2_U3014 = ~n33593 | ~n34877;
  assign n33595 = ~n33923 & ~P3_REIP_REG_22__SCAN_IN;
  assign n33599 = ~n33595 | ~n33594;
  assign n33597 = ~n39502 & ~n35945;
  assign n33603 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n33596 = ~n33603 & ~n35947;
  assign n33598 = ~n33597 & ~n33596;
  assign n33610 = ~n33599 | ~n33598;
  assign n33820 = ~n33772 | ~n33821;
  assign n33600 = ~n33822 | ~n33820;
  assign n33608 = ~n33600 | ~P3_REIP_REG_22__SCAN_IN;
  assign n33605 = ~n33601 & ~n34979;
  assign n37749 = ~n37754 | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n33604 = ~n33603 | ~n33602;
  assign n38154 = ~n37749 | ~n33604;
  assign n33606 = ~n33605 ^ n38154;
  assign n33607 = ~n33606 | ~n35930;
  assign n33609 = ~n33608 | ~n33607;
  assign n33614 = ~n33610 & ~n33609;
  assign n33611 = ~n39502 & ~n33823;
  assign n33612 = ~n33611 & ~n35642;
  assign n33613 = ~n33612 | ~n33802;
  assign P3_U2649 = ~n33614 | ~n33613;
  assign n36070 = P3_PHYADDRPOINTER_REG_8__SCAN_IN ^ n33615;
  assign n33616 = ~n33615 | ~n35924;
  assign n33617 = ~n41401 | ~n33616;
  assign n33618 = n36070 ^ n33617;
  assign n33635 = ~n33618 & ~n35942;
  assign n33629 = ~P3_REIP_REG_8__SCAN_IN & ~n33619;
  assign n33624 = ~n33621 & ~n33620;
  assign n33623 = ~n35944 | ~n33622;
  assign n33625 = ~n33624 & ~n33623;
  assign n33627 = ~n33625 & ~n34990;
  assign n33626 = ~n36154 | ~P3_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n33628 = ~n33627 | ~n33626;
  assign n33633 = ~n33629 & ~n33628;
  assign n33631 = ~n35951 & ~n33630;
  assign n33632 = ~n33631 | ~P3_REIP_REG_8__SCAN_IN;
  assign n33634 = ~n33633 | ~n33632;
  assign n33637 = ~n33635 & ~n33634;
  assign n33636 = ~P3_EBX_REG_8__SCAN_IN | ~n35935;
  assign P3_U2663 = ~n33637 | ~n33636;
  assign n33653 = ~n35945 & ~n34400;
  assign n33638 = ~n33647 | ~n33951;
  assign n33645 = ~n33638 & ~P3_REIP_REG_14__SCAN_IN;
  assign n33640 = ~n33688 & ~n34400;
  assign n33639 = ~n35944 | ~n33666;
  assign n33641 = ~n33640 & ~n33639;
  assign n33643 = ~n33641 & ~n34990;
  assign n33642 = ~n36154 | ~P3_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n33644 = ~n33643 | ~n33642;
  assign n33651 = ~n33645 & ~n33644;
  assign n33649 = ~n35951 & ~n33646;
  assign n33648 = ~n33647 | ~n33672;
  assign n33650 = ~n33649 | ~n33648;
  assign n33652 = ~n33651 | ~n33650;
  assign n33660 = ~n33653 & ~n33652;
  assign n33678 = ~n36222 & ~n36220;
  assign n36212 = ~n33678;
  assign n33654 = ~P3_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n33696 = ~n36182 | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n33655 = ~n33654 | ~n33696;
  assign n36181 = ~n36212 | ~n33655;
  assign n33656 = ~n33696 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n33657 = ~n33656 & ~n34979;
  assign n33658 = ~n36181 ^ n33657;
  assign n33659 = ~n33658 | ~n35930;
  assign P3_U2657 = ~n33660 | ~n33659;
  assign n33665 = ~P3_EBX_REG_15__SCAN_IN | ~n35935;
  assign n33663 = ~n33661 & ~n34545;
  assign n33664 = ~n33663 | ~n33662;
  assign n33677 = ~n33665 | ~n33664;
  assign n33668 = ~n33848 & ~n35642;
  assign n33667 = ~P3_EBX_REG_15__SCAN_IN | ~n33666;
  assign n33670 = ~n33668 | ~n33667;
  assign n33669 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN | ~n36154;
  assign n33671 = ~n33670 | ~n33669;
  assign n33675 = ~n34990 & ~n33671;
  assign n33673 = n33856 & n33672;
  assign n33862 = ~n33673 & ~n35951;
  assign n33674 = ~P3_REIP_REG_15__SCAN_IN | ~n33862;
  assign n33676 = ~n33675 | ~n33674;
  assign n33684 = ~n33677 & ~n33676;
  assign n33679 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN & ~n33678;
  assign n33844 = ~n37694 & ~n36212;
  assign n36216 = ~n33679 & ~n33844;
  assign n33680 = ~n36212 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n33681 = ~n33680 & ~n34979;
  assign n33682 = n36216 ^ n33681;
  assign n33683 = ~n35930 | ~n33682;
  assign P3_U2656 = ~n33684 | ~n33683;
  assign n33687 = ~P3_EBX_REG_13__SCAN_IN | ~n35935;
  assign n33685 = ~n33705 & ~n34545;
  assign n33686 = ~n33685 | ~n37088;
  assign n33704 = ~n33687 | ~n33686;
  assign n33690 = ~n33688 & ~n35642;
  assign n33689 = ~P3_EBX_REG_13__SCAN_IN | ~n33741;
  assign n33692 = ~n33690 | ~n33689;
  assign n33691 = ~P3_PHYADDRPOINTER_REG_13__SCAN_IN | ~n36154;
  assign n33693 = ~n33692 | ~n33691;
  assign n33702 = ~n34990 & ~n33693;
  assign n33694 = ~P3_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n33697 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN | ~n35849;
  assign n33695 = ~n33694 | ~n33697;
  assign n37096 = ~n33696 | ~n33695;
  assign n33698 = ~n33697 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n33699 = ~n33698 & ~n34979;
  assign n33700 = ~n37096 ^ n33699;
  assign n33701 = ~n35930 | ~n33700;
  assign n33703 = ~n33702 | ~n33701;
  assign n33708 = ~n33704 & ~n33703;
  assign n33706 = ~n33705 & ~n34536;
  assign n33753 = ~n33706 & ~n35951;
  assign n33707 = ~P3_REIP_REG_13__SCAN_IN | ~n33753;
  assign P3_U2658 = ~n33708 | ~n33707;
  assign n34070 = ~n35631 | ~n33709;
  assign n38058 = n34070 & n33710;
  assign n33713 = n34495 & n33711;
  assign n33712 = ~n34495 & ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n33729 = ~n33714 & ~P1_FLUSH_REG_SCAN_IN;
  assign n33715 = ~n33729 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n33722 = ~n33729;
  assign n33723 = ~n33722 & ~n33721;
  assign n33728 = ~n33727;
  assign n33730 = ~n33729 | ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n33732 = n35623 | P1_FLUSH_REG_SCAN_IN;
  assign P1_U3032 = ~n33734 & ~n34584;
  assign n33735 = ~P3_REIP_REG_12__SCAN_IN & ~n34545;
  assign n33737 = ~P3_REIP_REG_11__SCAN_IN | ~n33735;
  assign n33736 = ~P3_EBX_REG_12__SCAN_IN | ~n35935;
  assign n33752 = ~n33737 | ~n33736;
  assign n33744 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN | ~n36154;
  assign n33740 = ~n33739 & ~n33738;
  assign n33742 = ~n33740 & ~n35642;
  assign n33743 = ~n33742 | ~n33741;
  assign n33745 = ~n33744 | ~n33743;
  assign n33750 = ~n34990 & ~n33745;
  assign n37090 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n35845 = ~n35849 ^ n37090;
  assign n33746 = n35849 & n35924;
  assign n33747 = ~n33746 & ~n34979;
  assign n33748 = n35845 ^ n33747;
  assign n33749 = ~n35930 | ~n33748;
  assign n33751 = ~n33750 | ~n33749;
  assign n33755 = ~n33752 & ~n33751;
  assign n33754 = ~P3_REIP_REG_12__SCAN_IN | ~n33753;
  assign P3_U2659 = ~n33755 | ~n33754;
  assign n33780 = ~n33757 & ~n33756;
  assign n33760 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN & ~n33758;
  assign n36026 = ~n33760 & ~n33759;
  assign n33762 = ~n41401 | ~n33761;
  assign n33763 = n36026 ^ n33762;
  assign n33776 = ~n33763 & ~n35942;
  assign n33768 = ~n33765 & ~n33764;
  assign n33767 = ~n35944 | ~n33766;
  assign n33769 = ~n33768 & ~n33767;
  assign n33774 = ~n34990 & ~n33769;
  assign n33771 = ~P3_REIP_REG_6__SCAN_IN & ~n33770;
  assign n33773 = ~n33772 | ~n33771;
  assign n33775 = ~n33774 | ~n33773;
  assign n33778 = ~n33776 & ~n33775;
  assign n33777 = ~n36154 | ~P3_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n33779 = ~n33778 | ~n33777;
  assign n33782 = ~n33780 & ~n33779;
  assign n33781 = ~P3_EBX_REG_6__SCAN_IN | ~n35935;
  assign P3_U2665 = ~n33782 | ~n33781;
  assign n33788 = ~n36002 & ~n43111;
  assign n33785 = n33784 | n33783;
  assign n33787 = ~n42309 & ~n33786;
  assign n33790 = ~n33788 & ~n33787;
  assign n33789 = ~P2_EAX_REG_12__SCAN_IN | ~n43698;
  assign P2_U2907 = ~n33790 | ~n33789;
  assign n35503 = ~n33792 ^ n33791;
  assign n33798 = ~n35503 & ~n43298;
  assign n33796 = ~n34344;
  assign n33795 = ~n33794 | ~n33793;
  assign n33797 = ~n35517 & ~n44019;
  assign n33800 = ~n33798 & ~n33797;
  assign n33799 = ~P1_EBX_REG_4__SCAN_IN | ~n44023;
  assign P1_U2868 = ~n33800 | ~n33799;
  assign n33812 = ~n35947 & ~n37758;
  assign n33808 = ~n33892 & ~n37757;
  assign n33806 = ~P3_EBX_REG_23__SCAN_IN | ~n35935;
  assign n33804 = ~n33801 & ~n35642;
  assign n33803 = ~P3_EBX_REG_23__SCAN_IN | ~n33802;
  assign n33805 = ~n33804 | ~n33803;
  assign n33807 = ~n33806 | ~n33805;
  assign n33810 = ~n33808 & ~n33807;
  assign n33809 = ~n34659 | ~n37757;
  assign n33811 = ~n33810 | ~n33809;
  assign n33818 = ~n33812 & ~n33811;
  assign n33813 = ~n37758 | ~n37749;
  assign n37760 = n33894 & n33813;
  assign n33815 = ~n41401 | ~n33814;
  assign n33816 = ~n37760 ^ n33815;
  assign n33817 = ~n33816 | ~n35930;
  assign P3_U2648 = ~n33818 | ~n33817;
  assign n33834 = ~n33820 & ~n33819;
  assign n33830 = ~n33822 & ~n33821;
  assign n33828 = ~P3_EBX_REG_21__SCAN_IN | ~n35935;
  assign n33826 = ~n33823 & ~n35642;
  assign n33825 = ~P3_EBX_REG_21__SCAN_IN | ~n33824;
  assign n33827 = ~n33826 | ~n33825;
  assign n33829 = ~n33828 | ~n33827;
  assign n33832 = ~n33830 & ~n33829;
  assign n33831 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN | ~n36154;
  assign n33833 = ~n33832 | ~n33831;
  assign n33841 = ~n33834 & ~n33833;
  assign n38178 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN ^ n33835;
  assign n33837 = ~P3_PHYADDRPOINTER_REG_20__SCAN_IN | ~n33836;
  assign n33838 = ~n41401 | ~n33837;
  assign n33839 = n38178 ^ n33838;
  assign n33840 = ~n35930 | ~n33839;
  assign P3_U2650 = ~n33841 | ~n33840;
  assign n33843 = ~P3_PHYADDRPOINTER_REG_16__SCAN_IN & ~n33844;
  assign n34526 = ~n33842 & ~n36212;
  assign n37700 = ~n33843 & ~n34526;
  assign n33845 = ~n33844 | ~n35924;
  assign n33846 = ~n41401 | ~n33845;
  assign n33847 = n37700 ^ n33846;
  assign n33861 = ~n33847 & ~n35942;
  assign n33855 = ~n35945 & ~n35420;
  assign n33850 = ~n33848 & ~n35420;
  assign n33849 = ~n35944 | ~n34531;
  assign n33851 = ~n33850 & ~n33849;
  assign n33853 = ~n33851 & ~n34990;
  assign n33852 = ~n36154 | ~P3_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n33854 = ~n33853 | ~n33852;
  assign n33859 = ~n33855 & ~n33854;
  assign n33857 = ~P3_REIP_REG_16__SCAN_IN & ~n34545;
  assign n33858 = ~n33857 | ~n33856;
  assign n33860 = ~n33859 | ~n33858;
  assign n33864 = ~n33861 & ~n33860;
  assign n33863 = ~n33862 | ~P3_REIP_REG_16__SCAN_IN;
  assign P3_U2655 = ~n33864 | ~n33863;
  assign n33865 = ~n36963 | ~n33947;
  assign n36968 = ~n33866 | ~n33865;
  assign n33868 = ~n33867 & ~n34979;
  assign n33869 = n36968 ^ n33868;
  assign n33887 = ~n33869 & ~n35942;
  assign n33877 = ~n33871 & ~n33870;
  assign n33875 = ~n33925 & ~n33872;
  assign n33874 = ~n35944 | ~n33873;
  assign n33876 = ~n33875 & ~n33874;
  assign n33885 = ~n33877 & ~n33876;
  assign n33883 = ~n36963 & ~n35947;
  assign n33878 = ~n36311 & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n33879 = ~n34615 & ~n33878;
  assign n33881 = ~n34990 & ~n33879;
  assign n33880 = ~P3_EBX_REG_4__SCAN_IN | ~n35935;
  assign n33882 = ~n33881 | ~n33880;
  assign n33884 = ~n33883 & ~n33882;
  assign n33886 = ~n33885 | ~n33884;
  assign n33890 = ~n33887 & ~n33886;
  assign n33889 = ~P3_REIP_REG_4__SCAN_IN | ~n33888;
  assign P3_U2667 = ~n33890 | ~n33889;
  assign n33893 = ~n33892 | ~n33891;
  assign n33914 = ~n33893 | ~P3_REIP_REG_25__SCAN_IN;
  assign n40733 = ~n40738 | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n33896 = ~n40733;
  assign n33897 = ~n39426 & ~n33894;
  assign n33895 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN & ~n33897;
  assign n38913 = ~n33896 & ~n33895;
  assign n33898 = n33897 & n35924;
  assign n33899 = ~n38913 ^ n34637;
  assign n33912 = ~n33899 & ~n35942;
  assign n34624 = ~n33900 & ~n37757;
  assign n33901 = ~n34624 | ~n34659;
  assign n33905 = ~n33901 & ~P3_REIP_REG_25__SCAN_IN;
  assign n33903 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN | ~n36154;
  assign n33902 = ~P3_EBX_REG_25__SCAN_IN | ~n35935;
  assign n33904 = ~n33903 | ~n33902;
  assign n33910 = ~n33905 & ~n33904;
  assign n33908 = ~n34655 & ~n35642;
  assign n33907 = ~P3_EBX_REG_25__SCAN_IN | ~n33906;
  assign n33909 = ~n33908 | ~n33907;
  assign n33911 = ~n33910 | ~n33909;
  assign n33913 = ~n33912 & ~n33911;
  assign P3_U2646 = ~n33914 | ~n33913;
  assign n33916 = ~n33915 ^ n35253;
  assign n33920 = ~n33916 & ~n33538;
  assign n41172 = ~n33918 ^ n33917;
  assign n33919 = ~n41172 & ~n35967;
  assign n33922 = ~n33920 & ~n33919;
  assign n33921 = ~P2_EBX_REG_8__SCAN_IN | ~n35967;
  assign P2_U2879 = ~n33922 | ~n33921;
  assign n33924 = ~n35904 & ~P3_REIP_REG_3__SCAN_IN;
  assign n33931 = ~n33923 & ~n35979;
  assign n33929 = ~n33924 | ~n33931;
  assign n33927 = ~n33925 & ~n35642;
  assign n33926 = ~P3_EBX_REG_3__SCAN_IN | ~n35918;
  assign n33928 = ~n33927 | ~n33926;
  assign n33942 = ~n33929 | ~n33928;
  assign n35905 = ~n34626 & ~n33930;
  assign n35914 = ~n33931 | ~n35904;
  assign n33932 = ~n35905 | ~n35914;
  assign n33940 = ~n33932 | ~P3_REIP_REG_3__SCAN_IN;
  assign n33934 = ~n36040 & ~n33933;
  assign n36058 = ~n36294 & ~n33934;
  assign n33938 = ~n34615 & ~n36058;
  assign n33936 = ~P3_PHYADDRPOINTER_REG_3__SCAN_IN | ~n36154;
  assign n33935 = ~P3_EBX_REG_3__SCAN_IN | ~n35935;
  assign n33937 = ~n33936 | ~n33935;
  assign n33939 = ~n33938 & ~n33937;
  assign n33941 = ~n33940 | ~n33939;
  assign n33950 = ~n33942 & ~n33941;
  assign n33943 = ~n33944 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n35926 = ~n33943 & ~n34979;
  assign n33946 = ~n33945 | ~n33944;
  assign n36670 = ~n33947 | ~n33946;
  assign n33948 = ~n35926 ^ n36670;
  assign n33949 = ~n35930 | ~n33948;
  assign P3_U2668 = ~n33950 | ~n33949;
  assign n33952 = ~n33970 & ~P3_REIP_REG_19__SCAN_IN;
  assign n33957 = ~n33952 | ~n33951;
  assign n33955 = ~n33953 & ~n35642;
  assign n33954 = ~P3_EBX_REG_19__SCAN_IN | ~n34986;
  assign n33956 = ~n33955 | ~n33954;
  assign n33969 = ~n33957 | ~n33956;
  assign n33959 = ~P3_PHYADDRPOINTER_REG_19__SCAN_IN | ~n36154;
  assign n33958 = ~P3_EBX_REG_19__SCAN_IN | ~n35935;
  assign n33960 = ~n33959 | ~n33958;
  assign n33967 = ~n34990 & ~n33960;
  assign n33961 = ~P3_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n34976 = ~n37016 & ~n36220;
  assign n34978 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN | ~n34976;
  assign n33962 = ~n33961 | ~n34978;
  assign n38037 = ~n37578 | ~n33962;
  assign n33963 = ~n34978 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n33964 = ~n33963 & ~n34979;
  assign n33965 = ~n38037 ^ n33964;
  assign n33966 = ~n33965 | ~n35930;
  assign n33968 = ~n33967 | ~n33966;
  assign n33973 = ~n33969 & ~n33968;
  assign n33971 = ~n33970 & ~n34536;
  assign n34999 = ~n33971 & ~n35951;
  assign n33972 = ~P3_REIP_REG_19__SCAN_IN | ~n34999;
  assign P3_U2652 = ~n33973 | ~n33972;
  assign n40055 = ~BUF2_REG_22__SCAN_IN;
  assign n34007 = ~n36239 & ~n40055;
  assign n33975 = ~n22903 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n33974 = ~n22920 | ~P3_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n33979 = ~n33975 | ~n33974;
  assign n33977 = ~n36317 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n33976 = ~n36311 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n33978 = ~n33977 | ~n33976;
  assign n33983 = n33979 | n33978;
  assign n33981 = ~n36298 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n33980 = ~n22910 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n33982 = ~n33981 | ~n33980;
  assign n34003 = ~n33983 & ~n33982;
  assign n33985 = ~n22902 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n33984 = ~n36307 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n33989 = ~n33985 | ~n33984;
  assign n33987 = ~n22917 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n33986 = ~n35392 | ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n33988 = ~n33987 | ~n33986;
  assign n33997 = ~n33989 & ~n33988;
  assign n33991 = ~n22919 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n33990 = ~n22914 | ~P3_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n33995 = ~n33991 | ~n33990;
  assign n33993 = ~n22913 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n33992 = ~n36320 | ~P3_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n33994 = ~n33993 | ~n33992;
  assign n33996 = ~n33995 & ~n33994;
  assign n34001 = ~n33997 | ~n33996;
  assign n33999 = ~n36294 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n33998 = ~n22923 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n34000 = ~n33999 | ~n33998;
  assign n34002 = ~n34001 & ~n34000;
  assign n39500 = ~n34003 | ~n34002;
  assign n34005 = ~n36333 | ~n39500;
  assign n34004 = ~BUF2_REG_6__SCAN_IN | ~n36338;
  assign n34006 = ~n34005 | ~n34004;
  assign n34010 = ~n34007 & ~n34006;
  assign n34008 = ~n34011 ^ P3_EAX_REG_22__SCAN_IN;
  assign n34009 = ~n34008 | ~n36243;
  assign P3_U2713 = ~n34010 | ~n34009;
  assign n34015 = ~n34011;
  assign n34012 = ~n43967 & ~n34968;
  assign n34014 = ~n34013 & ~n34012;
  assign n34019 = ~n34015 & ~n34014;
  assign n34017 = ~n36282 | ~BUF2_REG_21__SCAN_IN;
  assign n34016 = ~n36338 | ~BUF2_REG_5__SCAN_IN;
  assign n34018 = ~n34017 | ~n34016;
  assign n34052 = ~n34019 & ~n34018;
  assign n34021 = ~n22902 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n34020 = ~n22914 | ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n34025 = ~n34021 | ~n34020;
  assign n34023 = ~n22913 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n34022 = ~n36320 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n34024 = ~n34023 | ~n34022;
  assign n34050 = ~n34025 & ~n34024;
  assign n34027 = ~n22919 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n34026 = ~n22903 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n34031 = ~n34027 | ~n34026;
  assign n34029 = ~n36310 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n34028 = ~n22917 | ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n34030 = ~n34029 | ~n34028;
  assign n34039 = ~n34031 & ~n34030;
  assign n34033 = ~n36317 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n34032 = ~n36307 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n34037 = ~n34033 | ~n34032;
  assign n34035 = ~n35392 | ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n34034 = ~n36311 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n34036 = ~n34035 | ~n34034;
  assign n34038 = ~n34037 & ~n34036;
  assign n34048 = ~n34039 | ~n34038;
  assign n34041 = n22901 | n34767;
  assign n34040 = ~n22923 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n34044 = ~n34041 | ~n34040;
  assign n34772 = ~P3_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n34043 = ~n34042 & ~n34772;
  assign n34046 = ~n34044 & ~n34043;
  assign n34045 = ~n36294 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n34047 = ~n34046 | ~n34045;
  assign n34049 = ~n34048 & ~n34047;
  assign n37918 = ~n34050 | ~n34049;
  assign n34051 = ~n36333 | ~n37918;
  assign P3_U2714 = ~n34052 | ~n34051;
  assign n34278 = ~n43033 & ~n35875;
  assign n34054 = ~n34278;
  assign n34053 = ~n43709 | ~P1_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n34062 = ~n34054 | ~n34053;
  assign n34056 = ~n34057;
  assign n34282 = n35323 ^ n35322;
  assign n34060 = ~n43707 | ~n34282;
  assign n34059 = ~n43362 | ~n35889;
  assign n34061 = ~n34060 | ~n34059;
  assign n34065 = ~n34062 & ~n34061;
  assign n35884 = ~n34063;
  assign n34064 = ~n35884 | ~n43367;
  assign P1_U2996 = ~n34065 | ~n34064;
  assign n34067 = ~n34898 & ~n34136;
  assign n34066 = ~n39934 & ~n35517;
  assign n34069 = ~n34067 & ~n34066;
  assign n34068 = ~P1_EAX_REG_4__SCAN_IN | ~n43732;
  assign P1_U2900 = ~n34069 | ~n34068;
  assign n34072 = ~n34241 & ~n39892;
  assign n34111 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~n37475;
  assign n38050 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n34111;
  assign n34073 = ~n38050 & ~n39937;
  assign n34079 = ~n34072 | ~n34073;
  assign n34077 = ~n43722 & ~n38050;
  assign n35475 = ~n34552;
  assign n34717 = ~n35475 & ~n35165;
  assign n34075 = ~n39302 & ~n34682;
  assign n34089 = ~n34075 & ~n34073;
  assign n34076 = ~n34089 & ~n39946;
  assign n34596 = n34077 | n34076;
  assign n34078 = ~n40017 | ~n34596;
  assign n34087 = ~n34079 | ~n34078;
  assign n34249 = ~n39901 & ~n43729;
  assign n34081 = ~n34249 | ~DATAI_31_;
  assign n34248 = ~n39896 & ~n43729;
  assign n34080 = ~n34248 | ~BUF1_REG_31__SCAN_IN;
  assign n34125 = ~n34270 | ~n34679;
  assign n34736 = ~n34560 | ~n34119;
  assign n38132 = ~n34125 & ~n34736;
  assign n34085 = ~n40014 | ~n38132;
  assign n34083 = ~n34248 | ~BUF1_REG_23__SCAN_IN;
  assign n34082 = ~n34249 | ~DATAI_23_;
  assign n34731 = ~n34560 | ~n34551;
  assign n39888 = ~n34125 & ~n34731;
  assign n34084 = ~n40022 | ~n39888;
  assign n34086 = ~n34085 | ~n34084;
  assign n34096 = ~n34087 & ~n34086;
  assign n34092 = ~n39946 & ~n34090;
  assign n34091 = ~n39307 & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n35185 = ~n37486 & ~n34091;
  assign n34093 = ~n38050 | ~n39946;
  assign n34095 = ~P1_INSTQUEUE_REG_11__7__SCAN_IN | ~n34599;
  assign P1_U3128 = ~n34096 | ~n34095;
  assign n34098 = ~n34241 & ~n34097;
  assign n34100 = ~n34098 | ~n34073;
  assign n34099 = ~n40043 | ~n34596;
  assign n34108 = ~n34100 | ~n34099;
  assign n34102 = ~n34248 | ~BUF1_REG_29__SCAN_IN;
  assign n34101 = ~n34249 | ~DATAI_29_;
  assign n34106 = ~n40038 | ~n38132;
  assign n34104 = ~n34249 | ~DATAI_21_;
  assign n34103 = ~n34248 | ~BUF1_REG_21__SCAN_IN;
  assign n34105 = ~n40049 | ~n39888;
  assign n34107 = ~n34106 | ~n34105;
  assign n34110 = ~n34108 & ~n34107;
  assign n34109 = ~P1_INSTQUEUE_REG_11__5__SCAN_IN | ~n34599;
  assign P1_U3126 = ~n34110 | ~n34109;
  assign n39298 = ~n34111 | ~n34677;
  assign n34112 = ~n39298 & ~n39937;
  assign n34118 = ~n34072 | ~n34112;
  assign n34116 = ~n43722 & ~n39298;
  assign n34113 = ~n35165;
  assign n34114 = ~n39302 & ~n34113;
  assign n34126 = ~n34114 & ~n34112;
  assign n34115 = ~n34126 & ~n39946;
  assign n34360 = n34116 | n34115;
  assign n34117 = ~n40017 | ~n34360;
  assign n34123 = ~n34118 | ~n34117;
  assign n38123 = ~n34125 & ~n35173;
  assign n34121 = ~n40022 | ~n38123;
  assign n39383 = ~n34125 & ~n35172;
  assign n34120 = ~n40014 | ~n39383;
  assign n34122 = ~n34121 | ~n34120;
  assign n34133 = ~n34123 & ~n34122;
  assign n34128 = ~n34125 & ~n35178;
  assign n34127 = ~n34126;
  assign n34129 = ~n34128 & ~n34127;
  assign n34130 = ~n39298 | ~n39946;
  assign n34132 = ~P1_INSTQUEUE_REG_9__7__SCAN_IN | ~n34363;
  assign P1_U3112 = ~n34133 | ~n34132;
  assign n34135 = ~n34241 & ~n34134;
  assign n34138 = ~n34135 | ~n34073;
  assign n34137 = ~n39984 | ~n34596;
  assign n34146 = ~n34138 | ~n34137;
  assign n34140 = ~n34249 | ~DATAI_28_;
  assign n34139 = ~n34248 | ~BUF1_REG_28__SCAN_IN;
  assign n34144 = ~n39981 | ~n38132;
  assign n34142 = ~n34249 | ~DATAI_20_;
  assign n34141 = ~n34248 | ~BUF1_REG_20__SCAN_IN;
  assign n34143 = ~n39989 | ~n39888;
  assign n34145 = ~n34144 | ~n34143;
  assign n34148 = ~n34146 & ~n34145;
  assign n34147 = ~P1_INSTQUEUE_REG_11__4__SCAN_IN | ~n34599;
  assign P1_U3125 = ~n34148 | ~n34147;
  assign n34150 = ~n34241 & ~n34149;
  assign n34153 = ~n34150 | ~n34112;
  assign n34152 = ~n40028 | ~n34360;
  assign n34161 = ~n34153 | ~n34152;
  assign n34155 = ~n34248 | ~BUF1_REG_22__SCAN_IN;
  assign n34154 = ~n34249 | ~DATAI_22_;
  assign n34159 = ~n40033 | ~n38123;
  assign n34157 = ~n34249 | ~DATAI_30_;
  assign n34156 = ~n34248 | ~BUF1_REG_30__SCAN_IN;
  assign n34158 = ~n40025 | ~n39383;
  assign n34160 = ~n34159 | ~n34158;
  assign n34163 = ~n34161 & ~n34160;
  assign n34162 = ~P1_INSTQUEUE_REG_9__6__SCAN_IN | ~n34363;
  assign P1_U3111 = ~n34163 | ~n34162;
  assign n34168 = ~n34165 | ~n34073;
  assign n34167 = ~n39995 | ~n34596;
  assign n34176 = ~n34168 | ~n34167;
  assign n34170 = ~n34249 | ~DATAI_27_;
  assign n34169 = ~n34248 | ~BUF1_REG_27__SCAN_IN;
  assign n34174 = ~n39992 | ~n38132;
  assign n34172 = ~n34248 | ~BUF1_REG_19__SCAN_IN;
  assign n34171 = ~n34249 | ~DATAI_19_;
  assign n34173 = ~n40000 | ~n39888;
  assign n34175 = ~n34174 | ~n34173;
  assign n34178 = ~n34176 & ~n34175;
  assign n34177 = ~P1_INSTQUEUE_REG_11__3__SCAN_IN | ~n34599;
  assign P1_U3124 = ~n34178 | ~n34177;
  assign n34180 = ~n34165 | ~n34112;
  assign n34179 = ~n39995 | ~n34360;
  assign n34184 = ~n34180 | ~n34179;
  assign n34182 = ~n40000 | ~n38123;
  assign n34181 = ~n39992 | ~n39383;
  assign n34183 = ~n34182 | ~n34181;
  assign n34186 = ~n34184 & ~n34183;
  assign n34185 = ~P1_INSTQUEUE_REG_9__3__SCAN_IN | ~n34363;
  assign P1_U3108 = ~n34186 | ~n34185;
  assign n34191 = ~n34188 | ~n34112;
  assign n34190 = ~n39973 | ~n34360;
  assign n34199 = ~n34191 | ~n34190;
  assign n34193 = ~n34249 | ~DATAI_17_;
  assign n34192 = ~n34248 | ~BUF1_REG_17__SCAN_IN;
  assign n34197 = ~n39978 | ~n38123;
  assign n34195 = ~n34248 | ~BUF1_REG_25__SCAN_IN;
  assign n34194 = ~n34249 | ~DATAI_25_;
  assign n34196 = ~n39970 | ~n39383;
  assign n34198 = ~n34197 | ~n34196;
  assign n34201 = ~n34199 & ~n34198;
  assign n34200 = ~P1_INSTQUEUE_REG_9__1__SCAN_IN | ~n34363;
  assign P1_U3106 = ~n34201 | ~n34200;
  assign n34203 = ~n34135 | ~n34112;
  assign n34202 = ~n39984 | ~n34360;
  assign n34207 = ~n34203 | ~n34202;
  assign n34205 = ~n39989 | ~n38123;
  assign n34204 = ~n39981 | ~n39383;
  assign n34206 = ~n34205 | ~n34204;
  assign n34209 = ~n34207 & ~n34206;
  assign n34208 = ~P1_INSTQUEUE_REG_9__4__SCAN_IN | ~n34363;
  assign P1_U3109 = ~n34209 | ~n34208;
  assign n34211 = ~n34098 | ~n34112;
  assign n34210 = ~n40043 | ~n34360;
  assign n34215 = ~n34211 | ~n34210;
  assign n34213 = ~n40049 | ~n38123;
  assign n34212 = ~n40038 | ~n39383;
  assign n34214 = ~n34213 | ~n34212;
  assign n34217 = ~n34215 & ~n34214;
  assign n34216 = ~P1_INSTQUEUE_REG_9__5__SCAN_IN | ~n34363;
  assign P1_U3110 = ~n34217 | ~n34216;
  assign n34219 = ~n34188 | ~n34073;
  assign n34218 = ~n39973 | ~n34596;
  assign n34223 = ~n34219 | ~n34218;
  assign n34221 = ~n39970 | ~n38132;
  assign n34220 = ~n39978 | ~n39888;
  assign n34222 = ~n34221 | ~n34220;
  assign n34225 = ~n34223 & ~n34222;
  assign n34224 = ~P1_INSTQUEUE_REG_11__1__SCAN_IN | ~n34599;
  assign P1_U3122 = ~n34225 | ~n34224;
  assign n34227 = ~n34241 & ~n34226;
  assign n34230 = ~n34227 | ~n34112;
  assign n34229 = ~n40006 | ~n34360;
  assign n34238 = ~n34230 | ~n34229;
  assign n34232 = ~n34249 | ~DATAI_18_;
  assign n34231 = ~n34248 | ~BUF1_REG_18__SCAN_IN;
  assign n34236 = ~n40011 | ~n38123;
  assign n34234 = ~n34248 | ~BUF1_REG_26__SCAN_IN;
  assign n34233 = ~n34249 | ~DATAI_26_;
  assign n34235 = ~n40003 | ~n39383;
  assign n34237 = ~n34236 | ~n34235;
  assign n34240 = ~n34238 & ~n34237;
  assign n34239 = ~P1_INSTQUEUE_REG_9__2__SCAN_IN | ~n34363;
  assign P1_U3107 = ~n34240 | ~n34239;
  assign n34245 = ~n34242 | ~n34073;
  assign n34244 = ~n39962 | ~n34596;
  assign n34255 = ~n34245 | ~n34244;
  assign n34247 = ~n34249 | ~DATAI_24_;
  assign n34246 = ~n34248 | ~BUF1_REG_24__SCAN_IN;
  assign n34253 = ~n39939 | ~n38132;
  assign n34251 = ~n34248 | ~BUF1_REG_16__SCAN_IN;
  assign n34250 = ~n34249 | ~DATAI_16_;
  assign n34252 = ~n39967 | ~n39888;
  assign n34254 = ~n34253 | ~n34252;
  assign n34257 = ~n34255 & ~n34254;
  assign n34256 = ~P1_INSTQUEUE_REG_11__0__SCAN_IN | ~n34599;
  assign P1_U3121 = ~n34257 | ~n34256;
  assign n35021 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n37474 = n34677 | n35021;
  assign n35010 = ~n37474 & ~n39937;
  assign n34263 = ~n34150 | ~n35010;
  assign n34261 = ~n43722 & ~n37474;
  assign n34409 = ~n34258;
  assign n34259 = ~n37476 & ~n34682;
  assign n34264 = ~n34259 & ~n35010;
  assign n34260 = ~n34264 & ~n39946;
  assign n35011 = n34261 | n34260;
  assign n34262 = ~n40028 | ~n35011;
  assign n34274 = ~n34263 | ~n34262;
  assign n34266 = ~n22916 & ~n34725;
  assign n34265 = ~n34264 | ~n39315;
  assign n34267 = ~n34266 & ~n34265;
  assign n34268 = ~n37474 | ~n39946;
  assign n34272 = ~P1_INSTQUEUE_REG_15__6__SCAN_IN | ~n35014;
  assign n35032 = ~n34270 | ~n34576;
  assign n40037 = ~n35032 & ~n34731;
  assign n34271 = ~n40033 | ~n40037;
  assign n34273 = ~n34272 | ~n34271;
  assign n34276 = ~n34274 & ~n34273;
  assign n38889 = ~n35032 & ~n34736;
  assign n34275 = ~n40025 | ~n38889;
  assign P1_U3159 = ~n34276 | ~n34275;
  assign n34277 = ~n43441 & ~n35869;
  assign n34297 = ~n34278 & ~n34277;
  assign n34281 = ~n34283 & ~n34279;
  assign n34280 = ~n41976 & ~n34290;
  assign n35364 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN & ~n35361;
  assign n34294 = ~n36906 | ~n34282;
  assign n34284 = ~n42922 & ~n34283;
  assign n34289 = ~n34285 & ~n34284;
  assign n34288 = ~n34287 & ~n34286;
  assign n34292 = ~n34289 & ~n34288;
  assign n34291 = ~n36891 | ~n34290;
  assign n35365 = ~n34292 | ~n34291;
  assign n34293 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN | ~n35365;
  assign n34295 = ~n34294 | ~n34293;
  assign n34296 = ~n35364 & ~n34295;
  assign P1_U3028 = ~n34297 | ~n34296;
  assign n34333 = BUF2_REG_27__SCAN_IN & n36282;
  assign n34299 = ~n36317 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n34298 = ~n36307 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n34303 = ~n34299 | ~n34298;
  assign n34301 = ~n22914 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n34300 = ~n22923 | ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n34302 = ~n34301 | ~n34300;
  assign n34311 = ~n34303 & ~n34302;
  assign n34305 = ~n22903 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n34304 = ~n36320 | ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n34309 = ~n34305 | ~n34304;
  assign n34307 = ~n36310 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n34306 = ~n22917 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n34308 = ~n34307 | ~n34306;
  assign n34310 = ~n34309 & ~n34308;
  assign n34327 = ~n34311 | ~n34310;
  assign n34313 = ~n22919 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n34312 = ~n36311 | ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n34317 = ~n34313 | ~n34312;
  assign n34315 = ~n22902 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n34314 = ~n36298 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n34316 = ~n34315 | ~n34314;
  assign n34325 = ~n34317 & ~n34316;
  assign n34319 = ~n22913 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n34318 = ~n22920 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n34323 = ~n34319 | ~n34318;
  assign n34321 = ~n36294 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n34320 = ~n35392 | ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n34322 = ~n34321 | ~n34320;
  assign n34324 = ~n34323 & ~n34322;
  assign n34326 = ~n34325 | ~n34324;
  assign n34764 = ~n34327 & ~n34326;
  assign n34763 = ~n34329 | ~n34328;
  assign n41388 = n34764 ^ n34763;
  assign n34331 = ~n36333 | ~n41388;
  assign n34330 = ~n36338 | ~BUF2_REG_11__SCAN_IN;
  assign n34332 = ~n34331 | ~n34330;
  assign n34338 = ~n34333 & ~n34332;
  assign n34334 = ~P3_EAX_REG_27__SCAN_IN | ~n36243;
  assign n34336 = ~n34334 | ~n34335;
  assign n34806 = ~n34808;
  assign n34337 = ~n34336 | ~n34806;
  assign P3_U2708 = ~n34338 | ~n34337;
  assign n34342 = ~n34818;
  assign n34341 = ~n34340 | ~n34339;
  assign n36119 = ~n34342 | ~n34341;
  assign n34347 = ~n36119 & ~n43298;
  assign n34345 = n34344 | n34343;
  assign n34346 = ~n36109 & ~n44019;
  assign n34349 = ~n34347 & ~n34346;
  assign n34348 = ~P1_EBX_REG_5__SCAN_IN | ~n44023;
  assign P1_U2867 = ~n34349 | ~n34348;
  assign n34353 = ~n35459 & ~n34350;
  assign n34352 = ~n34351 & ~n34843;
  assign n34359 = ~n34353 & ~n34352;
  assign n34354 = ~P3_EAX_REG_11__SCAN_IN | ~n36243;
  assign n34357 = ~n34354 | ~n34355;
  assign n34849 = ~n34356 & ~n34355;
  assign n34847 = ~n34849;
  assign n34358 = ~n34357 | ~n34847;
  assign P3_U2724 = ~n34359 | ~n34358;
  assign n34362 = ~n34242 | ~n34112;
  assign n34361 = ~n39962 | ~n34360;
  assign n34367 = ~n34362 | ~n34361;
  assign n34365 = ~P1_INSTQUEUE_REG_9__0__SCAN_IN | ~n34363;
  assign n34364 = ~n39967 | ~n38123;
  assign n34366 = ~n34365 | ~n34364;
  assign n34369 = ~n34367 & ~n34366;
  assign n34368 = ~n39939 | ~n39383;
  assign P1_U3105 = ~n34369 | ~n34368;
  assign n34371 = ~n22903 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n34370 = ~n36317 | ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n34375 = ~n34371 | ~n34370;
  assign n34373 = ~n22919 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n34372 = ~n36307 | ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n34374 = ~n34373 | ~n34372;
  assign n34379 = n34375 | n34374;
  assign n34377 = ~n22917 | ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n34376 = ~n35392 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n34378 = ~n34377 | ~n34376;
  assign n34399 = ~n34379 & ~n34378;
  assign n34381 = ~n22902 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n34380 = ~n22920 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n34385 = ~n34381 | ~n34380;
  assign n34383 = ~n36298 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n34382 = ~n36320 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n34384 = ~n34383 | ~n34382;
  assign n34393 = ~n34385 & ~n34384;
  assign n34387 = ~n36310 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n34386 = ~n22914 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n34391 = ~n34387 | ~n34386;
  assign n34389 = ~n36294 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n34388 = ~n22923 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n34390 = ~n34389 | ~n34388;
  assign n34392 = ~n34391 & ~n34390;
  assign n34397 = ~n34393 | ~n34392;
  assign n34395 = ~n22913 | ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n34394 = ~n36311 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n34396 = ~n34395 | ~n34394;
  assign n34398 = ~n34397 & ~n34396;
  assign n35308 = ~n34399 | ~n34398;
  assign n34407 = ~n42135 | ~n35308;
  assign n34403 = ~P3_EBX_REG_15__SCAN_IN | ~n43930;
  assign n34405 = ~n34403 | ~n34402;
  assign n34406 = ~n34405 | ~n35421;
  assign P3_U2688 = ~n34407 | ~n34406;
  assign n34408 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n38397 = ~n34408 | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n34749 = ~n38397 & ~n39937;
  assign n34415 = ~n34072 | ~n34749;
  assign n34420 = ~n38397;
  assign n34413 = ~n34420 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n34411 = ~n38482 | ~n35165;
  assign n34410 = ~n34749;
  assign n34412 = ~n39315 | ~n34421;
  assign n34414 = ~n40017 | ~n34748;
  assign n34419 = ~n34415 | ~n34414;
  assign n34737 = ~n22916 | ~n34576;
  assign n38469 = ~n34737 & ~n35172;
  assign n34417 = ~n40014 | ~n38469;
  assign n38557 = ~n34737 & ~n35173;
  assign n34416 = ~n40022 | ~n38557;
  assign n34418 = ~n34417 | ~n34416;
  assign n34427 = ~n34419 & ~n34418;
  assign n34424 = ~n34420 & ~n39315;
  assign n34422 = ~n34737 & ~n35178;
  assign n34423 = ~n34422 & ~n34421;
  assign n34426 = ~P1_INSTQUEUE_REG_5__7__SCAN_IN | ~n34752;
  assign P1_U3080 = ~n34427 | ~n34426;
  assign n34429 = ~n34098 | ~n34749;
  assign n34428 = ~n40043 | ~n34748;
  assign n34433 = ~n34429 | ~n34428;
  assign n34431 = ~n40038 | ~n38469;
  assign n34430 = ~n40049 | ~n38557;
  assign n34432 = ~n34431 | ~n34430;
  assign n34435 = ~n34433 & ~n34432;
  assign n34434 = ~P1_INSTQUEUE_REG_5__5__SCAN_IN | ~n34752;
  assign P1_U3078 = ~n34435 | ~n34434;
  assign n34437 = ~n34150 | ~n34749;
  assign n34436 = ~n40028 | ~n34748;
  assign n34441 = ~n34437 | ~n34436;
  assign n34439 = ~n40025 | ~n38469;
  assign n34438 = ~n40033 | ~n38557;
  assign n34440 = ~n34439 | ~n34438;
  assign n34443 = ~n34441 & ~n34440;
  assign n34442 = ~P1_INSTQUEUE_REG_5__6__SCAN_IN | ~n34752;
  assign P1_U3079 = ~n34443 | ~n34442;
  assign n34445 = ~n34165 | ~n34749;
  assign n34444 = ~n39995 | ~n34748;
  assign n34449 = ~n34445 | ~n34444;
  assign n34447 = ~n39992 | ~n38469;
  assign n34446 = ~n40000 | ~n38557;
  assign n34448 = ~n34447 | ~n34446;
  assign n34451 = ~n34449 & ~n34448;
  assign n34450 = ~P1_INSTQUEUE_REG_5__3__SCAN_IN | ~n34752;
  assign P1_U3076 = ~n34451 | ~n34450;
  assign n34453 = ~n34227 | ~n34749;
  assign n34452 = ~n40006 | ~n34748;
  assign n34457 = ~n34453 | ~n34452;
  assign n34455 = ~n40003 | ~n38469;
  assign n34454 = ~n40011 | ~n38557;
  assign n34456 = ~n34455 | ~n34454;
  assign n34459 = ~n34457 & ~n34456;
  assign n34458 = ~P1_INSTQUEUE_REG_5__2__SCAN_IN | ~n34752;
  assign P1_U3075 = ~n34459 | ~n34458;
  assign n34461 = ~n34188 | ~n34749;
  assign n34460 = ~n39973 | ~n34748;
  assign n34465 = ~n34461 | ~n34460;
  assign n34463 = ~n39970 | ~n38469;
  assign n34462 = ~n39978 | ~n38557;
  assign n34464 = ~n34463 | ~n34462;
  assign n34467 = ~n34465 & ~n34464;
  assign n34466 = ~P1_INSTQUEUE_REG_5__1__SCAN_IN | ~n34752;
  assign P1_U3074 = ~n34467 | ~n34466;
  assign n34469 = ~n34135 | ~n34749;
  assign n34468 = ~n39984 | ~n34748;
  assign n34473 = ~n34469 | ~n34468;
  assign n34471 = ~n39981 | ~n38469;
  assign n34470 = ~n39989 | ~n38557;
  assign n34472 = ~n34471 | ~n34470;
  assign n34475 = ~n34473 & ~n34472;
  assign n34474 = ~P1_INSTQUEUE_REG_5__4__SCAN_IN | ~n34752;
  assign P1_U3077 = ~n34475 | ~n34474;
  assign n34494 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n34489;
  assign n34483 = n34478 | n34476;
  assign n34481 = ~n34477 | ~n34495;
  assign n34479 = n34478 | n39937;
  assign n34480 = ~n34479 | ~n34677;
  assign n34482 = ~n34481 | ~n34480;
  assign n34484 = ~n34483 | ~n34482;
  assign n34488 = n34484 & P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n34486 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~n34484;
  assign n34487 = ~n34486 & ~n34485;
  assign n34491 = ~n34488 & ~n34487;
  assign n34490 = ~n34489 & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n34492 = ~n34491 & ~n34490;
  assign n34493 = ~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & ~n34492;
  assign n34506 = ~n34495 & ~n24830;
  assign n34497 = ~P1_FLUSH_REG_SCAN_IN & ~P1_MORE_REG_SCAN_IN;
  assign n34501 = ~n34497 & ~n34496;
  assign n34500 = n34499 | n34498;
  assign n34504 = ~n34501 & ~n34500;
  assign n34503 = ~n34502;
  assign n34510 = ~n35500 & ~n34509;
  assign n34516 = ~n34515 | ~n34514;
  assign n34519 = ~n34517 & ~n34516;
  assign n34520 = ~n34519 & ~n34518;
  assign n35622 = ~n34523;
  assign P1_U3466 = ~n34524 | ~n35622;
  assign n34525 = ~P3_PHYADDRPOINTER_REG_17__SCAN_IN & ~n34526;
  assign n36872 = ~n34525 & ~n34976;
  assign n34527 = ~n34526 | ~n35924;
  assign n34528 = ~n41401 | ~n34527;
  assign n34529 = n36872 ^ n34528;
  assign n34544 = ~n34529 & ~n35942;
  assign n36874 = ~P3_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n34530 = ~n36874 & ~n35947;
  assign n34542 = ~n34990 & ~n34530;
  assign n34533 = ~n34531 | ~P3_EBX_REG_17__SCAN_IN;
  assign n34532 = ~n34985 & ~n35642;
  assign n34535 = ~n34533 | ~n34532;
  assign n34534 = ~n35935 | ~P3_EBX_REG_17__SCAN_IN;
  assign n34540 = ~n34535 | ~n34534;
  assign n34538 = ~n34546 & ~n34536;
  assign n34537 = ~P3_REIP_REG_17__SCAN_IN | ~n35525;
  assign n34539 = ~n34538 & ~n34537;
  assign n34541 = ~n34540 & ~n34539;
  assign n34543 = ~n34542 | ~n34541;
  assign n34549 = ~n34544 & ~n34543;
  assign n34983 = ~n34546 & ~n34545;
  assign n34548 = ~n34983 | ~n34547;
  assign P3_U2654 = ~n34549 | ~n34548;
  assign n34556 = ~n35623 & ~n34550;
  assign n34554 = ~n34551 | ~n39315;
  assign n34579 = ~P1_STATE2_REG_1__SCAN_IN | ~n39307;
  assign n34553 = ~n34552 | ~n34579;
  assign n34555 = ~n34554 | ~n34553;
  assign n34557 = n34556 | n34555;
  assign n34559 = ~n34584 | ~n34557;
  assign n34558 = ~n34585 | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign P1_U3478 = ~n34559 | ~n34558;
  assign n34561 = ~n34560 | ~n39944;
  assign n34562 = ~n35178 | ~n34561;
  assign n34564 = ~n34562 | ~n39315;
  assign n34563 = ~n39301 | ~n34579;
  assign n34565 = ~n34564 | ~n34563;
  assign n34567 = ~n34584 | ~n34565;
  assign n34566 = ~n34585 | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign P1_U3477 = ~n34567 | ~n34566;
  assign n34568 = n22916 ^ n34725;
  assign n34571 = ~n34568 | ~n39315;
  assign n34570 = ~n34569 | ~n34579;
  assign n34572 = ~n34571 | ~n34570;
  assign n34574 = ~n34584 | ~n34572;
  assign n34573 = ~n34585 | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign P1_U3475 = ~n34574 | ~n34573;
  assign n34577 = ~n34576 & ~n34575;
  assign n34578 = ~n34577 & ~n39946;
  assign n34582 = ~n34578 | ~n34725;
  assign n34581 = ~n34580 | ~n34579;
  assign n34583 = ~n34582 | ~n34581;
  assign n34587 = ~n34584 | ~n34583;
  assign n34586 = ~n34585 | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign P1_U3476 = ~n34587 | ~n34586;
  assign n34589 = ~n34227 | ~n34073;
  assign n34588 = ~n40006 | ~n34596;
  assign n34593 = ~n34589 | ~n34588;
  assign n34591 = ~P1_INSTQUEUE_REG_11__2__SCAN_IN | ~n34599;
  assign n34590 = ~n40011 | ~n39888;
  assign n34592 = ~n34591 | ~n34590;
  assign n34595 = ~n34593 & ~n34592;
  assign n34594 = ~n40003 | ~n38132;
  assign P1_U3123 = ~n34595 | ~n34594;
  assign n34598 = ~n34150 | ~n34073;
  assign n34597 = ~n40028 | ~n34596;
  assign n34603 = ~n34598 | ~n34597;
  assign n34601 = ~P1_INSTQUEUE_REG_11__6__SCAN_IN | ~n34599;
  assign n34600 = ~n40025 | ~n38132;
  assign n34602 = ~n34601 | ~n34600;
  assign n34605 = ~n34603 & ~n34602;
  assign n34604 = ~n40033 | ~n39888;
  assign P1_U3127 = ~n34605 | ~n34604;
  assign n34608 = ~n34898 & ~n34606;
  assign n34607 = ~n39934 & ~n36109;
  assign n34610 = ~n34608 & ~n34607;
  assign n34609 = ~P1_EAX_REG_5__SCAN_IN | ~n43732;
  assign P1_U2899 = ~n34610 | ~n34609;
  assign n34613 = ~n36153 & ~n34611;
  assign n34612 = ~P3_EBX_REG_0__SCAN_IN;
  assign n34619 = ~n34613 & ~n34612;
  assign n34614 = ~n34626 & ~n35924;
  assign n34617 = ~n34614 | ~n35670;
  assign n35907 = ~n34615;
  assign n34616 = ~n35608 | ~n35907;
  assign n34618 = ~n34617 | ~n34616;
  assign n34621 = ~n34619 & ~n34618;
  assign n34620 = ~P3_REIP_REG_0__SCAN_IN | ~n35525;
  assign P3_U2671 = ~n34621 | ~n34620;
  assign n34623 = ~P3_PHYADDRPOINTER_REG_27__SCAN_IN | ~n36154;
  assign n34622 = ~P3_EBX_REG_27__SCAN_IN | ~n35935;
  assign n34636 = ~n34623 | ~n34622;
  assign n34661 = ~P3_REIP_REG_25__SCAN_IN | ~n34624;
  assign n34628 = ~n40723 & ~n34661;
  assign n34630 = ~P3_REIP_REG_27__SCAN_IN & ~n35541;
  assign n34627 = ~n34626 & ~n34625;
  assign n35523 = ~n34628 | ~n34627;
  assign n34664 = ~n35525 | ~n35523;
  assign n34629 = ~n35542 & ~n34664;
  assign n34634 = ~n34630 & ~n34629;
  assign n34632 = ~n35527 & ~n35642;
  assign n34631 = ~P3_EBX_REG_27__SCAN_IN | ~n34656;
  assign n34633 = ~n34632 | ~n34631;
  assign n34635 = ~n34634 | ~n34633;
  assign n34644 = ~n34636 & ~n34635;
  assign n41158 = ~P3_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n40725 = ~P3_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n34639 = ~n40725 | ~n40733;
  assign n40724 = ~n35529 | ~n34639;
  assign n34640 = ~n41156 & ~n34641;
  assign n34642 = ~n34640 & ~n35942;
  assign n34643 = ~n34642 | ~n35532;
  assign P3_U2644 = ~n34644 | ~n34643;
  assign n34647 = ~n34646 & ~n34645;
  assign n34648 = ~n34647 & ~n33538;
  assign n34650 = ~n34648 | ~n34917;
  assign n34649 = ~n35967 | ~P2_EBX_REG_9__SCAN_IN;
  assign n34654 = n34650 & n34649;
  assign n41707 = n34652 ^ n34651;
  assign n34653 = ~n41707 | ~n43525;
  assign P2_U2878 = ~n34654 | ~n34653;
  assign n34658 = ~n34655 & ~n41389;
  assign n34657 = ~n35944 | ~n34656;
  assign n34670 = ~n34658 & ~n34657;
  assign n34660 = ~n34659 | ~n40723;
  assign n34663 = ~n34661 & ~n34660;
  assign n34662 = ~n40725 & ~n35947;
  assign n34668 = ~n34663 & ~n34662;
  assign n34666 = ~n41389 & ~n35945;
  assign n34665 = ~n40723 & ~n34664;
  assign n34667 = ~n34666 & ~n34665;
  assign n34669 = ~n34668 | ~n34667;
  assign n34676 = ~n34670 & ~n34669;
  assign n34672 = ~n40724 & ~n34671;
  assign n34674 = ~n34672 & ~n35942;
  assign n34675 = ~n34674 | ~n34673;
  assign P3_U2645 = ~n34676 | ~n34675;
  assign n34678 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~n34677;
  assign n39028 = ~n34678 | ~n35163;
  assign n35152 = ~n39028 & ~n39937;
  assign n34681 = ~n34188 | ~n35152;
  assign n35179 = ~n22916 | ~n34679;
  assign n38478 = ~n35179 & ~n34731;
  assign n34680 = ~n39978 | ~n38478;
  assign n34698 = ~n34681 | ~n34680;
  assign n34683 = ~n39030 & ~n34682;
  assign n34692 = ~n34683 & ~n35152;
  assign n34686 = ~n34692;
  assign n34688 = ~n34686 & ~n34691;
  assign n34690 = ~n34688 & ~n34687;
  assign n34689 = ~n39028 | ~n39946;
  assign n34696 = ~P1_INSTQUEUE_REG_3__1__SCAN_IN | ~n35155;
  assign n34694 = ~n43722 & ~n39028;
  assign n34693 = ~n34692 & ~n34691;
  assign n35156 = n34694 | n34693;
  assign n34695 = ~n39973 | ~n35156;
  assign n34697 = ~n34696 | ~n34695;
  assign n34700 = ~n34698 & ~n34697;
  assign n39107 = ~n35179 & ~n34736;
  assign n34699 = ~n39970 | ~n39107;
  assign P1_U3058 = ~n34700 | ~n34699;
  assign n34702 = ~n34227 | ~n35152;
  assign n34701 = ~n40011 | ~n38478;
  assign n34706 = ~n34702 | ~n34701;
  assign n34704 = ~P1_INSTQUEUE_REG_3__2__SCAN_IN | ~n35155;
  assign n34703 = ~n40006 | ~n35156;
  assign n34705 = ~n34704 | ~n34703;
  assign n34708 = ~n34706 & ~n34705;
  assign n34707 = ~n40003 | ~n39107;
  assign P1_U3059 = ~n34708 | ~n34707;
  assign n34710 = ~n34150 | ~n35152;
  assign n34709 = ~n40033 | ~n38478;
  assign n34714 = ~n34710 | ~n34709;
  assign n34712 = ~P1_INSTQUEUE_REG_3__6__SCAN_IN | ~n35155;
  assign n34711 = ~n40028 | ~n35156;
  assign n34713 = ~n34712 | ~n34711;
  assign n34716 = ~n34714 & ~n34713;
  assign n34715 = ~n40025 | ~n39107;
  assign P1_U3063 = ~n34716 | ~n34715;
  assign n35350 = ~n34718;
  assign n34724 = ~n34165 | ~n35350;
  assign n34719 = ~n38482 | ~n34717;
  assign n34720 = ~n34719 | ~n34718;
  assign n34722 = ~n34720 | ~n39315;
  assign n34721 = ~n38481 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n34723 = ~n39995 | ~n35351;
  assign n34735 = ~n34724 | ~n34723;
  assign n34727 = ~n34725 & ~n39946;
  assign n34729 = ~n34727 | ~n22916;
  assign n34728 = ~n38481;
  assign n34733 = ~P1_INSTQUEUE_REG_7__3__SCAN_IN | ~n35354;
  assign n39374 = ~n34737 & ~n34731;
  assign n34732 = ~n40000 | ~n39374;
  assign n34734 = ~n34733 | ~n34732;
  assign n34739 = ~n34735 & ~n34734;
  assign n38562 = ~n34737 & ~n34736;
  assign n34738 = ~n39992 | ~n38562;
  assign P1_U3092 = ~n34739 | ~n34738;
  assign n34741 = ~n34150 | ~n35350;
  assign n34740 = ~n40028 | ~n35351;
  assign n34745 = ~n34741 | ~n34740;
  assign n34743 = ~P1_INSTQUEUE_REG_7__6__SCAN_IN | ~n35354;
  assign n34742 = ~n40033 | ~n39374;
  assign n34744 = ~n34743 | ~n34742;
  assign n34747 = ~n34745 & ~n34744;
  assign n34746 = ~n40025 | ~n38562;
  assign P1_U3095 = ~n34747 | ~n34746;
  assign n34751 = ~n39962 | ~n34748;
  assign n34750 = ~n34242 | ~n34749;
  assign n34756 = ~n34751 | ~n34750;
  assign n34754 = ~P1_INSTQUEUE_REG_5__0__SCAN_IN | ~n34752;
  assign n34753 = ~n39967 | ~n38557;
  assign n34755 = ~n34754 | ~n34753;
  assign n34758 = ~n34756 & ~n34755;
  assign n34757 = ~n39939 | ~n38469;
  assign P1_U3073 = ~n34758 | ~n34757;
  assign n34762 = ~n40325 | ~n43523;
  assign n34760 = ~n35720 | ~n43525;
  assign n34759 = n43525 | P2_EBX_REG_2__SCAN_IN;
  assign n34761 = ~n34760 | ~n34759;
  assign P2_U2885 = ~n34762 | ~n34761;
  assign n34805 = BUF2_REG_28__SCAN_IN & n36282;
  assign n35588 = ~n34764 & ~n34763;
  assign n34765 = ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n34770 = ~n34766 & ~n34765;
  assign n34769 = ~n34768 & ~n34767;
  assign n34777 = ~n34770 & ~n34769;
  assign n34771 = ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n34775 = ~n27301 & ~n34771;
  assign n34774 = ~n34773 & ~n34772;
  assign n34776 = ~n34775 & ~n34774;
  assign n34781 = ~n34777 | ~n34776;
  assign n34779 = ~n22913 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n34778 = ~n22920 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n34780 = ~n34779 | ~n34778;
  assign n34801 = ~n34781 & ~n34780;
  assign n34783 = ~n36294 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n34782 = ~n22919 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n34787 = ~n34783 | ~n34782;
  assign n34785 = ~n36298 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n34784 = ~n36310 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n34786 = ~n34785 | ~n34784;
  assign n34795 = ~n34787 & ~n34786;
  assign n34789 = ~n22903 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n34788 = ~n36317 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n34793 = ~n34789 | ~n34788;
  assign n34791 = ~n22914 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n34790 = ~n36320 | ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n34792 = ~n34791 | ~n34790;
  assign n34794 = ~n34793 & ~n34792;
  assign n34799 = ~n34795 | ~n34794;
  assign n34797 = ~n22917 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n34796 = ~n35392 | ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n34798 = ~n34797 | ~n34796;
  assign n34800 = ~n34799 & ~n34798;
  assign n35587 = ~n34801 | ~n34800;
  assign n41680 = n35588 ^ n35587;
  assign n34803 = ~n36333 | ~n41680;
  assign n34802 = ~n36338 | ~BUF2_REG_12__SCAN_IN;
  assign n34804 = ~n34803 | ~n34802;
  assign n34811 = ~n34805 & ~n34804;
  assign n34807 = ~P3_EAX_REG_28__SCAN_IN | ~n36243;
  assign n34809 = ~n34807 | ~n34806;
  assign n34810 = ~n34809 | ~n35594;
  assign P3_U2707 = ~n34811 | ~n34810;
  assign n34828 = ~n44013 & ~n43794;
  assign n36104 = ~n42185 & ~n35502;
  assign n34816 = ~P1_REIP_REG_5__SCAN_IN | ~n36104;
  assign n34822 = ~n34816 & ~P1_REIP_REG_6__SCAN_IN;
  assign n44014 = n34818 ^ n34817;
  assign n34820 = ~n44014 | ~n43803;
  assign n34819 = ~n43796 | ~P1_EBX_REG_6__SCAN_IN;
  assign n34821 = ~n34820 | ~n34819;
  assign n34826 = ~n34822 & ~n34821;
  assign n34824 = ~n41129 & ~n34823;
  assign n34825 = ~n34824 & ~n43469;
  assign n34827 = ~n34826 | ~n34825;
  assign n34834 = ~n34828 & ~n34827;
  assign n36982 = ~n34829 | ~n41894;
  assign n34832 = ~n34830 & ~n36990;
  assign n34831 = ~n35681 & ~n42175;
  assign n34833 = ~n34832 & ~n34831;
  assign P1_U2834 = ~n34834 | ~n34833;
  assign n34839 = ~n36002 & ~n43634;
  assign n34837 = n34836 & n34835;
  assign n34838 = n42117 & n35381;
  assign n34841 = ~n34839 & ~n34838;
  assign n34840 = ~P2_EAX_REG_13__SCAN_IN | ~n43698;
  assign P2_U2906 = ~n34841 | ~n34840;
  assign n34846 = ~n35459 & ~n34842;
  assign n34845 = ~n34844 & ~n34843;
  assign n34852 = ~n34846 & ~n34845;
  assign n34848 = ~P3_EAX_REG_12__SCAN_IN | ~n36243;
  assign n34850 = ~n34848 | ~n34847;
  assign n35456 = ~P3_EAX_REG_12__SCAN_IN | ~n34849;
  assign n34851 = ~n34850 | ~n35456;
  assign P3_U2723 = ~n34852 | ~n34851;
  assign n34855 = ~n43748 | ~n34853;
  assign n34854 = ~n43767 | ~n40306;
  assign n34873 = ~n34855 | ~n34854;
  assign n34868 = ~n43877 & ~n40311;
  assign n34856 = ~n43159 & ~n35796;
  assign n34857 = ~n43164 & ~n34856;
  assign n34862 = ~n34858 & ~n34857;
  assign n34860 = ~n36600 & ~n34859;
  assign n34861 = ~n34860 & ~n42699;
  assign n34866 = ~n34862 & ~n34861;
  assign n34864 = ~n34863 & ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n34865 = ~n43148 | ~n34864;
  assign n34867 = ~n34866 | ~n34865;
  assign n34871 = ~n34868 & ~n34867;
  assign n34870 = ~n43876 | ~n34869;
  assign n34872 = ~n34871 | ~n34870;
  assign n34875 = ~n34873 & ~n34872;
  assign n34874 = ~P2_REIP_REG_2__SCAN_IN | ~n43880;
  assign P2_U3044 = ~n34875 | ~n34874;
  assign n34878 = ~n43767 | ~n34876;
  assign n34893 = ~n34878 | ~n34877;
  assign n34882 = ~n43893 & ~n34879;
  assign n34881 = ~n43755 & ~n34880;
  assign n34883 = ~n34882 & ~n34881;
  assign n34884 = ~n34883 | ~n42110;
  assign n34891 = ~n34884 | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n34887 = ~n43893 & ~n34885;
  assign n34886 = ~n43755 & ~n37290;
  assign n34888 = ~n34887 & ~n34886;
  assign n34889 = ~n34888 | ~n42600;
  assign n34890 = ~n34889 | ~n33579;
  assign n34892 = ~n34891 | ~n34890;
  assign n34895 = ~n34893 & ~n34892;
  assign n34894 = ~n43583 | ~n37280;
  assign P2_U3046 = ~n34895 | ~n34894;
  assign n34897 = ~n39934 & ~n44013;
  assign n34896 = ~n44063 & ~n43734;
  assign n34900 = ~n34897 & ~n34896;
  assign n34899 = ~n40436 | ~n41773;
  assign P1_U2898 = ~n34900 | ~n34899;
  assign n34905 = ~n37131 & ~n34901;
  assign n36599 = n34903 ^ n34902;
  assign n34904 = ~n36599 & ~n39522;
  assign n34911 = ~n34905 & ~n34904;
  assign n34907 = ~n36744 & ~n36634;
  assign n34908 = ~n34907 | ~n37946;
  assign n34910 = ~n34909 | ~n34908;
  assign n34912 = ~n34911 | ~n34910;
  assign n34916 = ~n34913 | ~n34912;
  assign n34915 = ~n34914 | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign P2_U3602 = ~n34916 | ~n34915;
  assign n34919 = ~n34918 ^ n34917;
  assign n34922 = ~n34919 & ~n33538;
  assign n34921 = ~n34920 & ~n35967;
  assign n34924 = ~n34922 & ~n34921;
  assign n34923 = ~P2_EBX_REG_10__SCAN_IN | ~n35967;
  assign P2_U2877 = ~n34924 | ~n34923;
  assign n34926 = ~n34242 | ~n35010;
  assign n34925 = ~n39962 | ~n35011;
  assign n34930 = ~n34926 | ~n34925;
  assign n34928 = ~n39939 | ~n38889;
  assign n34927 = ~n39967 | ~n40037;
  assign n34929 = ~n34928 | ~n34927;
  assign n34932 = ~n34930 & ~n34929;
  assign n34931 = ~P1_INSTQUEUE_REG_15__0__SCAN_IN | ~n35014;
  assign P1_U3153 = ~n34932 | ~n34931;
  assign n34934 = ~n34165 | ~n35010;
  assign n34933 = ~n39995 | ~n35011;
  assign n34938 = ~n34934 | ~n34933;
  assign n34936 = ~n39992 | ~n38889;
  assign n34935 = ~n40000 | ~n40037;
  assign n34937 = ~n34936 | ~n34935;
  assign n34940 = ~n34938 & ~n34937;
  assign n34939 = ~P1_INSTQUEUE_REG_15__3__SCAN_IN | ~n35014;
  assign P1_U3156 = ~n34940 | ~n34939;
  assign n34942 = ~n34072 | ~n35010;
  assign n34941 = ~n40017 | ~n35011;
  assign n34946 = ~n34942 | ~n34941;
  assign n34944 = ~n40014 | ~n38889;
  assign n34943 = ~n40022 | ~n40037;
  assign n34945 = ~n34944 | ~n34943;
  assign n34948 = ~n34946 & ~n34945;
  assign n34947 = ~P1_INSTQUEUE_REG_15__7__SCAN_IN | ~n35014;
  assign P1_U3160 = ~n34948 | ~n34947;
  assign n34950 = ~n34188 | ~n35010;
  assign n34949 = ~n39973 | ~n35011;
  assign n34954 = ~n34950 | ~n34949;
  assign n34952 = ~n39970 | ~n38889;
  assign n34951 = ~n39978 | ~n40037;
  assign n34953 = ~n34952 | ~n34951;
  assign n34956 = ~n34954 & ~n34953;
  assign n34955 = ~P1_INSTQUEUE_REG_15__1__SCAN_IN | ~n35014;
  assign P1_U3154 = ~n34956 | ~n34955;
  assign n34958 = ~n34135 | ~n35010;
  assign n34957 = ~n39984 | ~n35011;
  assign n34962 = ~n34958 | ~n34957;
  assign n34960 = ~n39981 | ~n38889;
  assign n34959 = ~n39989 | ~n40037;
  assign n34961 = ~n34960 | ~n34959;
  assign n34964 = ~n34962 & ~n34961;
  assign n34963 = ~P1_INSTQUEUE_REG_15__4__SCAN_IN | ~n35014;
  assign P1_U3157 = ~n34964 | ~n34963;
  assign n34973 = ~n34965 & ~n35459;
  assign n35309 = ~n35307;
  assign n34970 = ~n34969 & ~n34968;
  assign n34971 = ~n35695 & ~n34970;
  assign n34972 = ~n35309 & ~n34971;
  assign n34975 = ~n34973 & ~n34972;
  assign n34974 = ~n35462 | ~BUF2_REG_14__SCAN_IN;
  assign P3_U2721 = ~n34975 | ~n34974;
  assign n38031 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n37011 = ~n34976;
  assign n34977 = ~n38031 | ~n37011;
  assign n37010 = ~n34978 | ~n34977;
  assign n34980 = ~n37011 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n34981 = ~n34980 & ~n34979;
  assign n34982 = n37010 ^ n34981;
  assign n34998 = ~n34982 & ~n35942;
  assign n34984 = ~P3_REIP_REG_17__SCAN_IN | ~n34983;
  assign n34994 = ~P3_REIP_REG_18__SCAN_IN & ~n34984;
  assign n34988 = ~n34985 & ~n36176;
  assign n34987 = ~n35944 | ~n34986;
  assign n34989 = ~n34988 & ~n34987;
  assign n34992 = ~n34990 & ~n34989;
  assign n34991 = ~P3_EBX_REG_18__SCAN_IN | ~n35935;
  assign n34993 = ~n34992 | ~n34991;
  assign n34996 = ~n34994 & ~n34993;
  assign n34995 = ~n36154 | ~P3_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n34997 = ~n34996 | ~n34995;
  assign n35001 = ~n34998 & ~n34997;
  assign n35000 = ~n34999 | ~P3_REIP_REG_18__SCAN_IN;
  assign P3_U2653 = ~n35001 | ~n35000;
  assign n35003 = ~n34227 | ~n35010;
  assign n35002 = ~n40006 | ~n35011;
  assign n35007 = ~n35003 | ~n35002;
  assign n35005 = ~P1_INSTQUEUE_REG_15__2__SCAN_IN | ~n35014;
  assign n35004 = ~n40003 | ~n38889;
  assign n35006 = ~n35005 | ~n35004;
  assign n35009 = ~n35007 & ~n35006;
  assign n35008 = ~n40011 | ~n40037;
  assign P1_U3155 = ~n35009 | ~n35008;
  assign n35013 = ~n34098 | ~n35010;
  assign n35012 = ~n40043 | ~n35011;
  assign n35018 = ~n35013 | ~n35012;
  assign n35016 = ~P1_INSTQUEUE_REG_15__5__SCAN_IN | ~n35014;
  assign n35015 = ~n40038 | ~n38889;
  assign n35017 = ~n35016 | ~n35015;
  assign n35020 = ~n35018 & ~n35017;
  assign n35019 = ~n40049 | ~n40037;
  assign P1_U3158 = ~n35020 | ~n35019;
  assign n39805 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n35021;
  assign n35022 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n39805;
  assign n35088 = ~n35022;
  assign n35027 = ~n34165 | ~n35088;
  assign n35025 = ~P1_STATE2_REG_2__SCAN_IN | ~n39805;
  assign n35023 = ~n39821 | ~n35165;
  assign n35024 = ~n39315 | ~n35033;
  assign n35026 = ~n39995 | ~n35089;
  assign n35031 = ~n35027 | ~n35026;
  assign n39879 = ~n35032 & ~n35172;
  assign n35029 = ~n39992 | ~n39879;
  assign n38894 = ~n35032 & ~n35173;
  assign n35028 = ~n40000 | ~n38894;
  assign n35030 = ~n35029 | ~n35028;
  assign n35039 = ~n35031 & ~n35030;
  assign n35036 = ~n39315 & ~n39805;
  assign n35034 = ~n35032 & ~n35178;
  assign n35035 = ~n35034 & ~n35033;
  assign n35037 = ~n35036 & ~n35035;
  assign n35038 = ~P1_INSTQUEUE_REG_13__3__SCAN_IN | ~n35096;
  assign P1_U3140 = ~n35039 | ~n35038;
  assign n35041 = ~n34098 | ~n35088;
  assign n35040 = ~n40043 | ~n35089;
  assign n35045 = ~n35041 | ~n35040;
  assign n35043 = ~n40038 | ~n39879;
  assign n35042 = ~n40049 | ~n38894;
  assign n35044 = ~n35043 | ~n35042;
  assign n35047 = ~n35045 & ~n35044;
  assign n35046 = ~P1_INSTQUEUE_REG_13__5__SCAN_IN | ~n35096;
  assign P1_U3142 = ~n35047 | ~n35046;
  assign n35049 = ~n39962 | ~n35089;
  assign n35048 = ~n34242 | ~n35088;
  assign n35053 = ~n35049 | ~n35048;
  assign n35051 = ~P1_INSTQUEUE_REG_13__0__SCAN_IN | ~n35096;
  assign n35050 = ~n39967 | ~n38894;
  assign n35052 = ~n35051 | ~n35050;
  assign n35055 = ~n35053 & ~n35052;
  assign n35054 = ~n39939 | ~n39879;
  assign P1_U3137 = ~n35055 | ~n35054;
  assign n35057 = ~n34150 | ~n35088;
  assign n35056 = ~n40028 | ~n35089;
  assign n35061 = ~n35057 | ~n35056;
  assign n35059 = ~n40025 | ~n39879;
  assign n35058 = ~n40033 | ~n38894;
  assign n35060 = ~n35059 | ~n35058;
  assign n35063 = ~n35061 & ~n35060;
  assign n35062 = ~P1_INSTQUEUE_REG_13__6__SCAN_IN | ~n35096;
  assign P1_U3143 = ~n35063 | ~n35062;
  assign n35065 = ~n34072 | ~n35088;
  assign n35064 = ~n40017 | ~n35089;
  assign n35069 = ~n35065 | ~n35064;
  assign n35067 = ~n40014 | ~n39879;
  assign n35066 = ~n40022 | ~n38894;
  assign n35068 = ~n35067 | ~n35066;
  assign n35071 = ~n35069 & ~n35068;
  assign n35070 = ~P1_INSTQUEUE_REG_13__7__SCAN_IN | ~n35096;
  assign P1_U3144 = ~n35071 | ~n35070;
  assign n35073 = ~n34227 | ~n35088;
  assign n35072 = ~n40006 | ~n35089;
  assign n35077 = ~n35073 | ~n35072;
  assign n35075 = ~n40003 | ~n39879;
  assign n35074 = ~n40011 | ~n38894;
  assign n35076 = ~n35075 | ~n35074;
  assign n35079 = ~n35077 & ~n35076;
  assign n35078 = ~P1_INSTQUEUE_REG_13__2__SCAN_IN | ~n35096;
  assign P1_U3139 = ~n35079 | ~n35078;
  assign n35081 = ~n34135 | ~n35088;
  assign n35080 = ~n39984 | ~n35089;
  assign n35085 = ~n35081 | ~n35080;
  assign n35083 = ~n39981 | ~n39879;
  assign n35082 = ~n39989 | ~n38894;
  assign n35084 = ~n35083 | ~n35082;
  assign n35087 = ~n35085 & ~n35084;
  assign n35086 = ~P1_INSTQUEUE_REG_13__4__SCAN_IN | ~n35096;
  assign P1_U3141 = ~n35087 | ~n35086;
  assign n35091 = ~n34188 | ~n35088;
  assign n35090 = ~n39973 | ~n35089;
  assign n35095 = ~n35091 | ~n35090;
  assign n35093 = ~n39970 | ~n39879;
  assign n35092 = ~n39978 | ~n38894;
  assign n35094 = ~n35093 | ~n35092;
  assign n35098 = ~n35095 & ~n35094;
  assign n35097 = ~P1_INSTQUEUE_REG_13__1__SCAN_IN | ~n35096;
  assign P1_U3138 = ~n35098 | ~n35097;
  assign n35103 = ~n36895 & ~n35099;
  assign n35101 = ~n36891 | ~n35100;
  assign n35102 = ~n36893 | ~n35101;
  assign n36120 = ~n35103 & ~n35102;
  assign n35107 = ~n35104 & ~n36120;
  assign n35689 = ~n43469 | ~P1_REIP_REG_6__SCAN_IN;
  assign n35105 = ~n44014 | ~n43344;
  assign n35106 = ~n35689 | ~n35105;
  assign n35119 = ~n35107 & ~n35106;
  assign n35111 = n35109 | n35108;
  assign n35117 = ~n43341 & ~n35682;
  assign n35115 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN & ~P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n36129 = ~n35361 & ~n35112;
  assign n35114 = ~n36129 | ~n35113;
  assign n35116 = ~n35115 & ~n35114;
  assign n35118 = ~n35117 & ~n35116;
  assign P1_U3025 = ~n35119 | ~n35118;
  assign n35121 = ~n34072 | ~n35152;
  assign n35120 = ~n40014 | ~n39107;
  assign n35125 = ~n35121 | ~n35120;
  assign n35123 = ~P1_INSTQUEUE_REG_3__7__SCAN_IN | ~n35155;
  assign n35122 = ~n40017 | ~n35156;
  assign n35124 = ~n35123 | ~n35122;
  assign n35127 = ~n35125 & ~n35124;
  assign n35126 = ~n40022 | ~n38478;
  assign P1_U3064 = ~n35127 | ~n35126;
  assign n35129 = ~n34098 | ~n35152;
  assign n35128 = ~n40038 | ~n39107;
  assign n35133 = ~n35129 | ~n35128;
  assign n35131 = ~P1_INSTQUEUE_REG_3__5__SCAN_IN | ~n35155;
  assign n35130 = ~n40043 | ~n35156;
  assign n35132 = ~n35131 | ~n35130;
  assign n35135 = ~n35133 & ~n35132;
  assign n35134 = ~n40049 | ~n38478;
  assign P1_U3062 = ~n35135 | ~n35134;
  assign n35137 = ~n34135 | ~n35152;
  assign n35136 = ~n39981 | ~n39107;
  assign n35141 = ~n35137 | ~n35136;
  assign n35139 = ~P1_INSTQUEUE_REG_3__4__SCAN_IN | ~n35155;
  assign n35138 = ~n39984 | ~n35156;
  assign n35140 = ~n35139 | ~n35138;
  assign n35143 = ~n35141 & ~n35140;
  assign n35142 = ~n39989 | ~n38478;
  assign P1_U3061 = ~n35143 | ~n35142;
  assign n35145 = ~n34165 | ~n35152;
  assign n35144 = ~n39992 | ~n39107;
  assign n35149 = ~n35145 | ~n35144;
  assign n35147 = ~P1_INSTQUEUE_REG_3__3__SCAN_IN | ~n35155;
  assign n35146 = ~n39995 | ~n35156;
  assign n35148 = ~n35147 | ~n35146;
  assign n35151 = ~n35149 & ~n35148;
  assign n35150 = ~n40000 | ~n38478;
  assign P1_U3060 = ~n35151 | ~n35150;
  assign n35154 = ~n34242 | ~n35152;
  assign n35153 = ~n39939 | ~n39107;
  assign n35160 = ~n35154 | ~n35153;
  assign n35158 = ~P1_INSTQUEUE_REG_3__0__SCAN_IN | ~n35155;
  assign n35157 = ~n39962 | ~n35156;
  assign n35159 = ~n35158 | ~n35157;
  assign n35162 = ~n35160 & ~n35159;
  assign n35161 = ~n39967 | ~n38478;
  assign P1_U3057 = ~n35162 | ~n35161;
  assign n35164 = ~n35163 | ~n37475;
  assign n39938 = ~n35164 & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n35166 = ~n39938 | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n35236 = ~n35166;
  assign n35171 = ~n34165 | ~n35236;
  assign n35169 = ~P1_STATE2_REG_2__SCAN_IN | ~n39938;
  assign n35167 = ~n39959 | ~n35165;
  assign n35168 = ~n39315 | ~n35180;
  assign n35170 = ~n39995 | ~n35237;
  assign n35177 = ~n35171 | ~n35170;
  assign n40048 = ~n35179 & ~n35172;
  assign n35175 = ~n39992 | ~n40048;
  assign n39102 = ~n35179 & ~n35173;
  assign n35174 = ~n40000 | ~n39102;
  assign n35176 = ~n35175 | ~n35174;
  assign n35187 = ~n35177 & ~n35176;
  assign n35183 = ~n39315 & ~n39938;
  assign n35181 = ~n35179 & ~n35178;
  assign n35182 = ~n35181 & ~n35180;
  assign n35184 = ~n35183 & ~n35182;
  assign n35186 = ~P1_INSTQUEUE_REG_1__3__SCAN_IN | ~n35244;
  assign P1_U3044 = ~n35187 | ~n35186;
  assign n35189 = ~n34188 | ~n35236;
  assign n35188 = ~n39973 | ~n35237;
  assign n35193 = ~n35189 | ~n35188;
  assign n35191 = ~n39970 | ~n40048;
  assign n35190 = ~n39978 | ~n39102;
  assign n35192 = ~n35191 | ~n35190;
  assign n35195 = ~n35193 & ~n35192;
  assign n35194 = ~P1_INSTQUEUE_REG_1__1__SCAN_IN | ~n35244;
  assign P1_U3042 = ~n35195 | ~n35194;
  assign n35197 = ~n34150 | ~n35236;
  assign n35196 = ~n40028 | ~n35237;
  assign n35201 = ~n35197 | ~n35196;
  assign n35199 = ~n40025 | ~n40048;
  assign n35198 = ~n40033 | ~n39102;
  assign n35200 = ~n35199 | ~n35198;
  assign n35203 = ~n35201 & ~n35200;
  assign n35202 = ~P1_INSTQUEUE_REG_1__6__SCAN_IN | ~n35244;
  assign P1_U3047 = ~n35203 | ~n35202;
  assign n35205 = ~n34098 | ~n35236;
  assign n35204 = ~n40043 | ~n35237;
  assign n35209 = ~n35205 | ~n35204;
  assign n35207 = ~n40038 | ~n40048;
  assign n35206 = ~n40049 | ~n39102;
  assign n35208 = ~n35207 | ~n35206;
  assign n35211 = ~n35209 & ~n35208;
  assign n35210 = ~P1_INSTQUEUE_REG_1__5__SCAN_IN | ~n35244;
  assign P1_U3046 = ~n35211 | ~n35210;
  assign n35213 = ~n39962 | ~n35237;
  assign n35212 = ~n34242 | ~n35236;
  assign n35217 = ~n35213 | ~n35212;
  assign n35215 = ~n39939 | ~n40048;
  assign n35214 = ~n39967 | ~n39102;
  assign n35216 = ~n35215 | ~n35214;
  assign n35219 = ~n35217 & ~n35216;
  assign n35218 = ~P1_INSTQUEUE_REG_1__0__SCAN_IN | ~n35244;
  assign P1_U3041 = ~n35219 | ~n35218;
  assign n35221 = ~n34135 | ~n35236;
  assign n35220 = ~n39984 | ~n35237;
  assign n35225 = ~n35221 | ~n35220;
  assign n35223 = ~n39981 | ~n40048;
  assign n35222 = ~n39989 | ~n39102;
  assign n35224 = ~n35223 | ~n35222;
  assign n35227 = ~n35225 & ~n35224;
  assign n35226 = ~P1_INSTQUEUE_REG_1__4__SCAN_IN | ~n35244;
  assign P1_U3045 = ~n35227 | ~n35226;
  assign n35229 = ~n34072 | ~n35236;
  assign n35228 = ~n40017 | ~n35237;
  assign n35233 = ~n35229 | ~n35228;
  assign n35231 = ~n40014 | ~n40048;
  assign n35230 = ~n40022 | ~n39102;
  assign n35232 = ~n35231 | ~n35230;
  assign n35235 = ~n35233 & ~n35232;
  assign n35234 = ~P1_INSTQUEUE_REG_1__7__SCAN_IN | ~n35244;
  assign P1_U3048 = ~n35235 | ~n35234;
  assign n35239 = ~n34227 | ~n35236;
  assign n35238 = ~n40006 | ~n35237;
  assign n35243 = ~n35239 | ~n35238;
  assign n35241 = ~n40003 | ~n40048;
  assign n35240 = ~n40011 | ~n39102;
  assign n35242 = ~n35241 | ~n35240;
  assign n35246 = ~n35243 & ~n35242;
  assign n35245 = ~P1_INSTQUEUE_REG_1__2__SCAN_IN | ~n35244;
  assign P1_U3043 = ~n35246 | ~n35245;
  assign n35248 = ~n40580 | ~n43523;
  assign n35247 = ~n35967 | ~P2_EBX_REG_4__SCAN_IN;
  assign n35252 = n35248 & n35247;
  assign n40565 = n35250 ^ n35249;
  assign n35251 = ~n40565 | ~n43525;
  assign P2_U2883 = ~n35252 | ~n35251;
  assign n35257 = ~n35253 | ~n43523;
  assign n35255 = ~n36253 & ~n35254;
  assign n35256 = ~n35255 & ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n35260 = ~n35257 & ~n35256;
  assign n35258 = ~P2_EBX_REG_7__SCAN_IN;
  assign n35259 = ~n43525 & ~n35258;
  assign n35264 = ~n35260 & ~n35259;
  assign n40943 = ~n35262 ^ n35261;
  assign n37339 = ~n40943;
  assign n35263 = ~n37339 | ~n43525;
  assign P2_U2880 = ~n35264 | ~n35263;
  assign n35266 = ~n42011 & ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n35265 = ~n35452 & ~P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n35271 = ~n35266 & ~n35265;
  assign n35269 = ~n40968 | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n35610 = ~n35267 & ~n42320;
  assign n35268 = n35610 | P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n35270 = ~n36057 | ~n41345;
  assign n35272 = ~n35271 | ~n35270;
  assign n35274 = ~n36061 | ~n35272;
  assign n35273 = ~n36063 | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign P3_U3290 = ~n35274 | ~n35273;
  assign n35276 = ~n34098 | ~n35350;
  assign n35275 = ~n40043 | ~n35351;
  assign n35280 = ~n35276 | ~n35275;
  assign n35278 = ~n40038 | ~n38562;
  assign n35277 = ~n40049 | ~n39374;
  assign n35279 = ~n35278 | ~n35277;
  assign n35282 = ~n35280 & ~n35279;
  assign n35281 = ~P1_INSTQUEUE_REG_7__5__SCAN_IN | ~n35354;
  assign P1_U3094 = ~n35282 | ~n35281;
  assign n35284 = ~n34188 | ~n35350;
  assign n35283 = ~n39973 | ~n35351;
  assign n35288 = ~n35284 | ~n35283;
  assign n35286 = ~n39970 | ~n38562;
  assign n35285 = ~n39978 | ~n39374;
  assign n35287 = ~n35286 | ~n35285;
  assign n35290 = ~n35288 & ~n35287;
  assign n35289 = ~P1_INSTQUEUE_REG_7__1__SCAN_IN | ~n35354;
  assign P1_U3090 = ~n35290 | ~n35289;
  assign n35292 = ~n34135 | ~n35350;
  assign n35291 = ~n39984 | ~n35351;
  assign n35296 = ~n35292 | ~n35291;
  assign n35294 = ~n39981 | ~n38562;
  assign n35293 = ~n39989 | ~n39374;
  assign n35295 = ~n35294 | ~n35293;
  assign n35298 = ~n35296 & ~n35295;
  assign n35297 = ~P1_INSTQUEUE_REG_7__4__SCAN_IN | ~n35354;
  assign P1_U3093 = ~n35298 | ~n35297;
  assign n35300 = ~n34227 | ~n35350;
  assign n35299 = ~n40006 | ~n35351;
  assign n35304 = ~n35300 | ~n35299;
  assign n35302 = ~n40003 | ~n38562;
  assign n35301 = ~n40011 | ~n39374;
  assign n35303 = ~n35302 | ~n35301;
  assign n35306 = ~n35304 & ~n35303;
  assign n35305 = ~P1_INSTQUEUE_REG_7__2__SCAN_IN | ~n35354;
  assign P1_U3091 = ~n35306 | ~n35305;
  assign n35698 = ~n36243 | ~n35307;
  assign n35313 = ~n35697 & ~n35698;
  assign n35311 = ~n36333 | ~n35308;
  assign n35310 = ~n35309 | ~n35697;
  assign n35312 = ~n35311 | ~n35310;
  assign n35315 = ~n35313 & ~n35312;
  assign n35314 = ~n35462 | ~BUF2_REG_15__SCAN_IN;
  assign P3_U2720 = ~n35315 | ~n35314;
  assign n35319 = n42219 & n35381;
  assign n35318 = ~n36002 & ~n35317;
  assign n35320 = ~P2_EAX_REG_15__SCAN_IN | ~n43698;
  assign P2_U2904 = ~n35321 | ~n35320;
  assign n35328 = ~n35327;
  assign n35333 = ~n35331;
  assign n35337 = ~n43358 & ~n35363;
  assign n35370 = ~P1_REIP_REG_4__SCAN_IN | ~n43469;
  assign n35335 = ~n43709 | ~P1_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n35336 = ~n35370 | ~n35335;
  assign n35341 = ~n35337 & ~n35336;
  assign n35339 = ~n35518 & ~n43713;
  assign n35338 = ~n35517 & ~n43729;
  assign n35340 = ~n35339 & ~n35338;
  assign P1_U2995 = ~n35341 | ~n35340;
  assign n35343 = ~n34242 | ~n35350;
  assign n35342 = ~n39962 | ~n35351;
  assign n35347 = ~n35343 | ~n35342;
  assign n35345 = ~P1_INSTQUEUE_REG_7__0__SCAN_IN | ~n35354;
  assign n35344 = ~n39939 | ~n38562;
  assign n35346 = ~n35345 | ~n35344;
  assign n35349 = ~n35347 & ~n35346;
  assign n35348 = ~n39967 | ~n39374;
  assign P1_U3089 = ~n35349 | ~n35348;
  assign n35353 = ~n34072 | ~n35350;
  assign n35352 = ~n40017 | ~n35351;
  assign n35358 = ~n35353 | ~n35352;
  assign n35356 = ~P1_INSTQUEUE_REG_7__7__SCAN_IN | ~n35354;
  assign n35355 = ~n40014 | ~n38562;
  assign n35357 = ~n35356 | ~n35355;
  assign n35360 = ~n35358 & ~n35357;
  assign n35359 = ~n40022 | ~n39374;
  assign P1_U3096 = ~n35360 | ~n35359;
  assign n35362 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN & ~n35361;
  assign n35375 = ~n35362 | ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n35373 = ~n43341 & ~n35363;
  assign n35369 = ~n43441 & ~n35503;
  assign n35367 = ~n35365 & ~n35364;
  assign n35368 = ~n35367 & ~n35366;
  assign n35371 = ~n35369 & ~n35368;
  assign n35372 = ~n35371 | ~n35370;
  assign n35374 = ~n35373 & ~n35372;
  assign P1_U3027 = ~n35375 | ~n35374;
  assign n35383 = ~n36002 & ~n43696;
  assign n35379 = ~n35378 & ~n35377;
  assign n35382 = n42665 & n35381;
  assign n35385 = ~n35383 & ~n35382;
  assign n35384 = ~P2_EAX_REG_14__SCAN_IN | ~n43698;
  assign P2_U2905 = ~n35385 | ~n35384;
  assign n35387 = ~n36320 | ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n35386 = ~n22923 | ~P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n35391 = ~n35387 | ~n35386;
  assign n35389 = ~n22909 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n35388 = ~n22913 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n35390 = ~n35389 | ~n35388;
  assign n35418 = ~n35391 & ~n35390;
  assign n35394 = ~n22902 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n35393 = ~n35392 | ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n35398 = ~n35394 | ~n35393;
  assign n35396 = ~n36294 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n35395 = ~n22917 | ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n35397 = ~n35396 | ~n35395;
  assign n35406 = ~n35398 & ~n35397;
  assign n35400 = ~n22903 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n35399 = ~n36317 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n35404 = ~n35400 | ~n35399;
  assign n35402 = ~n36307 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n35401 = ~n36311 | ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n35403 = ~n35402 | ~n35401;
  assign n35405 = ~n35404 & ~n35403;
  assign n35416 = ~n35406 | ~n35405;
  assign n35410 = n22922 | n35407;
  assign n35409 = ~n22910 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n35414 = ~n35410 | ~n35409;
  assign n35412 = ~n22919 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n35411 = ~n22914 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n35413 = ~n35412 | ~n35411;
  assign n35415 = n35414 | n35413;
  assign n35417 = ~n35416 & ~n35415;
  assign n35691 = ~n35418 | ~n35417;
  assign n35424 = ~n42135 | ~n35691;
  assign n35419 = ~P3_EBX_REG_16__SCAN_IN | ~n43930;
  assign n35422 = ~n35419 | ~n35421;
  assign n35423 = ~n35422 | ~n35551;
  assign P3_U2687 = ~n35424 | ~n35423;
  assign n35427 = ~n35426 & ~n35425;
  assign n35428 = ~n35427 & ~n33538;
  assign n35430 = ~n35428 | ~n35599;
  assign n35429 = ~n35967 | ~P2_EBX_REG_11__SCAN_IN;
  assign n35434 = n35430 & n35429;
  assign n35433 = ~n42565 | ~n43525;
  assign P2_U2876 = ~n35434 | ~n35433;
  assign n36527 = ~n40865 & ~n35904;
  assign n37089 = ~n41095;
  assign n35441 = ~n37089 & ~P3_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n35438 = ~n35437 | ~n35436;
  assign n36515 = ~n35439 | ~n35438;
  assign n35440 = ~n41397 & ~n36515;
  assign n35450 = ~n35441 & ~n35440;
  assign n35444 = ~P3_STATE2_REG_0__SCAN_IN & ~n35442;
  assign n37753 = ~n35444 & ~n35443;
  assign n35448 = ~n40734 & ~n36661;
  assign n36516 = ~n35446 ^ n35445;
  assign n35447 = ~n36914 & ~n36516;
  assign n35449 = ~n35448 & ~n35447;
  assign n35451 = ~n35450 | ~n35449;
  assign n35454 = ~n36527 & ~n35451;
  assign n40731 = ~P3_STATE2_REG_1__SCAN_IN | ~P3_STATEBS16_REG_SCAN_IN;
  assign n41400 = ~n35452 & ~n36660;
  assign n35923 = ~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~n36661;
  assign n35925 = ~P3_PHYADDRPOINTER_REG_2__SCAN_IN | ~n36220;
  assign n35910 = ~n35923 | ~n35925;
  assign n35453 = ~n36871 | ~n35910;
  assign P3_U2828 = ~n35454 | ~n35453;
  assign n35455 = ~P3_EAX_REG_13__SCAN_IN | ~n36243;
  assign n35457 = n35456 & n35455;
  assign n35461 = ~n35695 & ~n35457;
  assign n35460 = ~n35459 & ~n35458;
  assign n35464 = ~n35461 & ~n35460;
  assign n35463 = ~BUF2_REG_13__SCAN_IN | ~n35462;
  assign P3_U2722 = ~n35464 | ~n35463;
  assign n35467 = ~n35466 & ~n35465;
  assign n35481 = ~n35468 & ~n36143;
  assign n35469 = ~n41129 | ~n42175;
  assign n35479 = ~n35469 | ~P1_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n35472 = ~n35470 | ~n43803;
  assign n35471 = ~n43796 | ~P1_EBX_REG_0__SCAN_IN;
  assign n35477 = ~n35472 | ~n35471;
  assign n36135 = ~n35474 | ~n35473;
  assign n35476 = ~n35475 & ~n36135;
  assign n35478 = ~n35477 & ~n35476;
  assign n35480 = ~n35479 | ~n35478;
  assign n35483 = ~n35481 & ~n35480;
  assign n35482 = ~P1_REIP_REG_0__SCAN_IN | ~n35512;
  assign P1_U2840 = ~n35483 | ~n35482;
  assign n35491 = ~n35484 & ~n36143;
  assign n35487 = ~n43570 & ~n35485;
  assign n35486 = ~n39942 & ~n36135;
  assign n35489 = ~n35487 & ~n35486;
  assign n35488 = ~P1_EBX_REG_1__SCAN_IN | ~n43796;
  assign n35490 = ~n35489 | ~n35488;
  assign n35499 = ~n35491 & ~n35490;
  assign n35497 = ~P1_PHYADDRPOINTER_REG_1__SCAN_IN & ~n42175;
  assign n35493 = ~n41894 & ~n35494;
  assign n35492 = P1_PHYADDRPOINTER_REG_1__SCAN_IN & n43797;
  assign n35495 = ~n35493 & ~n35492;
  assign n36141 = ~n42405 | ~n35494;
  assign n35496 = ~n35495 | ~n36141;
  assign n35498 = ~n35497 & ~n35496;
  assign P1_U2839 = ~n35499 | ~n35498;
  assign n35516 = ~n36135 & ~n35500;
  assign n35511 = ~n35501 | ~n41894;
  assign n36107 = ~n42405 | ~n35502;
  assign n35510 = ~n35511 & ~n36107;
  assign n35506 = ~n43570 & ~n35503;
  assign n35504 = ~P1_PHYADDRPOINTER_REG_4__SCAN_IN | ~n43797;
  assign n35505 = ~n35504 | ~n43033;
  assign n35508 = ~n35506 & ~n35505;
  assign n35507 = ~P1_EBX_REG_4__SCAN_IN | ~n43796;
  assign n35509 = ~n35508 | ~n35507;
  assign n35514 = ~n35510 & ~n35509;
  assign n35878 = n35512 & n35511;
  assign n35513 = ~P1_REIP_REG_4__SCAN_IN | ~n35878;
  assign n35522 = ~n35516 & ~n35515;
  assign n35520 = ~n35517 & ~n36143;
  assign n35519 = ~n35518 & ~n42175;
  assign n35521 = ~n35520 & ~n35519;
  assign P1_U2836 = ~n35522 | ~n35521;
  assign n35524 = ~n35542 & ~n35523;
  assign n35949 = ~P3_REIP_REG_28__SCAN_IN | ~n35524;
  assign n35547 = ~n35543 & ~n35644;
  assign n41682 = ~P3_EBX_REG_28__SCAN_IN;
  assign n35540 = ~n35945 & ~n41682;
  assign n35526 = ~n41682 & ~n35527;
  assign n35528 = ~n35526 & ~n35642;
  assign n35538 = ~n35528 | ~n35641;
  assign n35530 = ~n41158 & ~n35529;
  assign n35531 = ~P3_PHYADDRPOINTER_REG_28__SCAN_IN & ~n35530;
  assign n40864 = ~n35531 & ~n35654;
  assign n35535 = ~n40864;
  assign n35533 = ~n35535 & ~n35534;
  assign n35536 = ~n35533 & ~n35942;
  assign n35537 = ~n35536 | ~n35656;
  assign n35539 = ~n35538 | ~n35537;
  assign n35545 = ~n35540 & ~n35539;
  assign n35640 = ~n35542 & ~n35541;
  assign n35544 = ~n35640 | ~n35543;
  assign n35549 = ~n35547 & ~n35546;
  assign n35548 = ~n36154 | ~P3_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign P3_U2643 = ~n35549 | ~n35548;
  assign n35556 = ~n42135 | ~n35550;
  assign n35552 = ~P3_EBX_REG_17__SCAN_IN | ~n43930;
  assign n35554 = ~n35552 | ~n35551;
  assign P3_U2686 = ~n35556 | ~n35555;
  assign n35592 = BUF2_REG_29__SCAN_IN & n36282;
  assign n35558 = ~n22919 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n35557 = ~n22903 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n35562 = ~n35558 | ~n35557;
  assign n35560 = ~n22914 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n35559 = ~n36307 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n35561 = ~n35560 | ~n35559;
  assign n35570 = ~n35562 & ~n35561;
  assign n35564 = ~n22902 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n35563 = ~n36317 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n35568 = ~n35564 | ~n35563;
  assign n35566 = ~n36320 | ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n35565 = ~n22920 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n35567 = ~n35566 | ~n35565;
  assign n35569 = ~n35568 & ~n35567;
  assign n35586 = ~n35570 | ~n35569;
  assign n35572 = ~n36294 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n35571 = ~n36298 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n35576 = ~n35572 | ~n35571;
  assign n35574 = ~n36310 | ~P3_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n35573 = ~n22913 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n35575 = ~n35574 | ~n35573;
  assign n35584 = ~n35576 & ~n35575;
  assign n35578 = ~n35392 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n35577 = ~n36311 | ~P3_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n35582 = ~n35578 | ~n35577;
  assign n35580 = ~n22917 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n35579 = ~n22923 | ~P3_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n35581 = ~n35580 | ~n35579;
  assign n35583 = ~n35582 & ~n35581;
  assign n35585 = ~n35584 | ~n35583;
  assign n36330 = ~n35586 & ~n35585;
  assign n36329 = ~n35588 | ~n35587;
  assign n41862 = n36330 ^ n36329;
  assign n35590 = ~n36333 | ~n41862;
  assign n35589 = ~n36338 | ~BUF2_REG_13__SCAN_IN;
  assign n35591 = ~n35590 | ~n35589;
  assign n35597 = ~n35592 & ~n35591;
  assign n35593 = ~P3_EAX_REG_29__SCAN_IN | ~n36243;
  assign n35595 = ~n35593 | ~n35594;
  assign n35596 = ~n35595 | ~n36283;
  assign P3_U2706 = ~n35597 | ~n35596;
  assign n35600 = ~n35599 ^ n35598;
  assign n35605 = ~n35600 & ~n33538;
  assign n35603 = ~n42452;
  assign n35604 = ~n35603 & ~n35967;
  assign n35607 = ~n35605 & ~n35604;
  assign n35606 = ~P2_EBX_REG_12__SCAN_IN | ~n35967;
  assign P2_U2875 = ~n35607 | ~n35606;
  assign n35612 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~n36038;
  assign n35611 = ~n35610 & ~n35613;
  assign n35615 = ~n35670 & ~n41342;
  assign n35614 = ~n42011 & ~n35613;
  assign n35618 = ~n35615 & ~n35614;
  assign n35671 = ~P3_STATE2_REG_1__SCAN_IN | ~P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n35616 = ~n35671;
  assign n35672 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN ^ P3_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n35617 = ~n35616 | ~n35672;
  assign n35619 = ~n35618 | ~n35617;
  assign n35621 = ~n36061 | ~n35619;
  assign n35620 = ~n36063 | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign P3_U3289 = ~n35621 | ~n35620;
  assign n35625 = ~n35623 & ~n35622;
  assign n35639 = ~n35625 & ~n35624;
  assign n35637 = ~n35627 & ~n35626;
  assign n35628 = P1_STATE2_REG_0__SCAN_IN & n44100;
  assign n35629 = ~n35628 | ~n43722;
  assign n35635 = ~n44106 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n35632 = ~n35631 & ~n35630;
  assign n35633 = ~n35632 & ~P1_STATE2_REG_0__SCAN_IN;
  assign n35634 = ~n35633 | ~n44098;
  assign n35636 = ~n35635 | ~n35634;
  assign n35638 = ~n35637 & ~n35636;
  assign P1_U3161 = ~n35639 | ~n35638;
  assign n35653 = ~P3_REIP_REG_29__SCAN_IN & ~n36158;
  assign n35643 = ~P3_EBX_REG_29__SCAN_IN | ~n35641;
  assign n35943 = ~P3_EBX_REG_29__SCAN_IN & ~n35641;
  assign n35960 = ~n35943 & ~n35642;
  assign n35651 = ~n35643 | ~n35960;
  assign n35649 = ~n35645 & ~n35644;
  assign n35647 = ~P3_PHYADDRPOINTER_REG_29__SCAN_IN | ~n36154;
  assign n35646 = ~P3_EBX_REG_29__SCAN_IN | ~n35935;
  assign n35648 = ~n35647 | ~n35646;
  assign n35650 = ~n35649 & ~n35648;
  assign n35652 = ~n35651 | ~n35650;
  assign n35661 = ~n35653 & ~n35652;
  assign n41096 = ~P3_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n41099 = ~n35654;
  assign n35655 = ~n41096 | ~n41099;
  assign n41105 = ~n41402 | ~n35655;
  assign n35657 = ~n41105 & ~n35658;
  assign n35659 = ~n35657 & ~n35942;
  assign P3_U2642 = ~n35661 | ~n35660;
  assign n35662 = ~n36048 & ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n35906 = ~n35662 & ~n36040;
  assign n35669 = ~n40442 & ~n35906;
  assign n35664 = n35663 ^ P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n35665 = ~n36049 | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n35666 = ~n41537 & ~n35665;
  assign n35668 = n35667 | n35666;
  assign n35674 = ~n35670 & ~n41329;
  assign n35673 = ~n35672 & ~n35671;
  assign n35677 = ~n35674 & ~n35673;
  assign n35675 = ~n42011;
  assign n35676 = ~n35906 | ~n35675;
  assign n35678 = ~n35677 | ~n35676;
  assign n35680 = ~n36061 | ~n35678;
  assign n35679 = ~n36063 | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign P3_U3288 = ~n35680 | ~n35679;
  assign n35688 = ~n43713 & ~n35681;
  assign n35684 = ~n44013 & ~n43729;
  assign n35683 = ~n43358 & ~n35682;
  assign n35686 = ~n35684 & ~n35683;
  assign n35685 = ~P1_PHYADDRPOINTER_REG_6__SCAN_IN | ~n43709;
  assign n35690 = ~n35688 & ~n35687;
  assign P1_U2993 = ~n35690 | ~n35689;
  assign n35693 = ~BUF2_REG_16__SCAN_IN | ~n36282;
  assign n35692 = ~n36333 | ~n35691;
  assign n35704 = ~n35693 | ~n35692;
  assign n35696 = ~n35694 & ~P3_EAX_REG_16__SCAN_IN;
  assign n35702 = ~n35696 | ~n35695;
  assign n35699 = ~n36242 | ~n35697;
  assign n35700 = ~n35699 | ~n35698;
  assign n35701 = ~n35700 | ~P3_EAX_REG_16__SCAN_IN;
  assign n35703 = ~n35702 | ~n35701;
  assign n35706 = ~n35704 & ~n35703;
  assign n35705 = ~BUF2_REG_0__SCAN_IN | ~n36338;
  assign P3_U2719 = ~n35706 | ~n35705;
  assign n35713 = ~n35707 & ~n41877;
  assign n35710 = ~n35709;
  assign n35712 = ~n35711 | ~n35710;
  assign n36358 = ~n35713 & ~n35712;
  assign n35717 = ~n35719 | ~n35714;
  assign n35716 = ~n35766 | ~n35715;
  assign n35736 = ~n35719 & ~n35718;
  assign n35734 = ~n35720 & ~n35750;
  assign n35723 = ~n43484 & ~n35721;
  assign n35727 = ~n35722 | ~n35723;
  assign n35724 = ~n35723;
  assign n35726 = ~n35725 | ~n35724;
  assign n35732 = ~n35727 | ~n35726;
  assign n35730 = ~n35729 & ~n35728;
  assign n35731 = ~n35752 | ~n35730;
  assign n35733 = ~n35732 | ~n35731;
  assign n36497 = ~n35734 & ~n35733;
  assign n35735 = ~n35766 & ~n36497;
  assign n35748 = ~n35772 & ~n35769;
  assign n35737 = ~P2_FLUSH_REG_SCAN_IN & ~P2_MORE_REG_SCAN_IN;
  assign n35739 = ~n35738 & ~n35737;
  assign n35741 = ~n35740 & ~n35739;
  assign n35743 = ~n35742 | ~n35741;
  assign n35746 = ~n35744 & ~n35743;
  assign n35745 = ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n35766;
  assign n35747 = ~n35746 | ~n35745;
  assign n35779 = ~n35748 & ~n35747;
  assign n35768 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~n35769;
  assign n35761 = ~n39114 & ~n35749;
  assign n35764 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n35761;
  assign n35760 = ~n37302 & ~n35750;
  assign n35754 = ~n35751 | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n35753 = n35752 | P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n35758 = ~n35754 | ~n35753;
  assign n35757 = ~n35756 | ~n35755;
  assign n35759 = ~n35758 | ~n35757;
  assign n36531 = ~n35760 & ~n35759;
  assign n35762 = P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & n35761;
  assign n35763 = ~n36531 & ~n35762;
  assign n35765 = ~n35764 & ~n35763;
  assign n35767 = ~n35766 & ~n35765;
  assign n35770 = P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | n35769;
  assign n35773 = ~n35774 | ~n38277;
  assign n35775 = ~n35774 & ~n38277;
  assign n35776 = ~n35775 & ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign P2_U3593 = ~n35800 | ~n35781;
  assign n35783 = ~n43164 | ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n35794 = ~n35783 | ~n35782;
  assign n35789 = ~n43893 & ~n35784;
  assign n35787 = ~n43583 | ~n37303;
  assign n35786 = ~n43876 | ~n35785;
  assign n35788 = ~n35787 | ~n35786;
  assign n35792 = ~n35789 & ~n35788;
  assign n35791 = ~n43767 | ~n35790;
  assign n35793 = ~n35792 | ~n35791;
  assign n35799 = ~n35794 & ~n35793;
  assign n35795 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN & ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n35797 = ~n35796 & ~n35795;
  assign n35798 = ~n35797 | ~n43165;
  assign P2_U3045 = ~n35799 | ~n35798;
  assign n35810 = ~n35801 & ~n35800;
  assign n35803 = ~n39511 | ~n35802;
  assign n36360 = ~n35803 & ~n36357;
  assign n35808 = ~n35804 & ~n36360;
  assign n35807 = ~n35806 | ~n35805;
  assign n35809 = ~n35808 | ~n35807;
  assign n35818 = ~n35810 & ~n35809;
  assign n35813 = ~n36358;
  assign n35812 = n35811 | n36533;
  assign n35814 = ~n35813 | ~n35812;
  assign n35815 = ~n35814 | ~n36357;
  assign n35817 = ~n35816 | ~n35815;
  assign P2_U3176 = ~n35818 | ~n35817;
  assign n35827 = ~n36269 & ~n44019;
  assign n35825 = ~n35821;
  assign n35824 = ~n35823 | ~n35822;
  assign n36981 = ~n35825 | ~n35824;
  assign n35826 = ~n36981 & ~n43298;
  assign n35829 = ~n35827 & ~n35826;
  assign n35828 = ~P1_EBX_REG_7__SCAN_IN | ~n44023;
  assign P1_U2865 = ~n35829 | ~n35828;
  assign n36263 = ~n43033 & ~n36991;
  assign n35830 = ~n43441 & ~n36981;
  assign n35839 = ~n36263 & ~n35830;
  assign n35837 = ~P1_INSTADDRPOINTER_REG_7__SCAN_IN & ~n36890;
  assign n35835 = ~n36906 | ~n36264;
  assign n35834 = ~P1_INSTADDRPOINTER_REG_7__SCAN_IN | ~n35833;
  assign P1_U3024 = ~n35839 | ~n35838;
  assign n40961 = ~n40981 & ~n40403;
  assign n40969 = ~n40961;
  assign n36447 = ~n40959;
  assign n40387 = ~n40969 & ~n40503;
  assign n35841 = ~n41408 & ~n40387;
  assign n35840 = ~n41397 & ~n40388;
  assign n35855 = ~n40403 & ~n37085;
  assign n36068 = ~n41095 | ~n36415;
  assign n36434 = ~n36068;
  assign n35851 = ~n35842 | ~n36434;
  assign n35844 = n36660 & n35851;
  assign n35843 = ~n41403 & ~n35849;
  assign n37092 = ~n35844 & ~n35843;
  assign n35848 = ~n37092 & ~n37090;
  assign n35846 = ~n35845 | ~n41400;
  assign n40406 = ~n41145 | ~P3_REIP_REG_12__SCAN_IN;
  assign n35847 = ~n35846 | ~n40406;
  assign n35853 = ~n35848 & ~n35847;
  assign n35850 = ~n40726 | ~n35849;
  assign n37094 = ~n35851 | ~n35850;
  assign n35852 = ~n37094 | ~n37090;
  assign n35854 = ~n35853 | ~n35852;
  assign n35868 = ~n35855 & ~n35854;
  assign n40377 = ~n40127 | ~n40403;
  assign n35857 = ~n41397 & ~n40371;
  assign n35856 = ~n41408 & ~n40451;
  assign n35866 = ~n40377 & ~n36459;
  assign n40857 = ~n36914 & ~n35858;
  assign n35860 = ~n35859 & ~P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n35862 = ~n35861 | ~n35860;
  assign n35864 = ~n36193 | ~n35862;
  assign n35863 = n41149 ^ n40403;
  assign n40378 = n35864 ^ n35863;
  assign n35865 = ~n41531 & ~n40378;
  assign n35867 = ~n35866 & ~n35865;
  assign P3_U2818 = ~n35868 | ~n35867;
  assign n35872 = ~n43570 & ~n35869;
  assign n35871 = ~n35870 & ~n36135;
  assign n35874 = ~n35872 & ~n35871;
  assign n35873 = ~P1_PHYADDRPOINTER_REG_3__SCAN_IN | ~n43797;
  assign n35888 = ~n35874 | ~n35873;
  assign n35876 = ~n42405 | ~n35875;
  assign n35882 = ~n35877 & ~n35876;
  assign n35880 = ~n35878 | ~P1_REIP_REG_3__SCAN_IN;
  assign n35879 = ~n43796 | ~P1_EBX_REG_3__SCAN_IN;
  assign n35881 = ~n35880 | ~n35879;
  assign n35886 = ~n35882 & ~n35881;
  assign n35883 = ~n36143;
  assign n35885 = ~n35884 | ~n35883;
  assign n35890 = ~n35889 | ~n43559;
  assign P1_U2837 = ~n35891 | ~n35890;
  assign n35892 = ~n35893;
  assign n35898 = ~n40202 & ~n35892;
  assign n35895 = ~n41235 & ~n35893;
  assign n35894 = ~n40418 & ~n41540;
  assign n35896 = ~n35895 & ~n35894;
  assign n36342 = ~n40418 | ~n41535;
  assign n35897 = ~n35896 | ~n36342;
  assign n35899 = ~n35898 & ~n35897;
  assign n35901 = ~n42336 & ~n35899;
  assign n35900 = ~n42338 & ~n40418;
  assign n35903 = ~n35901 & ~n35900;
  assign P3_U2862 = ~n35903 | ~n35902;
  assign n35934 = ~n35905 & ~n35904;
  assign n35909 = ~n35907 | ~n35906;
  assign n35908 = ~n36154 | ~P3_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n35913 = ~n35909 | ~n35908;
  assign n35911 = ~n35930 | ~n35910;
  assign n35912 = ~n41401 & ~n35911;
  assign n35915 = ~n35913 & ~n35912;
  assign n35922 = ~n35915 | ~n35914;
  assign n35920 = ~n35917 & ~n35916;
  assign n35919 = ~n35944 | ~n35918;
  assign n35921 = ~n35920 & ~n35919;
  assign n35932 = ~n35922 & ~n35921;
  assign n35928 = ~n35924 & ~n35923;
  assign n35927 = ~n35926 | ~n35925;
  assign n35929 = ~n35928 & ~n35927;
  assign n35931 = ~n35930 | ~n35929;
  assign n35933 = ~n35932 | ~n35931;
  assign n35937 = ~n35934 & ~n35933;
  assign n35936 = ~P3_EBX_REG_2__SCAN_IN | ~n35935;
  assign P3_U2669 = ~n35937 | ~n35936;
  assign n35938 = ~n41518 | ~n41402;
  assign n41519 = ~n35939 | ~n35938;
  assign n35946 = ~n35945 | ~n36161;
  assign n35957 = ~n35946 | ~P3_EBX_REG_30__SCAN_IN;
  assign n35955 = ~n41518 & ~n35947;
  assign n35948 = ~P3_REIP_REG_30__SCAN_IN & ~n36158;
  assign n35953 = ~n35948 | ~P3_REIP_REG_29__SCAN_IN;
  assign n36157 = ~P3_REIP_REG_30__SCAN_IN | ~P3_REIP_REG_29__SCAN_IN;
  assign n35950 = ~n35949 & ~n36157;
  assign n36171 = ~n35951 & ~n35950;
  assign n35952 = ~n36171 | ~P3_REIP_REG_30__SCAN_IN;
  assign n35954 = ~n35953 | ~n35952;
  assign n35956 = ~n35955 & ~n35954;
  assign n42130 = ~P3_EBX_REG_30__SCAN_IN;
  assign n35961 = ~n35960 | ~n42130;
  assign P3_U2641 = ~n35962 | ~n35961;
  assign n35965 = ~n35964 & ~n35963;
  assign n35966 = ~n35965 & ~n33538;
  assign n35969 = ~n35966 | ~n36203;
  assign n35968 = ~n35967 | ~P2_EBX_REG_13__SCAN_IN;
  assign n35973 = n35969 & n35968;
  assign n40620 = ~n42140;
  assign n35972 = ~n40620 | ~n43525;
  assign P2_U2874 = ~n35973 | ~n35972;
  assign n36345 = ~n35974 ^ n35976;
  assign n35978 = ~n41397 & ~n36345;
  assign n36346 = ~n35976 ^ n35975;
  assign n35977 = ~n36914 & ~n36346;
  assign n35985 = ~n35978 & ~n35977;
  assign n41098 = ~n36660;
  assign n35983 = ~n36220 & ~n41098;
  assign n36353 = ~n40865 & ~n35979;
  assign n35981 = ~n36353;
  assign n35980 = ~n36871 | ~n36220;
  assign n35982 = ~n35981 | ~n35980;
  assign n35984 = ~n35983 & ~n35982;
  assign P3_U2829 = ~n35985 | ~n35984;
  assign n40280 = ~P3_REIP_REG_7__SCAN_IN | ~n41145;
  assign n35987 = ~n35986 | ~n36871;
  assign n35994 = ~n40280 | ~n35987;
  assign n40260 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n40263 = ~n35988 ^ n40260;
  assign n35992 = ~n36975 | ~n40263;
  assign n35990 = ~n22937 | ~n35989;
  assign n40261 = ~n35990 ^ P3_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n35991 = ~n40261 | ~n40743;
  assign n35993 = ~n35992 | ~n35991;
  assign n36000 = ~n35994 & ~n35993;
  assign n35996 = ~P3_PHYADDRPOINTER_REG_7__SCAN_IN | ~n36660;
  assign n36031 = ~n37089 & ~n35995;
  assign n36034 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN | ~n36031;
  assign n35998 = ~n35996 | ~n36034;
  assign n36066 = ~n35997 | ~n36031;
  assign n35999 = ~n35998 | ~n36066;
  assign P3_U2823 = ~n36000 | ~n35999;
  assign n36012 = ~n36002 & ~n36001;
  assign n36006 = ~n37638 | ~n40311;
  assign n36005 = ~n36004 | ~n36003;
  assign n36947 = ~n36006 | ~n36005;
  assign n36948 = ~n37131 | ~n36599;
  assign n38815 = ~n36599;
  assign n36946 = ~n23700 | ~n38815;
  assign n36007 = ~n36948 | ~n36946;
  assign n36008 = n36947 ^ n36007;
  assign n36010 = ~n36008 | ~n43693;
  assign n36009 = ~n41756 | ~n38815;
  assign n36014 = ~n36012 & ~n36011;
  assign n36013 = ~P2_EAX_REG_3__SCAN_IN | ~n43698;
  assign P2_U2916 = ~n36014 | ~n36013;
  assign n36016 = ~n39934 & ~n36269;
  assign n36015 = ~n24862 & ~n43734;
  assign n36018 = ~n36016 & ~n36015;
  assign n36017 = ~n40436 | ~n41688;
  assign P1_U2897 = ~n36018 | ~n36017;
  assign n40208 = ~P3_REIP_REG_6__SCAN_IN | ~n41145;
  assign n36030 = ~n40208;
  assign n40201 = ~n36020 ^ n36019;
  assign n36025 = ~n36914 & ~n40201;
  assign n36023 = ~n36022 & ~n36021;
  assign n40193 = ~n36023 ^ P3_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n36024 = ~n41397 & ~n40193;
  assign n36028 = ~n36025 & ~n36024;
  assign n36027 = ~n36026 | ~n36871;
  assign n36029 = ~n36028 | ~n36027;
  assign n36037 = ~n36030 & ~n36029;
  assign n36033 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN | ~n36660;
  assign n36032 = ~n36031;
  assign n36035 = ~n36033 | ~n36032;
  assign n36036 = ~n36035 | ~n36034;
  assign P3_U2824 = ~n36037 | ~n36036;
  assign n36044 = ~n41537 & ~n36040;
  assign n36056 = n36046 | n36045;
  assign n36051 = ~n36048 & ~n36047;
  assign n36050 = ~n36049 & ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n36053 = ~n36051 & ~n36050;
  assign n36054 = ~n36053 & ~n36052;
  assign n36060 = ~n36057 | ~n41326;
  assign n36059 = n42011 | n36058;
  assign n36062 = ~n36060 | ~n36059;
  assign n36065 = ~n36062 | ~n36061;
  assign n36064 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n36063;
  assign P3_U3285 = ~n36065 | ~n36064;
  assign n39638 = ~n41145 | ~P3_REIP_REG_8__SCAN_IN;
  assign n36074 = ~n39638;
  assign n36067 = ~P3_PHYADDRPOINTER_REG_8__SCAN_IN | ~n36660;
  assign n36069 = ~n36067 | ~n36066;
  assign n36072 = ~n36069 | ~n36068;
  assign n36071 = ~n36070 | ~n36871;
  assign n36073 = ~n36072 | ~n36071;
  assign n36085 = ~n36074 & ~n36073;
  assign n36076 = ~n36429 & ~n36075;
  assign n39616 = ~n40372 & ~n36076;
  assign n36083 = ~n41531 & ~n39616;
  assign n36081 = ~n39616 | ~n40744;
  assign n36079 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN & ~n36077;
  assign n39618 = ~n36079 & ~n36078;
  assign n36080 = ~n39618 | ~n40743;
  assign n36082 = ~n36081 | ~n36080;
  assign n36084 = ~n36083 & ~n36082;
  assign P3_U2822 = ~n36085 | ~n36084;
  assign n36098 = ~n43713 & ~n36110;
  assign n36087 = ~n36086;
  assign n36089 = ~n36088 & ~n36087;
  assign n36121 = ~n36092 | ~n36091;
  assign n36094 = ~n43358 & ~n36121;
  assign n36093 = ~n36109 & ~n43729;
  assign n36096 = ~n36094 & ~n36093;
  assign n36095 = ~P1_PHYADDRPOINTER_REG_5__SCAN_IN | ~n43709;
  assign n36124 = ~n43469 | ~P1_REIP_REG_5__SCAN_IN;
  assign P1_U2994 = ~n36099 | ~n36124;
  assign n36102 = ~n43570 & ~n36119;
  assign n36100 = ~P1_PHYADDRPOINTER_REG_5__SCAN_IN | ~n43797;
  assign n36101 = ~n36100 | ~n43033;
  assign n36106 = ~n36102 & ~n36101;
  assign n36105 = ~n36104 | ~n36103;
  assign n36108 = ~n41894 | ~n36107;
  assign n36114 = ~n36108 | ~P1_REIP_REG_5__SCAN_IN;
  assign n36112 = ~n36109 & ~n36143;
  assign n36111 = ~n36110 & ~n42175;
  assign n36113 = ~n36112 & ~n36111;
  assign n36117 = ~P1_EBX_REG_5__SCAN_IN | ~n43796;
  assign P1_U2835 = ~n36118 | ~n36117;
  assign n36127 = ~n43441 & ~n36119;
  assign n36123 = ~n36128 & ~n36120;
  assign n36130 = ~n36129 | ~n36128;
  assign P1_U3026 = ~n36131 | ~n36130;
  assign n36132 = ~n42185 & ~P1_REIP_REG_2__SCAN_IN;
  assign n36140 = ~n36132 | ~P1_REIP_REG_1__SCAN_IN;
  assign n36134 = ~n44022 | ~n43803;
  assign n36133 = ~n43797 | ~P1_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n36138 = ~n36134 | ~n36133;
  assign n36137 = ~n36136 & ~n36135;
  assign n36139 = ~n36138 & ~n36137;
  assign n36142 = ~n41894 | ~n36141;
  assign n36148 = ~n36142 | ~P1_REIP_REG_2__SCAN_IN;
  assign n36146 = ~n44020 & ~n36143;
  assign n36145 = ~n36144 & ~n42175;
  assign n36147 = ~n36146 & ~n36145;
  assign n36151 = ~P1_EBX_REG_2__SCAN_IN | ~n43796;
  assign P1_U2838 = ~n36152 | ~n36151;
  assign n36156 = ~n36153 | ~P3_EBX_REG_31__SCAN_IN;
  assign n36155 = ~n36154 | ~P3_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n36170 = ~n36156 | ~n36155;
  assign n36160 = ~n36158 & ~n36157;
  assign n36166 = ~n36161 & ~P3_EBX_REG_30__SCAN_IN;
  assign n36163 = ~n41519 | ~n36162;
  assign n36165 = ~n36164 & ~n36163;
  assign n36172 = ~P3_REIP_REG_31__SCAN_IN | ~n36171;
  assign P3_U2640 = ~n36173 | ~n36172;
  assign n36180 = ~n42135 | ~n36174;
  assign n36175 = ~P3_EBX_REG_18__SCAN_IN | ~n43930;
  assign n36178 = ~n36175 | ~n36177;
  assign P3_U2685 = ~n36180 | ~n36179;
  assign n36189 = ~n36181 & ~n36967;
  assign n40150 = ~n41145 | ~P3_REIP_REG_14__SCAN_IN;
  assign n36185 = ~n40150;
  assign n36183 = ~n36182 & ~P3_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n36214 = ~n41095 | ~n36222;
  assign n36184 = ~n36183 & ~n36214;
  assign n36187 = ~n36185 & ~n36184;
  assign n36186 = ~P3_PHYADDRPOINTER_REG_14__SCAN_IN | ~n37753;
  assign n36188 = ~n36187 | ~n36186;
  assign n36201 = ~n36189 & ~n36188;
  assign n40144 = ~n36227 ^ P3_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n36199 = ~n41408 & ~n40144;
  assign n36191 = ~n41149 | ~n36190;
  assign n36194 = ~n36192 | ~n36191;
  assign n40134 = ~n36195 ^ P3_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n36197 = ~n40134 | ~n40857;
  assign n40135 = ~n36230 ^ n40132;
  assign n36196 = ~n40135 | ~n40743;
  assign n36198 = ~n36197 | ~n36196;
  assign n36200 = ~n36199 & ~n36198;
  assign P3_U2816 = ~n36201 | ~n36200;
  assign n36204 = ~n36203 ^ n36202;
  assign n36208 = ~n36204 & ~n33538;
  assign n36207 = ~n42842 & ~n35967;
  assign n36210 = ~n36208 & ~n36207;
  assign n36209 = ~P2_EBX_REG_14__SCAN_IN | ~n35967;
  assign P2_U2873 = ~n36210 | ~n36209;
  assign n36226 = ~n41531 & ~n40229;
  assign n36213 = ~n41100 | ~n36212;
  assign n36215 = ~n36214 | ~n36213;
  assign n37696 = ~n37753 & ~n36215;
  assign n36219 = ~n37696 & ~n37694;
  assign n36217 = ~n36216 | ~n41400;
  assign n40235 = ~n41145 | ~P3_REIP_REG_15__SCAN_IN;
  assign n36218 = ~n36217 | ~n40235;
  assign n36224 = ~n36219 & ~n36218;
  assign n36221 = ~n41403 & ~n36220;
  assign n37698 = ~n36222 & ~n40872;
  assign n36223 = ~n37698 | ~n37694;
  assign n36225 = ~n36224 | ~n36223;
  assign n36236 = ~n36226 & ~n36225;
  assign n40339 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n36228 = ~n36227 | ~P3_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n40214 = ~n40339 | ~n36228;
  assign n36229 = ~n40214;
  assign n36234 = ~n36868 & ~n36229;
  assign n36231 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN | ~n36230;
  assign n40216 = ~n40339 | ~n36231;
  assign n36232 = ~n40216;
  assign n36233 = ~n36869 & ~n36232;
  assign n36235 = ~n36234 & ~n36233;
  assign P3_U2815 = ~n36236 | ~n36235;
  assign n36238 = ~n36237 | ~P3_EAX_REG_30__SCAN_IN;
  assign n36241 = ~n36238 & ~P3_EAX_REG_31__SCAN_IN;
  assign n41481 = ~BUF2_REG_31__SCAN_IN;
  assign n36240 = ~n41481 & ~n36239;
  assign n36247 = ~n36241 & ~n36240;
  assign n36244 = ~n36242 | ~n36280;
  assign n36245 = ~n36244 | ~n36281;
  assign n36246 = ~n36245 | ~P3_EAX_REG_31__SCAN_IN;
  assign P3_U2704 = ~n36247 | ~n36246;
  assign n36252 = ~n36248 & ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n36250 = ~n36249 | ~n43091;
  assign n36251 = ~n43523 | ~n36250;
  assign n36254 = ~n36252 & ~n36251;
  assign n36256 = ~n36254 | ~n36253;
  assign n36255 = ~n35967 | ~P2_EBX_REG_5__SCAN_IN;
  assign n36260 = n36256 & n36255;
  assign n40368 = n36258 ^ n36257;
  assign n36259 = ~n40368 | ~n43525;
  assign P2_U2882 = ~n36260 | ~n36259;
  assign n36262 = ~n43362 | ~n36992;
  assign n36261 = ~n43709 | ~P1_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n36268 = ~n36262 | ~n36261;
  assign n36266 = ~n36263;
  assign n36265 = ~n43707 | ~n36264;
  assign n36267 = ~n36266 | ~n36265;
  assign n36271 = ~n36268 & ~n36267;
  assign n36270 = ~n36993 | ~n43367;
  assign P1_U2992 = ~n36271 | ~n36270;
  assign n36275 = ~n37500;
  assign n36277 = ~n37242 & ~n44019;
  assign n36276 = ~n37246 & ~n43298;
  assign n36278 = ~P1_EBX_REG_8__SCAN_IN | ~n44023;
  assign P1_U2864 = ~n36279 | ~n36278;
  assign n36337 = ~n36281 & ~n36280;
  assign n36285 = BUF2_REG_30__SCAN_IN & n36282;
  assign n36284 = ~P3_EAX_REG_30__SCAN_IN & ~n36283;
  assign n36335 = ~n36285 & ~n36284;
  assign n36288 = ~n22917 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n36287 = ~n22920 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n36293 = ~n36288 | ~n36287;
  assign n36291 = ~n22902 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n36290 = ~n22913 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n36292 = ~n36291 | ~n36290;
  assign n36305 = ~n36293 & ~n36292;
  assign n36297 = ~n36294 | ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n36296 = ~n22914 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n36303 = ~n36297 | ~n36296;
  assign n36301 = ~n36298 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n36300 = ~n22923 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n36302 = ~n36301 | ~n36300;
  assign n36304 = ~n36303 & ~n36302;
  assign n36328 = ~n36305 | ~n36304;
  assign n36309 = ~n22919 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n36308 = ~n36307 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n36315 = ~n36309 | ~n36308;
  assign n36313 = ~n36310 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n36312 = ~n36311 | ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n36314 = ~n36313 | ~n36312;
  assign n36326 = ~n36315 & ~n36314;
  assign n36319 = ~n22903 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n36318 = ~n36317 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n36324 = ~n36319 | ~n36318;
  assign n36322 = ~n35392 | ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n36321 = ~n36320 | ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n36323 = ~n36322 | ~n36321;
  assign n36325 = ~n36324 & ~n36323;
  assign n36327 = ~n36326 | ~n36325;
  assign n36332 = ~n36328 & ~n36327;
  assign n36331 = ~n36330 & ~n36329;
  assign n42134 = ~n36332 ^ n36331;
  assign n36334 = ~n36333 | ~n42134;
  assign n36336 = ~n36335 | ~n36334;
  assign n36340 = ~n36337 & ~n36336;
  assign n36339 = ~BUF2_REG_14__SCAN_IN | ~n36338;
  assign P3_U2705 = ~n36340 | ~n36339;
  assign n36341 = ~n36352 | ~n41005;
  assign n36344 = ~n36341 & ~n36509;
  assign n36343 = ~n36352 & ~n36342;
  assign n36350 = ~n36344 & ~n36343;
  assign n36348 = ~n41235 & ~n36345;
  assign n36347 = ~n40202 & ~n36346;
  assign n36349 = ~n36348 & ~n36347;
  assign n36351 = ~n36350 | ~n36349;
  assign n36356 = ~n36351 | ~n41257;
  assign n36354 = ~n42338 & ~n36352;
  assign n36355 = ~n36354 & ~n36353;
  assign P3_U2861 = ~n36356 | ~n36355;
  assign n36361 = ~n36359 & ~n36360;
  assign n36362 = ~n31055 & ~n36361;
  assign n36372 = ~n36363 & ~n36362;
  assign n36367 = ~n36365 | ~n36364;
  assign n36368 = ~n36367 | ~n36366;
  assign n36369 = n36368 & P2_STATE2_REG_0__SCAN_IN;
  assign n36371 = ~n36370 | ~n36369;
  assign P2_U3177 = ~n36372 | ~n36371;
  assign n36394 = n42287 & n40602;
  assign n36378 = ~n39222 | ~n41718;
  assign n36379 = n36378 ^ n42438;
  assign n36389 = ~n36379 & ~n41919;
  assign n36383 = ~n40350 & ~n36380;
  assign n36381 = ~P2_EBX_REG_18__SCAN_IN | ~n41935;
  assign n36382 = ~n36381 | ~n40668;
  assign n36387 = ~n36383 & ~n36382;
  assign n36386 = ~n42285 | ~n41934;
  assign n36388 = ~n36387 | ~n36386;
  assign n36392 = ~n36389 & ~n36388;
  assign n36391 = ~P2_PHYADDRPOINTER_REG_18__SCAN_IN | ~n41921;
  assign n36397 = ~n42439;
  assign P2_U2837 = ~n36399 | ~n36398;
  assign n36406 = ~n42135 | ~n36400;
  assign n36402 = ~P3_EBX_REG_19__SCAN_IN | ~n43930;
  assign n36404 = ~n36402 | ~n36401;
  assign P3_U2684 = ~n36406 | ~n36405;
  assign n36408 = ~n39934 & ~n37242;
  assign n36407 = ~n44054 & ~n43734;
  assign n36410 = ~n36408 & ~n36407;
  assign n36409 = ~n40436 | ~n42043;
  assign P1_U2896 = ~n36410 | ~n36409;
  assign n36426 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN & ~n36459;
  assign n36414 = ~n36411 | ~n36871;
  assign n36413 = ~n36434 | ~n36412;
  assign n36419 = ~n36414 | ~n36413;
  assign n40463 = ~n41145 | ~P3_REIP_REG_9__SCAN_IN;
  assign n37748 = ~n40731;
  assign n36462 = ~n36415 | ~P3_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n36416 = ~n37748 | ~n36462;
  assign n36465 = ~n40734 | ~n36416;
  assign n36417 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN | ~n36465;
  assign n36418 = ~n40463 | ~n36417;
  assign n36424 = ~n36419 & ~n36418;
  assign n36421 = ~n40743 | ~n40371;
  assign n36420 = ~n40744 | ~n40451;
  assign n36422 = ~n36421 | ~n36420;
  assign n36423 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN | ~n36422;
  assign n36425 = ~n36424 | ~n36423;
  assign n36432 = ~n36426 & ~n36425;
  assign n36428 = ~n41147 & ~n39620;
  assign n36430 = n36444 & n36446;
  assign n40455 = ~n36430 ^ P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n36431 = ~n40857 | ~n40455;
  assign P3_U2821 = ~n36432 | ~n36431;
  assign n36435 = ~n36433 & ~P3_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n36443 = ~n36435 | ~n36434;
  assign n40987 = ~n41145 | ~P3_REIP_REG_11__SCAN_IN;
  assign n36437 = ~n36436 | ~n36871;
  assign n36441 = ~n40987 | ~n36437;
  assign n36463 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN & ~n37089;
  assign n36438 = ~n36463 & ~n36465;
  assign n36440 = ~n36439 & ~n36438;
  assign n36442 = ~n36441 & ~n36440;
  assign n36454 = ~n36443 | ~n36442;
  assign n36470 = ~n36444;
  assign n36445 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN & ~P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n36449 = ~n36470 | ~n36445;
  assign n36471 = ~n36446;
  assign n36448 = ~n36471 | ~n36447;
  assign n36450 = ~n36449 | ~n36448;
  assign n40979 = ~n40981 ^ n36450;
  assign n36452 = ~n40857 | ~n40979;
  assign n37086 = ~n36459 & ~n40959;
  assign n36451 = ~n37086 | ~n40981;
  assign n36453 = ~n36452 | ~n36451;
  assign n36458 = ~n36454 & ~n36453;
  assign n36456 = ~n40743 | ~n40500;
  assign n36455 = ~n40744 | ~n40503;
  assign n36457 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN | ~n36479;
  assign P3_U2819 = ~n36458 | ~n36457;
  assign n40513 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN | ~n27697;
  assign n36478 = ~n36459 & ~n40513;
  assign n40519 = ~n41145 | ~P3_REIP_REG_10__SCAN_IN;
  assign n36461 = ~n36460 | ~n36871;
  assign n36469 = ~n40519 | ~n36461;
  assign n36464 = ~n36462;
  assign n36467 = ~n36464 | ~n36463;
  assign n36466 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN | ~n36465;
  assign n36468 = ~n36467 | ~n36466;
  assign n36476 = ~n36469 & ~n36468;
  assign n36473 = ~n36470 | ~n27696;
  assign n36472 = ~n36471 | ~P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n36474 = ~n36473 | ~n36472;
  assign n40510 = n36474 ^ P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n36475 = ~n40857 | ~n40510;
  assign n36477 = ~n36476 | ~n36475;
  assign n36481 = ~n36478 & ~n36477;
  assign n36480 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN | ~n36479;
  assign P3_U2820 = ~n36481 | ~n36480;
  assign n36484 = ~n43911 & ~n38829;
  assign n36604 = ~n43880 | ~P2_REIP_REG_3__SCAN_IN;
  assign n36482 = ~n43917 | ~P2_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n36483 = ~n36604 | ~n36482;
  assign n36496 = ~n36484 & ~n36483;
  assign n36494 = ~n36612 & ~n43924;
  assign n36851 = ~n36490;
  assign n36491 = ~n43813 | ~n36607;
  assign n36495 = ~n36494 & ~n36493;
  assign P2_U3011 = ~n36496 | ~n36495;
  assign n36499 = ~n36532 & ~n36497;
  assign n36498 = ~n37638 & ~n36533;
  assign n36505 = ~n36499 & ~n36498;
  assign n36537 = ~n31055 & ~n36500;
  assign n37315 = n37285 ^ n36501;
  assign n36503 = ~n37315 | ~n41718;
  assign n36502 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN | ~n41204;
  assign n36536 = ~n36503 | ~n36502;
  assign n36504 = ~n36537 | ~n36536;
  assign n36506 = ~n36505 | ~n36504;
  assign n36508 = ~n36542 | ~n36506;
  assign n36507 = ~n36543 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign P2_U3599 = ~n36508 | ~n36507;
  assign n36510 = ~n39404 | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n36514 = ~n36526 | ~n36510;
  assign n40445 = ~n42322;
  assign n40247 = ~n40418 | ~n42320;
  assign n36511 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN | ~n40247;
  assign n36512 = ~n40445 | ~n36511;
  assign n36513 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN | ~n36512;
  assign n36524 = ~n36514 | ~n36513;
  assign n40384 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~n40168;
  assign n36522 = ~n40384 & ~n40442;
  assign n36518 = ~n41235 & ~n36515;
  assign n36517 = ~n40202 & ~n36516;
  assign n36520 = ~n36518 & ~n36517;
  assign n38598 = ~n40422 | ~n36519;
  assign n36521 = ~n36520 | ~n38598;
  assign n36523 = ~n36522 & ~n36521;
  assign n36525 = ~n36524 | ~n36523;
  assign n36530 = ~n36525 | ~n41257;
  assign n36528 = ~n42338 & ~n36526;
  assign n36529 = ~n36528 & ~n36527;
  assign P3_U2860 = ~n36530 | ~n36529;
  assign n36535 = ~n36532 & ~n36531;
  assign n36534 = ~n37945 & ~n36533;
  assign n36540 = ~n36535 & ~n36534;
  assign n36538 = ~n36536;
  assign n36539 = ~n36538 | ~n36537;
  assign n36541 = ~n36540 | ~n36539;
  assign n36545 = ~n36542 | ~n36541;
  assign n36544 = ~n36543 | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign P2_U3600 = ~n36545 | ~n36544;
  assign n36551 = P2_EBX_REG_15__SCAN_IN & n35967;
  assign n36548 = ~n36547 & ~n36546;
  assign n36549 = ~n36548 & ~n33538;
  assign n36550 = n36549 & n37120;
  assign n36555 = ~n36551 & ~n36550;
  assign n36554 = ~n42424 | ~n43525;
  assign P2_U2872 = ~n36555 | ~n36554;
  assign n36577 = ~n37131 | ~n36556;
  assign n39021 = ~n36577 & ~n38279;
  assign n36802 = ~n36557 & ~n43915;
  assign n36803 = ~n36558 & ~n43915;
  assign n36564 = ~n38221 & ~n40906;
  assign n36778 = ~n38334 & ~n39522;
  assign n37132 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n37610 = ~n36562 & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n36563 = ~n39230 & ~n37596;
  assign n36585 = ~n36564 & ~n36563;
  assign n38235 = ~n37596;
  assign n36566 = ~n36569 & ~n38235;
  assign n36567 = ~n36566 & ~n39511;
  assign n36583 = ~n40908 & ~n37597;
  assign n36570 = ~n36569 | ~n39522;
  assign n36571 = ~n36570 | ~n39524;
  assign n36572 = ~n38235 & ~n36571;
  assign n36576 = ~n38334 & ~n36572;
  assign n36573 = ~n37610;
  assign n36581 = ~P2_INSTQUEUE_REG_1__2__SCAN_IN | ~n37604;
  assign n39233 = ~n36579 | ~n36578;
  assign n36580 = ~n37839 | ~n39233;
  assign n36582 = ~n36581 | ~n36580;
  assign n36584 = ~n36583 & ~n36582;
  assign P2_U3058 = ~n36585 | ~n36584;
  assign n36589 = ~n38221 & ~n41290;
  assign n39601 = ~n23415 | ~n36778;
  assign n36588 = ~n39601 & ~n37596;
  assign n36598 = ~n36589 & ~n36588;
  assign n36596 = ~n41289 & ~n37597;
  assign n36594 = ~P2_INSTQUEUE_REG_1__7__SCAN_IN | ~n37604;
  assign n39606 = ~n36592 | ~n36591;
  assign n36593 = ~n37839 | ~n39606;
  assign n36595 = ~n36594 | ~n36593;
  assign n36597 = ~n36596 & ~n36595;
  assign P2_U3063 = ~n36598 | ~n36597;
  assign n36611 = ~n43877 & ~n36599;
  assign n36603 = ~n42699 & ~n36600;
  assign n36602 = ~n43159 & ~n36601;
  assign n36841 = ~n36603 & ~n36602;
  assign n36606 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN & ~n36841;
  assign n36605 = ~n36604;
  assign n36609 = ~n36606 & ~n36605;
  assign n36608 = ~n43767 | ~n36607;
  assign n36610 = ~n36609 | ~n36608;
  assign n36619 = ~n36611 & ~n36610;
  assign n36617 = ~n36612 & ~n43893;
  assign n36614 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN | ~n36846;
  assign n36618 = ~n36617 & ~n36616;
  assign P2_U3043 = ~n36619 | ~n36618;
  assign n36623 = ~n38221 & ~n39549;
  assign n36622 = ~n39251 & ~n37596;
  assign n36631 = ~n36623 & ~n36622;
  assign n36629 = ~n39540 & ~n37597;
  assign n36627 = ~P2_INSTQUEUE_REG_1__1__SCAN_IN | ~n37604;
  assign n39542 = ~n36625 | ~n36624;
  assign n36626 = ~n37839 | ~n39542;
  assign n36628 = ~n36627 | ~n36626;
  assign n36630 = ~n36629 & ~n36628;
  assign P2_U3057 = ~n36631 | ~n36630;
  assign n39244 = ~n36633 | ~n36632;
  assign n36647 = ~n39535 & ~n38305;
  assign n37944 = ~n36635 & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n36651 = ~n36796;
  assign n36636 = ~n36648 & ~n36651;
  assign n36639 = ~n36636 & ~n39511;
  assign n36637 = ~n37944;
  assign n36638 = ~n36637 & ~n39524;
  assign n36641 = ~n39515 & ~n36793;
  assign n36640 = ~n39241 & ~n36796;
  assign n36645 = ~n36641 & ~n36640;
  assign n38773 = ~n36652 & ~n38279;
  assign n39517 = ~n36643 | ~n36642;
  assign n36644 = ~n38773 | ~n39517;
  assign n36646 = ~n36645 | ~n36644;
  assign n36658 = ~n36647 & ~n36646;
  assign n36649 = ~n36648 | ~n39522;
  assign n36650 = ~n36649 | ~n39524;
  assign n36655 = ~n36651 & ~n36650;
  assign n36657 = ~P2_INSTQUEUE_REG_13__0__SCAN_IN | ~n36801;
  assign P2_U3152 = ~n36658 | ~n36657;
  assign n36962 = ~n36659 | ~n40734;
  assign n36917 = ~n36660 | ~n36962;
  assign n36662 = ~n37089 & ~n36661;
  assign n36663 = ~P3_PHYADDRPOINTER_REG_3__SCAN_IN & ~n36662;
  assign n36674 = ~n36917 & ~n36663;
  assign n38724 = ~n36665 ^ n36664;
  assign n36669 = ~n36914 & ~n38724;
  assign n38723 = ~n36667 ^ n36666;
  assign n36668 = ~n41397 & ~n38723;
  assign n36672 = ~n36669 & ~n36668;
  assign n36671 = n36967 | n36670;
  assign n36675 = ~n36674 & ~n36673;
  assign n38735 = ~n41145 | ~P3_REIP_REG_3__SCAN_IN;
  assign P3_U2827 = ~n36675 | ~n38735;
  assign n39153 = ~n41873 | ~n36778;
  assign n36681 = ~n39153 & ~n37596;
  assign n39156 = ~n36677 | ~n36676;
  assign n36679 = ~n37839 | ~n39156;
  assign n36678 = ~P2_INSTQUEUE_REG_1__5__SCAN_IN | ~n37604;
  assign n36687 = ~n36681 & ~n36680;
  assign n36685 = ~n38221 & ~n40883;
  assign n36684 = ~n40882 & ~n37597;
  assign n36686 = ~n36685 & ~n36684;
  assign P2_U3061 = ~n36687 | ~n36686;
  assign n36690 = ~n41301 & ~n36793;
  assign n36689 = ~n39200 & ~n36796;
  assign n36700 = ~n36690 & ~n36689;
  assign n39201 = ~n36692 | ~n36691;
  assign n36698 = ~n38305 & ~n41295;
  assign n36696 = ~P2_INSTQUEUE_REG_13__6__SCAN_IN | ~n36801;
  assign n36695 = ~n38773 | ~n38696;
  assign n36699 = ~n36698 & ~n36697;
  assign P2_U3158 = ~n36700 | ~n36699;
  assign n36702 = ~n40882 & ~n36793;
  assign n36701 = ~n39153 & ~n36796;
  assign n36708 = ~n36702 & ~n36701;
  assign n36706 = ~n38305 & ~n40881;
  assign n36704 = ~P2_INSTQUEUE_REG_13__5__SCAN_IN | ~n36801;
  assign n36703 = ~n38773 | ~n38687;
  assign n36707 = ~n36706 & ~n36705;
  assign P2_U3157 = ~n36708 | ~n36707;
  assign n36710 = ~n41289 & ~n36793;
  assign n36709 = ~n39601 & ~n36796;
  assign n36716 = ~n36710 & ~n36709;
  assign n36714 = ~n38305 & ~n41283;
  assign n36712 = ~P2_INSTQUEUE_REG_13__7__SCAN_IN | ~n36801;
  assign n36711 = ~n38773 | ~n37808;
  assign n36715 = ~n36714 & ~n36713;
  assign P2_U3159 = ~n36716 | ~n36715;
  assign n36718 = ~n39540 & ~n36793;
  assign n36717 = ~n39251 & ~n36796;
  assign n36724 = ~n36718 & ~n36717;
  assign n36722 = ~n38305 & ~n38703;
  assign n36720 = ~P2_INSTQUEUE_REG_13__1__SCAN_IN | ~n36801;
  assign n36719 = ~n38773 | ~n38706;
  assign n36721 = ~n36720 | ~n36719;
  assign n36723 = ~n36722 & ~n36721;
  assign P2_U3153 = ~n36724 | ~n36723;
  assign n36726 = ~n40908 & ~n36793;
  assign n36725 = ~n39230 & ~n36796;
  assign n36732 = ~n36726 & ~n36725;
  assign n36730 = ~n38305 & ~n40907;
  assign n36728 = ~P2_INSTQUEUE_REG_13__2__SCAN_IN | ~n36801;
  assign n36727 = ~n38773 | ~n38715;
  assign n36731 = ~n36730 & ~n36729;
  assign P2_U3154 = ~n36732 | ~n36731;
  assign n36743 = ~n41295 & ~n39187;
  assign n36733 = ~n36746 | ~n39522;
  assign n36734 = ~n36733 | ~n39524;
  assign n36735 = ~n37542 & ~n36734;
  assign n36739 = ~n36735 & ~n38334;
  assign n36741 = ~P2_INSTQUEUE_REG_7__6__SCAN_IN | ~n37547;
  assign n36740 = ~n41296 | ~n37542;
  assign n36742 = ~n36741 | ~n36740;
  assign n36753 = ~n36743 & ~n36742;
  assign n36751 = ~n37854 & ~n41302;
  assign n36747 = ~n36746 & ~n37542;
  assign n36748 = ~n36747 & ~n39511;
  assign n36750 = ~n41301 & ~n37539;
  assign n36752 = ~n36751 & ~n36750;
  assign P2_U3110 = ~n36753 | ~n36752;
  assign n36757 = ~n40883 & ~n37854;
  assign n36755 = ~P2_INSTQUEUE_REG_7__5__SCAN_IN | ~n37547;
  assign n40886 = ~n39153;
  assign n36754 = ~n40886 | ~n37542;
  assign n36756 = ~n36755 | ~n36754;
  assign n36761 = ~n36757 & ~n36756;
  assign n36759 = ~n39187 & ~n40881;
  assign n36758 = ~n40882 & ~n37539;
  assign n36760 = ~n36759 & ~n36758;
  assign P2_U3109 = ~n36761 | ~n36760;
  assign n36765 = ~n41290 & ~n37854;
  assign n36763 = ~P2_INSTQUEUE_REG_7__7__SCAN_IN | ~n37547;
  assign n36762 = ~n41284 | ~n37542;
  assign n36764 = ~n36763 | ~n36762;
  assign n36769 = ~n36765 & ~n36764;
  assign n36767 = ~n39187 & ~n41283;
  assign n36766 = ~n41289 & ~n37539;
  assign n36768 = ~n36767 & ~n36766;
  assign P2_U3111 = ~n36769 | ~n36768;
  assign n36773 = ~n39549 & ~n37854;
  assign n36771 = ~P2_INSTQUEUE_REG_7__1__SCAN_IN | ~n37547;
  assign n36770 = ~n39541 | ~n37542;
  assign n36772 = ~n36771 | ~n36770;
  assign n36777 = ~n36773 & ~n36772;
  assign n36775 = ~n39187 & ~n38703;
  assign n36774 = ~n39540 & ~n37539;
  assign n36776 = ~n36775 & ~n36774;
  assign P2_U3105 = ~n36777 | ~n36776;
  assign n36781 = ~n41317 & ~n36793;
  assign n39268 = ~n36779 | ~n36778;
  assign n36780 = ~n39268 & ~n36796;
  assign n36791 = ~n36781 & ~n36780;
  assign n39271 = ~n36783 | ~n36782;
  assign n36789 = ~n38305 & ~n41308;
  assign n36787 = ~P2_INSTQUEUE_REG_13__4__SCAN_IN | ~n36801;
  assign n38678 = ~n36785 | ~n36784;
  assign n36786 = ~n38773 | ~n38678;
  assign n36790 = ~n36789 & ~n36788;
  assign P2_U3156 = ~n36791 | ~n36790;
  assign n36798 = ~n40896 & ~n36793;
  assign n36797 = ~n39280 & ~n36796;
  assign n36811 = ~n36798 & ~n36797;
  assign n39285 = ~n36800 | ~n36799;
  assign n36809 = ~n38305 & ~n40895;
  assign n36807 = ~P2_INSTQUEUE_REG_13__3__SCAN_IN | ~n36801;
  assign n38669 = ~n36805 | ~n36804;
  assign n36806 = ~n38773 | ~n38669;
  assign n36810 = ~n36809 & ~n36808;
  assign P2_U3155 = ~n36811 | ~n36810;
  assign n36815 = ~n40894 & ~n37854;
  assign n36813 = ~P2_INSTQUEUE_REG_7__3__SCAN_IN | ~n37547;
  assign n36812 = ~n40899 | ~n37542;
  assign n36814 = ~n36813 | ~n36812;
  assign n36819 = ~n36815 & ~n36814;
  assign n36817 = ~n39187 & ~n40895;
  assign n36816 = ~n40896 & ~n37539;
  assign n36818 = ~n36817 & ~n36816;
  assign P2_U3107 = ~n36819 | ~n36818;
  assign n36821 = ~n38221 & ~n40894;
  assign n36820 = ~n39280 & ~n37596;
  assign n36827 = ~n36821 & ~n36820;
  assign n36825 = ~n40896 & ~n37597;
  assign n36823 = ~P2_INSTQUEUE_REG_1__3__SCAN_IN | ~n37604;
  assign n36822 = ~n37839 | ~n39285;
  assign n36824 = ~n36823 | ~n36822;
  assign n36826 = ~n36825 & ~n36824;
  assign P2_U3059 = ~n36827 | ~n36826;
  assign n40354 = ~n36829 ^ n36828;
  assign n36837 = ~n40354 & ~n43695;
  assign n40559 = ~n36831 ^ n36830;
  assign n36832 = ~n40559;
  assign n36953 = ~n36832 | ~n40580;
  assign n36833 = ~n36953 | ~n40354;
  assign n36835 = ~n36833 | ~n43693;
  assign n36834 = ~n36955 | ~n39675;
  assign n36836 = ~n36835 | ~n36834;
  assign n36839 = ~n36837 & ~n36836;
  assign n36838 = ~P2_EAX_REG_5__SCAN_IN | ~n43698;
  assign P2_U2914 = ~n36839 | ~n36838;
  assign n36843 = ~n43767 | ~n40565;
  assign n39658 = ~n36841 & ~n36840;
  assign n36842 = ~n39658 | ~n39656;
  assign n36850 = ~n36843 | ~n36842;
  assign n36845 = ~n43877 & ~n40559;
  assign n37558 = ~n43880 | ~P2_REIP_REG_4__SCAN_IN;
  assign n36844 = ~n37558;
  assign n36848 = ~n36845 & ~n36844;
  assign n36847 = ~P2_INSTADDRPOINTER_REG_4__SCAN_IN | ~n36846;
  assign n36849 = ~n36848 | ~n36847;
  assign n36865 = ~n36850 & ~n36849;
  assign n36856 = ~n36852 & ~n36851;
  assign n36855 = ~n36854 | ~n36853;
  assign n36858 = n36856 | n36855;
  assign n36863 = ~n37557 & ~n43755;
  assign n36864 = ~n36863 & ~n36862;
  assign P2_U3042 = ~n36865 | ~n36864;
  assign n37706 = ~n36867 & ~n36866;
  assign n36870 = ~n39450 & ~n37706;
  assign n36884 = ~n37021 & ~n39440;
  assign n39392 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN | ~n39440;
  assign n36881 = ~n37706 & ~n39392;
  assign n36879 = ~n36872 | ~n36871;
  assign n36875 = ~n36873 | ~n41095;
  assign n36877 = ~n36875 | ~n36874;
  assign n36876 = ~n37748 | ~n37016;
  assign n37012 = ~n40734 | ~n36876;
  assign n36878 = ~n36877 | ~n37012;
  assign n36880 = ~n36879 | ~n36878;
  assign n36882 = ~n36881 & ~n36880;
  assign n39418 = ~n41145 | ~P3_REIP_REG_17__SCAN_IN;
  assign n36883 = ~n36882 | ~n39418;
  assign n36888 = ~n36884 & ~n36883;
  assign n36886 = n36885 | n39440;
  assign P3_U2813 = ~n36888 | ~n36887;
  assign n36899 = n39557 | P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n36892 = ~n36891 | ~n38648;
  assign n36897 = ~n36893 | ~n36892;
  assign n36896 = ~n36895 & ~n36894;
  assign n39559 = ~n36897 & ~n36896;
  assign n36898 = ~n39559 | ~P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n36912 = ~n36899 | ~n36898;
  assign n36903 = ~n37220;
  assign n36902 = ~n36901 | ~n36900;
  assign n36910 = ~n43441 & ~n37550;
  assign n37496 = ~n43033 & ~n37508;
  assign n36907 = ~n37496;
  assign P1_U3022 = ~n36912 | ~n36911;
  assign n40183 = ~n36913 ^ P3_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n36926 = ~n36914 & ~n40183;
  assign n36923 = ~n36967 & ~n36915;
  assign n36916 = ~n37748 | ~n36963;
  assign n36964 = ~n36917 | ~n36916;
  assign n36919 = ~n36964 & ~n40731;
  assign n36921 = ~n36919 | ~n36918;
  assign n36920 = ~n36964 | ~P3_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n36922 = ~n36921 | ~n36920;
  assign n36924 = ~n36923 & ~n36922;
  assign n40189 = ~P3_REIP_REG_5__SCAN_IN | ~n41145;
  assign n36925 = ~n36924 | ~n40189;
  assign n36929 = ~n36926 & ~n36925;
  assign n40180 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN ^ n36927;
  assign n36928 = ~n40180 | ~n40743;
  assign P3_U2825 = ~n36929 | ~n36928;
  assign n36933 = ~n41308 & ~n39187;
  assign n36931 = ~P2_INSTQUEUE_REG_7__4__SCAN_IN | ~n37547;
  assign n41311 = ~n39268;
  assign n36930 = ~n41311 | ~n37542;
  assign n36932 = ~n36931 | ~n36930;
  assign n36937 = ~n36933 & ~n36932;
  assign n36935 = ~n37854 & ~n41318;
  assign n36934 = ~n41317 & ~n37539;
  assign n36936 = ~n36935 & ~n36934;
  assign P2_U3108 = ~n36937 | ~n36936;
  assign n36941 = ~n39241 & ~n37596;
  assign n36939 = ~n37839 | ~n39244;
  assign n36938 = ~P2_INSTQUEUE_REG_1__0__SCAN_IN | ~n37604;
  assign n36945 = ~n36941 & ~n36940;
  assign n36943 = ~n38221 & ~n39240;
  assign n36942 = ~n39515 & ~n37597;
  assign n36944 = ~n36943 & ~n36942;
  assign P2_U3056 = ~n36945 | ~n36944;
  assign n36959 = ~n40559 & ~n43695;
  assign n36949 = ~n36947 | ~n36946;
  assign n36951 = ~n36949 | ~n36948;
  assign n36950 = ~n40580 & ~n36832;
  assign n36952 = ~n36951 | ~n36950;
  assign n36954 = n36952 & n43693;
  assign n36956 = ~n36955 | ~n38972;
  assign n36961 = ~n36959 & ~n36958;
  assign n36960 = ~P2_EAX_REG_4__SCAN_IN | ~n43698;
  assign P2_U2915 = ~n36961 | ~n36960;
  assign n36965 = ~n36963 | ~n36962;
  assign n36980 = ~n36965 | ~n36964;
  assign n38590 = ~n40865 & ~n36966;
  assign n36972 = ~n36968 & ~n36967;
  assign n38593 = ~n36970 ^ n36969;
  assign n36971 = ~n41397 & ~n38593;
  assign n36977 = ~n36972 & ~n36971;
  assign n38592 = n36974 ^ n36973;
  assign n36976 = ~n36975 | ~n38592;
  assign n36979 = ~n38590 & ~n36978;
  assign P3_U2826 = ~n36980 | ~n36979;
  assign n36989 = ~n36981 & ~n43570;
  assign n37238 = ~n42405 | ~n37235;
  assign n36985 = ~n37238 & ~n36982;
  assign n36983 = ~P1_PHYADDRPOINTER_REG_7__SCAN_IN | ~n43797;
  assign n36984 = ~n36983 | ~n43033;
  assign n36987 = ~n36985 & ~n36984;
  assign n36986 = ~P1_EBX_REG_7__SCAN_IN | ~n43796;
  assign n36988 = ~n36987 | ~n36986;
  assign n36999 = ~n36989 & ~n36988;
  assign n36997 = ~n36991 & ~n36990;
  assign n36995 = ~n36992 | ~n43559;
  assign n36994 = ~n36993 | ~n41453;
  assign n36996 = ~n36995 | ~n36994;
  assign n36998 = ~n36997 & ~n36996;
  assign P1_U2833 = ~n36999 | ~n36998;
  assign n37005 = n43709 & P1_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n37008 = ~n43713 & ~n37243;
  assign P1_U2991 = n37009 | n37008;
  assign n37020 = ~n37010 & ~n41520;
  assign n37013 = n41100 & n37011;
  assign n38033 = ~n37013 & ~n37012;
  assign n37015 = ~n38031 & ~n38033;
  assign n39459 = ~n41145 | ~P3_REIP_REG_18__SCAN_IN;
  assign n37014 = ~n39459;
  assign n37018 = ~n37015 & ~n37014;
  assign n38035 = ~n37016 & ~n40872;
  assign n37017 = ~n38035 | ~n38031;
  assign n37019 = ~n37018 | ~n37017;
  assign n37029 = ~n37020 & ~n37019;
  assign n37027 = ~n40421 & ~n37021;
  assign n37022 = ~n38143 | ~n37568;
  assign n38142 = ~n37706 & ~n37023;
  assign P3_U2812 = ~n37029 | ~n37028;
  assign n38208 = ~n37045 | ~n38279;
  assign n37032 = ~n38208 & ~n39535;
  assign n37030 = ~n37635 | ~n37634;
  assign n37076 = ~n37851 | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n37031 = ~n39241 & ~n37076;
  assign n37051 = ~n37032 & ~n37031;
  assign n37034 = ~n37851;
  assign n37035 = ~n37039 & ~n38294;
  assign n37036 = ~n37035 & ~n39511;
  assign n37049 = ~n39515 & ~n37416;
  assign n37040 = ~n37039 | ~n39522;
  assign n37041 = ~n37040 | ~n39524;
  assign n37042 = ~n38294 & ~n37041;
  assign n37047 = ~P2_INSTQUEUE_REG_9__0__SCAN_IN | ~n37423;
  assign n37046 = ~n39286 | ~n39517;
  assign n37050 = ~n37049 & ~n37048;
  assign P2_U3120 = ~n37051 | ~n37050;
  assign n37053 = ~n38208 & ~n41295;
  assign n37052 = ~n39200 & ~n37076;
  assign n37059 = ~n37053 & ~n37052;
  assign n37057 = ~n41301 & ~n37416;
  assign n37055 = ~P2_INSTQUEUE_REG_9__6__SCAN_IN | ~n37423;
  assign n37054 = ~n39286 | ~n38696;
  assign n37058 = ~n37057 & ~n37056;
  assign P2_U3126 = ~n37059 | ~n37058;
  assign n37061 = ~n38208 & ~n41308;
  assign n37060 = ~n39268 & ~n37076;
  assign n37067 = ~n37061 & ~n37060;
  assign n37065 = ~n41317 & ~n37416;
  assign n37063 = ~P2_INSTQUEUE_REG_9__4__SCAN_IN | ~n37423;
  assign n37062 = ~n39286 | ~n38678;
  assign n37066 = ~n37065 & ~n37064;
  assign P2_U3124 = ~n37067 | ~n37066;
  assign n37069 = ~n38208 & ~n40881;
  assign n37068 = ~n39153 & ~n37076;
  assign n37075 = ~n37069 & ~n37068;
  assign n37073 = ~n40882 & ~n37416;
  assign n37071 = ~P2_INSTQUEUE_REG_9__5__SCAN_IN | ~n37423;
  assign n37070 = ~n39286 | ~n38687;
  assign n37074 = ~n37073 & ~n37072;
  assign P2_U3125 = ~n37075 | ~n37074;
  assign n37078 = ~n38208 & ~n40895;
  assign n37077 = ~n39280 & ~n37076;
  assign n37084 = ~n37078 & ~n37077;
  assign n37082 = ~n40896 & ~n37416;
  assign n37080 = ~P2_INSTQUEUE_REG_9__3__SCAN_IN | ~n37423;
  assign n37079 = ~n39286 | ~n38669;
  assign n37083 = ~n37082 & ~n37081;
  assign P2_U3123 = ~n37084 | ~n37083;
  assign n40962 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n37105 = ~n37085 & ~n40962;
  assign n37087 = ~n40969 & ~P3_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n37103 = ~n37087 | ~n37086;
  assign n40956 = ~n40865 & ~n37088;
  assign n38155 = ~n37089 | ~n41403;
  assign n37091 = ~n37090 | ~n38155;
  assign n37093 = ~n37092 | ~n37091;
  assign n37100 = ~n37093 | ~P3_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n37095 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN | ~n37094;
  assign n37098 = ~n37095 & ~P3_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n37097 = ~n37096 & ~n41520;
  assign n37099 = ~n37098 & ~n37097;
  assign n37101 = ~n37100 | ~n37099;
  assign n37102 = ~n40956 & ~n37101;
  assign n37104 = ~n37103 | ~n37102;
  assign n37111 = ~n37105 & ~n37104;
  assign n37109 = ~n37106;
  assign n37108 = ~n37107 | ~P3_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n37110 = ~n40857 | ~n40958;
  assign P3_U2817 = ~n37111 | ~n37110;
  assign n37114 = ~P2_EAX_REG_16__SCAN_IN | ~n43698;
  assign n37113 = ~n42804 | ~n37112;
  assign n37118 = ~n37114 | ~n37113;
  assign n37116 = ~BUF2_REG_16__SCAN_IN | ~n43689;
  assign n37115 = ~BUF1_REG_16__SCAN_IN | ~n43690;
  assign n37117 = ~n37116 | ~n37115;
  assign n37129 = ~n37118 & ~n37117;
  assign n37122 = ~n37442;
  assign n37127 = ~n37352 & ~n41754;
  assign n37125 = n37124 | n37123;
  assign n37126 = ~n42633 & ~n43695;
  assign P2_U2903 = ~n37129 | ~n37128;
  assign n39193 = ~n37147 & ~n38279;
  assign n37134 = ~n39110 & ~n39240;
  assign n39123 = ~n38316 & ~n39114;
  assign n37202 = ~n39123;
  assign n37133 = ~n39241 & ~n37202;
  assign n37153 = ~n37134 & ~n37133;
  assign n37135 = n38321 | n37147;
  assign n37136 = ~n37139 & ~n39123;
  assign n37137 = ~n37136 & ~n39511;
  assign n37151 = ~n39515 & ~n37205;
  assign n37140 = ~n37139 | ~n39522;
  assign n37141 = ~n37140 | ~n39524;
  assign n37142 = ~n39123 & ~n37141;
  assign n37146 = ~n38334 & ~n37142;
  assign n37149 = ~P2_INSTQUEUE_REG_5__0__SCAN_IN | ~n37206;
  assign n37148 = ~n38319 | ~n39244;
  assign P2_U3088 = ~n37153 | ~n37152;
  assign n37155 = ~n39602 & ~n41308;
  assign n37154 = ~n39268 & ~n37202;
  assign n37161 = ~n37155 & ~n37154;
  assign n37159 = ~n41317 & ~n37205;
  assign n37157 = ~P2_INSTQUEUE_REG_5__4__SCAN_IN | ~n37206;
  assign n37156 = ~n39193 | ~n38678;
  assign P2_U3092 = ~n37161 | ~n37160;
  assign n37163 = ~n39110 & ~n41302;
  assign n37162 = ~n39200 & ~n37202;
  assign n37169 = ~n37163 & ~n37162;
  assign n37167 = ~n41301 & ~n37205;
  assign n37165 = ~P2_INSTQUEUE_REG_5__6__SCAN_IN | ~n37206;
  assign n37164 = ~n38319 | ~n39201;
  assign P2_U3094 = ~n37169 | ~n37168;
  assign n37171 = ~n39602 & ~n40895;
  assign n37170 = ~n39280 & ~n37202;
  assign n37177 = ~n37171 & ~n37170;
  assign n37175 = ~n40896 & ~n37205;
  assign n37173 = ~P2_INSTQUEUE_REG_5__3__SCAN_IN | ~n37206;
  assign n37172 = ~n39193 | ~n38669;
  assign P2_U3091 = ~n37177 | ~n37176;
  assign n37179 = ~n39110 & ~n40883;
  assign n37178 = ~n39153 & ~n37202;
  assign n37185 = ~n37179 & ~n37178;
  assign n37183 = ~n40882 & ~n37205;
  assign n37181 = ~P2_INSTQUEUE_REG_5__5__SCAN_IN | ~n37206;
  assign n37180 = ~n38319 | ~n39156;
  assign P2_U3093 = ~n37185 | ~n37184;
  assign n37187 = ~n39110 & ~n41290;
  assign n37186 = ~n39601 & ~n37202;
  assign n37193 = ~n37187 & ~n37186;
  assign n37191 = ~n41289 & ~n37205;
  assign n37189 = ~P2_INSTQUEUE_REG_5__7__SCAN_IN | ~n37206;
  assign n37188 = ~n38319 | ~n39606;
  assign P2_U3095 = ~n37193 | ~n37192;
  assign n37195 = ~n39110 & ~n40906;
  assign n37194 = ~n39230 & ~n37202;
  assign n37201 = ~n37195 & ~n37194;
  assign n37199 = ~n40908 & ~n37205;
  assign n37197 = ~P2_INSTQUEUE_REG_5__2__SCAN_IN | ~n37206;
  assign n37196 = ~n38319 | ~n39233;
  assign P2_U3090 = ~n37201 | ~n37200;
  assign n37204 = ~n39602 & ~n38703;
  assign n37203 = ~n39251 & ~n37202;
  assign n37212 = ~n37204 & ~n37203;
  assign n37210 = ~n39540 & ~n37205;
  assign n37208 = ~P2_INSTQUEUE_REG_5__1__SCAN_IN | ~n37206;
  assign n37207 = ~n39193 | ~n38706;
  assign P2_U3089 = ~n37212 | ~n37211;
  assign n37216 = ~n37536;
  assign n37217 = ~n38804 & ~n42175;
  assign n44008 = n37220 ^ n37219;
  assign n37222 = ~n44008 | ~n43803;
  assign n37221 = ~n43796 | ~P1_EBX_REG_10__SCAN_IN;
  assign n37223 = ~n37222 | ~n37221;
  assign n37225 = ~n43469 & ~n37223;
  assign n37224 = ~n43797 | ~P1_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n37232 = ~n37225 | ~n37224;
  assign n37226 = ~n42400 & ~n37227;
  assign n37229 = n37228 & n38781;
  assign n37230 = ~n38781 & ~P1_REIP_REG_10__SCAN_IN;
  assign n37231 = ~n38790 & ~n37230;
  assign n37233 = ~n37232 & ~n37231;
  assign P1_U2830 = ~n37234 | ~n37233;
  assign n37236 = n42185 | n37235;
  assign n37240 = ~n37237 | ~n37236;
  assign n37239 = ~n42400 & ~n37237;
  assign n37255 = ~n37240 | ~n37507;
  assign n37253 = ~n41129 & ~n37241;
  assign n37244 = ~n37243 & ~n42175;
  assign n37249 = ~n43570 & ~n37246;
  assign n37247 = ~P1_EBX_REG_8__SCAN_IN | ~n43796;
  assign n37248 = ~n37247 | ~n43033;
  assign n37250 = ~n37249 & ~n37248;
  assign P1_U2832 = ~n37255 | ~n37254;
  assign n37257 = ~n41920 | ~P2_REIP_REG_20__SCAN_IN;
  assign n37256 = ~n41921 | ~P2_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n37263 = ~n37257 | ~n37256;
  assign n37258 = ~n37717 | ~n41718;
  assign n37259 = ~n37258 ^ n42473;
  assign n37261 = ~n37259 | ~n41206;
  assign n37260 = ~P2_EBX_REG_20__SCAN_IN | ~n41935;
  assign n37262 = ~n37261 | ~n37260;
  assign n37268 = ~n37263 & ~n37262;
  assign n37266 = ~n42516;
  assign n37276 = ~n42517 | ~n40602;
  assign P2_U2835 = n37278 | n37277;
  assign n37284 = ~n37279 & ~n41888;
  assign n37282 = ~n37280 | ~n40602;
  assign n37281 = ~P2_EBX_REG_0__SCAN_IN | ~n41935;
  assign n37283 = ~n37282 | ~n37281;
  assign n37301 = ~n37284 & ~n37283;
  assign n37299 = ~n40669 & ~n37285;
  assign n37287 = ~n41921 & ~n39732;
  assign n37295 = ~n37287 & ~n37286;
  assign n37293 = ~n37947 | ~n40579;
  assign n37291 = ~n37290;
  assign n37292 = ~n37291 | ~n41934;
  assign n37294 = ~n37293 | ~n37292;
  assign n37297 = ~n37295 & ~n37294;
  assign n37296 = ~n41920 | ~P2_REIP_REG_0__SCAN_IN;
  assign n37298 = ~n37297 | ~n37296;
  assign n37300 = ~n37299 & ~n37298;
  assign P2_U2855 = ~n37301 | ~n37300;
  assign n37307 = ~n37302 & ~n41888;
  assign n37305 = ~n37303 | ~n40602;
  assign n37304 = ~P2_EBX_REG_1__SCAN_IN | ~n41935;
  assign n37306 = ~n37305 | ~n37304;
  assign n37321 = ~n37307 & ~n37306;
  assign n37319 = ~n41926 & ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n37309 = ~n37637 | ~n40579;
  assign n37308 = ~n41921 | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n37314 = ~n37309 | ~n37308;
  assign n37312 = ~n37310 | ~n41934;
  assign n37311 = ~n41920 | ~P2_REIP_REG_1__SCAN_IN;
  assign n37313 = ~n37312 | ~n37311;
  assign n37317 = ~n37314 & ~n37313;
  assign n37316 = ~n41869 | ~n37315;
  assign n37318 = ~n37317 | ~n37316;
  assign n37320 = ~n37319 & ~n37318;
  assign P2_U2854 = ~n37321 | ~n37320;
  assign n37328 = ~n42135 | ~n37322;
  assign n37323 = ~P3_EBX_REG_20__SCAN_IN | ~n43930;
  assign n37326 = ~n37323 | ~n37325;
  assign n37921 = ~n37325 & ~n37324;
  assign P3_U2683 = ~n37328 | ~n37327;
  assign n37331 = ~n37329 | ~n41934;
  assign n37330 = ~n41935 | ~P2_EBX_REG_7__SCAN_IN;
  assign n37333 = ~n37331 | ~n37330;
  assign n37332 = ~n40948 & ~n41926;
  assign n37334 = ~n37333 & ~n37332;
  assign n37336 = ~n41920 | ~P2_REIP_REG_7__SCAN_IN;
  assign n37335 = ~n41921 | ~P2_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n37337 = ~n37336 | ~n37335;
  assign n37347 = ~n37338 & ~n37337;
  assign n37345 = n40775 & n40602;
  assign n37343 = ~n37339 | ~n41942;
  assign n37340 = ~n40948 & ~n39721;
  assign n37341 = ~n37340 & ~n40669;
  assign n37342 = ~n37341 | ~n38941;
  assign n37344 = ~n37343 | ~n37342;
  assign n37346 = ~n37345 & ~n37344;
  assign P2_U2848 = ~n37347 | ~n37346;
  assign n37348 = ~n44044 & ~n43734;
  assign n37350 = ~n40436 | ~n42688;
  assign P1_U2894 = ~n37351 | ~n37350;
  assign n37354 = P2_EBX_REG_16__SCAN_IN & n35967;
  assign n37353 = ~n37352 & ~n33538;
  assign n37358 = ~n37354 & ~n37353;
  assign n37357 = ~n42637 | ~n43525;
  assign P2_U2871 = ~n37358 | ~n37357;
  assign n37375 = ~n39529 & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n37371 = ~n39241 & ~n38769;
  assign n37369 = ~n38773 | ~n39244;
  assign n37361 = ~n37375 & ~n37360;
  assign n37609 = ~n37852;
  assign n38778 = ~n37367 | ~n37366;
  assign n37381 = ~n41307 & ~n39240;
  assign n37377 = ~n37376 & ~n37375;
  assign n37378 = ~n37377 & ~n39511;
  assign n37380 = ~n39515 & ~n38770;
  assign P2_U3160 = ~n37383 | ~n37382;
  assign n37387 = ~n39153 & ~n38769;
  assign n37385 = ~n38773 | ~n39156;
  assign n37389 = ~n41307 & ~n40883;
  assign n37388 = ~n40882 & ~n38770;
  assign P2_U3165 = ~n37391 | ~n37390;
  assign n37395 = ~n39251 & ~n38769;
  assign n37393 = ~n38773 | ~n39542;
  assign n37397 = ~n41307 & ~n39549;
  assign n37396 = ~n39540 & ~n38770;
  assign P2_U3161 = ~n37399 | ~n37398;
  assign n37405 = ~n41290 & ~n38280;
  assign n37401 = ~n38208 & ~n41283;
  assign n37400 = ~n41289 & ~n37416;
  assign n37403 = ~n37401 & ~n37400;
  assign n37402 = ~n41284 | ~n38294;
  assign P2_U3127 = ~n37407 | ~n37406;
  assign n37413 = ~n39549 & ~n38280;
  assign n37409 = ~n38208 & ~n38703;
  assign n37408 = ~n39540 & ~n37416;
  assign n37411 = ~n37409 & ~n37408;
  assign n37410 = ~n39541 | ~n38294;
  assign n37415 = ~n37413 & ~n37412;
  assign P2_U3121 = ~n37415 | ~n37414;
  assign n37422 = ~n40906 & ~n38280;
  assign n37418 = ~n38208 & ~n40907;
  assign n37417 = ~n40908 & ~n37416;
  assign n37420 = ~n37418 & ~n37417;
  assign n37419 = ~n40911 | ~n38294;
  assign P2_U3122 = ~n37425 | ~n37424;
  assign n37431 = ~n40906 & ~n37854;
  assign n37427 = ~n39187 & ~n40907;
  assign n37426 = ~n40908 & ~n37539;
  assign n37429 = ~n37427 & ~n37426;
  assign n37428 = ~n40911 | ~n37542;
  assign n37432 = ~P2_INSTQUEUE_REG_7__2__SCAN_IN | ~n37547;
  assign P2_U3106 = ~n37433 | ~n37432;
  assign n37436 = ~P2_EAX_REG_17__SCAN_IN | ~n43698;
  assign n37435 = ~n42804 | ~n37434;
  assign n37440 = ~n37436 | ~n37435;
  assign n37438 = ~BUF2_REG_17__SCAN_IN | ~n43689;
  assign n37437 = ~BUF1_REG_17__SCAN_IN | ~n43690;
  assign n37439 = ~n37438 | ~n37437;
  assign n37449 = ~n37440 & ~n37439;
  assign n37443 = n37442 | n37441;
  assign n37447 = ~n37827 & ~n41754;
  assign n37446 = ~n42612 & ~n43695;
  assign P2_U2902 = ~n37449 | ~n37448;
  assign n37451 = ~n41920 | ~P2_REIP_REG_21__SCAN_IN;
  assign n37450 = ~n41921 | ~P2_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n37458 = ~n37451 | ~n37450;
  assign n37453 = ~n41204 & ~n37452;
  assign n37454 = ~n37453 ^ n42856;
  assign n37456 = ~n37454 | ~n41206;
  assign n37455 = ~P2_EBX_REG_21__SCAN_IN | ~n41935;
  assign n37457 = ~n37456 | ~n37455;
  assign n37463 = ~n37458 & ~n37457;
  assign n37462 = ~n37461 | ~n41942;
  assign n37465 = ~n37464;
  assign n42723 = ~n39701 & ~n37467;
  assign n37471 = ~n42723 | ~n40602;
  assign P2_U2834 = n37473 | n37472;
  assign n37480 = ~n34242 | ~n38884;
  assign n38057 = ~n37485 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n39819 = ~n38057;
  assign n38062 = ~n39310 & ~n37475;
  assign n37478 = ~n39819 | ~n38062;
  assign n37477 = ~n39315 | ~n37488;
  assign n37479 = ~n39962 | ~n38885;
  assign n37484 = ~n37480 | ~n37479;
  assign n37482 = ~n39939 | ~n38894;
  assign n37481 = ~n39967 | ~n38889;
  assign n37483 = ~n37482 | ~n37481;
  assign n37495 = ~n37484 & ~n37483;
  assign n39956 = ~n37485 & ~n43722;
  assign P1_U3145 = ~n37495 | ~n37494;
  assign n37497 = n43362 & n37516;
  assign n37506 = ~n37497 & ~n37496;
  assign n37504 = n43709 & P1_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign P1_U2990 = ~n37506 | ~n37505;
  assign n37510 = ~n37508 | ~n37507;
  assign n37522 = ~n37510 | ~n37509;
  assign n37514 = ~n43570 & ~n37550;
  assign n37512 = ~n43796 | ~P1_EBX_REG_9__SCAN_IN;
  assign n37511 = ~n43797 | ~P1_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n37513 = ~n37512 | ~n37511;
  assign n37515 = ~n37514 & ~n37513;
  assign n37518 = ~n37551 | ~n41453;
  assign n37517 = ~n43559 | ~n37516;
  assign P1_U2831 = ~n37522 | ~n37521;
  assign n37528 = ~n39200 & ~n37596;
  assign n37524 = ~n38221 & ~n41302;
  assign n37523 = ~n41301 & ~n37597;
  assign n37526 = ~n37524 & ~n37523;
  assign n37525 = ~n37839 | ~n39201;
  assign P2_U3062 = ~n37530 | ~n37529;
  assign n39646 = n37532 ^ n37531;
  assign n37534 = ~n39646 | ~n44021;
  assign n37533 = ~P1_EBX_REG_11__SCAN_IN | ~n44023;
  assign n37538 = n37534 & n37533;
  assign P1_U2861 = ~n37538 | ~n37537;
  assign n37546 = ~n39240 & ~n37854;
  assign n37541 = ~n39187 & ~n39535;
  assign n37540 = ~n39515 & ~n37539;
  assign n37544 = ~n37541 & ~n37540;
  assign n37543 = ~n39516 | ~n37542;
  assign n37548 = ~P2_INSTQUEUE_REG_7__0__SCAN_IN | ~n37547;
  assign P2_U3104 = ~n37549 | ~n37548;
  assign n37553 = ~n37550 & ~n43298;
  assign n37552 = ~n37846 & ~n44019;
  assign n37554 = ~P1_EBX_REG_9__SCAN_IN | ~n44023;
  assign P1_U2863 = ~n37555 | ~n37554;
  assign n37565 = ~n37556 & ~n43924;
  assign n37559 = ~n40574 | ~n43896;
  assign n37560 = ~n37559 | ~n37558;
  assign n37562 = ~n43917 | ~P2_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n37566 = ~n43813 | ~n40565;
  assign P2_U3010 = ~n37567 | ~n37566;
  assign n40470 = ~n40421 & ~n40431;
  assign n37576 = ~n41095 | ~n37575;
  assign n37582 = ~n37577 | ~n37576;
  assign n37579 = n37578 & n41100;
  assign n37581 = ~n37753 & ~n37579;
  assign n37580 = ~n37748 | ~n38140;
  assign n38156 = ~n37581 | ~n37580;
  assign n37586 = ~n37582 | ~n38156;
  assign n38157 = ~n41403 & ~P3_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n37583 = n41400 | n38157;
  assign n37585 = ~n37584 | ~n37583;
  assign n37587 = ~n37586 | ~n37585;
  assign n37592 = ~n40744 | ~n40410;
  assign P3_U2810 = ~n37595 | ~n37594;
  assign n37603 = ~n39268 & ~n37596;
  assign n37599 = ~n38221 & ~n41318;
  assign n37598 = ~n41317 & ~n37597;
  assign n37601 = ~n37599 & ~n37598;
  assign n37600 = ~n37839 | ~n39271;
  assign P2_U3060 = ~n37606 | ~n37605;
  assign n39548 = ~n39507 & ~n38279;
  assign n37607 = n39548 | n37839;
  assign n38323 = ~n37853 & ~n37609;
  assign n37611 = ~n37834;
  assign n37613 = ~n37612 & ~n37611;
  assign n37614 = ~n37613 & ~n39511;
  assign n37617 = ~n37835 & ~n39515;
  assign n37616 = ~n39241 & ~n37834;
  assign n37619 = ~n37617 & ~n37616;
  assign n37618 = ~n37839 | ~n39517;
  assign n37622 = ~n37620;
  assign n37632 = ~n39548 | ~n39244;
  assign P2_U3048 = ~n37633 | ~n37632;
  assign n37636 = ~n37634 | ~n38277;
  assign n37649 = ~n39268 & ~n37933;
  assign n37647 = ~n39607 | ~n38678;
  assign n37646 = ~P2_INSTQUEUE_REG_3__4__SCAN_IN | ~n37941;
  assign n37661 = ~n37649 & ~n37648;
  assign n37659 = ~n39015 & ~n41308;
  assign n37652 = ~n38220;
  assign n37653 = ~n37933;
  assign n37655 = ~n37654 & ~n37653;
  assign n37656 = ~n37655 & ~n39511;
  assign n37658 = ~n41317 & ~n37934;
  assign n37660 = ~n37659 & ~n37658;
  assign P2_U3076 = ~n37661 | ~n37660;
  assign n37663 = ~n39015 & ~n40895;
  assign n37662 = ~n39280 & ~n37933;
  assign n37669 = ~n37663 & ~n37662;
  assign n37667 = ~n40896 & ~n37934;
  assign n37665 = ~P2_INSTQUEUE_REG_3__3__SCAN_IN | ~n37941;
  assign n37664 = ~n39607 | ~n38669;
  assign n37666 = ~n37665 | ~n37664;
  assign n37668 = ~n37667 & ~n37666;
  assign P2_U3075 = ~n37669 | ~n37668;
  assign n37671 = ~n39015 & ~n38703;
  assign n37670 = ~n39251 & ~n37933;
  assign n37677 = ~n37671 & ~n37670;
  assign n37675 = ~n39540 & ~n37934;
  assign n37673 = ~P2_INSTQUEUE_REG_3__1__SCAN_IN | ~n37941;
  assign n37672 = ~n39607 | ~n38706;
  assign n37674 = ~n37673 | ~n37672;
  assign n37676 = ~n37675 & ~n37674;
  assign P2_U3073 = ~n37677 | ~n37676;
  assign n37679 = ~n39015 & ~n41283;
  assign n37678 = ~n39601 & ~n37933;
  assign n37685 = ~n37679 & ~n37678;
  assign n37683 = ~n41289 & ~n37934;
  assign n37681 = ~P2_INSTQUEUE_REG_3__7__SCAN_IN | ~n37941;
  assign n37680 = ~n39607 | ~n37808;
  assign n37682 = ~n37681 | ~n37680;
  assign n37684 = ~n37683 & ~n37682;
  assign P2_U3079 = ~n37685 | ~n37684;
  assign n37687 = ~n39015 & ~n41295;
  assign n37686 = ~n39200 & ~n37933;
  assign n37693 = ~n37687 & ~n37686;
  assign n37691 = ~n41301 & ~n37934;
  assign n37689 = ~P2_INSTQUEUE_REG_3__6__SCAN_IN | ~n37941;
  assign n37688 = ~n39607 | ~n38696;
  assign n37690 = ~n37689 | ~n37688;
  assign n37692 = ~n37691 & ~n37690;
  assign P2_U3078 = ~n37693 | ~n37692;
  assign n37695 = ~n37694 | ~n38155;
  assign n37697 = ~n37696 | ~n37695;
  assign n37705 = ~n37697 | ~P3_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n37699 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN | ~n37698;
  assign n37703 = ~n37699 & ~P3_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n37701 = ~n37700 | ~n41400;
  assign n40348 = ~n41145 | ~P3_REIP_REG_16__SCAN_IN;
  assign n37702 = ~n37701 | ~n40348;
  assign n37704 = ~n37703 & ~n37702;
  assign n37708 = ~n37705 | ~n37704;
  assign n37707 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN & ~n37706;
  assign n37712 = ~n37708 & ~n37707;
  assign n37709 = n41149 ^ P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n37711 = ~n40857 | ~n40335;
  assign n37715 = n37712 & n37711;
  assign n37714 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN | ~n37713;
  assign P3_U2814 = ~n37715 | ~n37714;
  assign n37719 = ~n37716 & ~n42345;
  assign n37718 = ~n41869 | ~n37717;
  assign n37734 = ~n37719 & ~n37718;
  assign n37722 = ~n41926 & ~n42345;
  assign n37720 = ~P2_REIP_REG_19__SCAN_IN | ~n41920;
  assign n37721 = ~n37720 | ~n40668;
  assign n37724 = ~n37722 & ~n37721;
  assign n37723 = ~P2_PHYADDRPOINTER_REG_19__SCAN_IN | ~n41921;
  assign n37737 = ~n42352 | ~n41934;
  assign P2_U2836 = ~n37738 | ~n37737;
  assign n37741 = ~n37835 & ~n40908;
  assign n37740 = ~n39230 & ~n37834;
  assign n37742 = ~n37839 | ~n38715;
  assign n37746 = ~n39548 | ~n39233;
  assign P2_U3050 = ~n37747 | ~n37746;
  assign n37770 = ~n39420 & ~n40820;
  assign n37751 = ~n37748 | ~n38909;
  assign n37750 = ~n41100 | ~n37749;
  assign n37752 = ~n37751 | ~n37750;
  assign n38918 = ~n37753 & ~n37752;
  assign n37755 = n41095 & n37754;
  assign n37756 = ~P3_PHYADDRPOINTER_REG_23__SCAN_IN & ~n37755;
  assign n37764 = ~n38918 & ~n37756;
  assign n40237 = ~n40865 & ~n37757;
  assign n37762 = ~n40237;
  assign n38917 = ~n40726 | ~n37758;
  assign n37759 = ~n41520 | ~n38917;
  assign n37761 = ~n37760 | ~n37759;
  assign n37763 = ~n37762 | ~n37761;
  assign n37768 = ~n37764 & ~n37763;
  assign n37771 = ~n39785;
  assign n37773 = ~n39790;
  assign n37775 = ~n37774 | ~n37773;
  assign P3_U2807 = ~n37779 | ~n37778;
  assign n37785 = ~n39251 & ~n37834;
  assign n37781 = ~n39540 & ~n37835;
  assign n37780 = ~n37836 & ~n41597;
  assign n37786 = ~n39548 | ~n39542;
  assign P2_U3049 = ~n37787 | ~n37786;
  assign n37793 = ~n39200 & ~n37834;
  assign n37789 = ~n41301 & ~n37835;
  assign n37788 = ~n35254 & ~n37836;
  assign n37794 = ~n39548 | ~n39201;
  assign P2_U3054 = ~n37795 | ~n37794;
  assign n37802 = ~n39280 & ~n37834;
  assign n37798 = ~n40896 & ~n37835;
  assign n37797 = ~n37836 & ~n37796;
  assign n37803 = ~n39548 | ~n39285;
  assign P2_U3051 = ~n37804 | ~n37803;
  assign n37812 = ~n39601 & ~n37834;
  assign n37807 = ~n41289 & ~n37835;
  assign n37806 = ~n37805 & ~n37836;
  assign n37813 = ~n39548 | ~n39606;
  assign P2_U3055 = ~n37814 | ~n37813;
  assign n37820 = ~n39153 & ~n37834;
  assign n37816 = ~n40882 & ~n37835;
  assign n37815 = ~n37836 & ~n43091;
  assign n37821 = ~n39548 | ~n39156;
  assign P2_U3053 = ~n37822 | ~n37821;
  assign n37824 = ~n40436 | ~n42736;
  assign n37823 = ~P1_EAX_REG_11__SCAN_IN | ~n43732;
  assign n37826 = n37824 & n37823;
  assign P1_U2893 = ~n37826 | ~n37825;
  assign n37829 = P2_EBX_REG_17__SCAN_IN & n35967;
  assign n37828 = ~n37827 & ~n33538;
  assign n37833 = ~n37829 & ~n37828;
  assign n37832 = ~n42616 | ~n43525;
  assign P2_U2870 = ~n37833 | ~n37832;
  assign n37843 = ~n39268 & ~n37834;
  assign n37838 = ~n41317 & ~n37835;
  assign n37837 = ~n37836 & ~n42782;
  assign n37844 = ~n39548 | ~n39271;
  assign P2_U3052 = ~n37845 | ~n37844;
  assign n37847 = ~n44049 & ~n43734;
  assign n37849 = ~n40436 | ~n42029;
  assign P1_U2895 = ~n37850 | ~n37849;
  assign n37865 = ~n39230 & ~n38207;
  assign n37863 = ~n38212 | ~n39233;
  assign n38324 = ~n37951;
  assign n37950 = ~n37853 | ~n37852;
  assign n37866 = ~n38324 & ~n37950;
  assign n37869 = ~n38207;
  assign n37875 = ~n38208 & ~n40906;
  assign n37867 = ~n37866;
  assign n37871 = ~n37870 & ~n37869;
  assign n37872 = ~n37871 & ~n39511;
  assign n37874 = ~n40908 & ~n38209;
  assign P2_U3114 = ~n37877 | ~n37876;
  assign n37881 = ~n39251 & ~n38207;
  assign n37879 = ~n38212 | ~n39542;
  assign n37883 = ~n38208 & ~n39549;
  assign n37882 = ~n39540 & ~n38209;
  assign P2_U3113 = ~n37885 | ~n37884;
  assign n37889 = ~n39241 & ~n38207;
  assign n37887 = ~n38212 | ~n39244;
  assign n37891 = ~n38208 & ~n39240;
  assign n37890 = ~n39515 & ~n38209;
  assign P2_U3112 = ~n37893 | ~n37892;
  assign n37897 = ~n39200 & ~n38207;
  assign n37895 = ~n38212 | ~n39201;
  assign n37899 = ~n38208 & ~n41302;
  assign n37898 = ~n41301 & ~n38209;
  assign P2_U3118 = ~n37901 | ~n37900;
  assign n37907 = ~n39230 & ~n37933;
  assign n37903 = ~n39015 & ~n40907;
  assign n37902 = ~n40908 & ~n37934;
  assign n37905 = ~n37903 & ~n37902;
  assign n37904 = ~n39607 | ~n38715;
  assign n37908 = ~P2_INSTQUEUE_REG_3__2__SCAN_IN | ~n37941;
  assign P2_U3074 = ~n37909 | ~n37908;
  assign n37915 = ~n39241 & ~n37933;
  assign n37911 = ~n39015 & ~n39535;
  assign n37910 = ~n39515 & ~n37934;
  assign n37913 = ~n37911 & ~n37910;
  assign n37912 = ~n39607 | ~n39517;
  assign n37916 = ~P2_INSTQUEUE_REG_3__0__SCAN_IN | ~n37941;
  assign P2_U3072 = ~n37917 | ~n37916;
  assign n37924 = ~n42135 | ~n37918;
  assign n37920 = ~P3_EBX_REG_21__SCAN_IN | ~n43930;
  assign n39503 = ~n37921 | ~P3_EBX_REG_21__SCAN_IN;
  assign n37923 = ~n37922 | ~n39503;
  assign P3_U2682 = ~n37924 | ~n37923;
  assign n37928 = ~n39153 & ~n38207;
  assign n37926 = ~n38212 | ~n39156;
  assign n37930 = ~n38208 & ~n40883;
  assign n37929 = ~n40882 & ~n38209;
  assign P2_U3117 = ~n37932 | ~n37931;
  assign n37940 = ~n39153 & ~n37933;
  assign n37936 = ~n39015 & ~n40881;
  assign n37935 = ~n40882 & ~n37934;
  assign n37938 = ~n37936 & ~n37935;
  assign n37937 = ~n39607 | ~n38687;
  assign n37943 = ~n37940 & ~n37939;
  assign n37942 = ~P2_INSTQUEUE_REG_3__5__SCAN_IN | ~n37941;
  assign P2_U3077 = ~n37943 | ~n37942;
  assign n37960 = ~n39251 & ~n38304;
  assign n37958 = ~n38933 | ~n39542;
  assign n37961 = ~n37951 & ~n37950;
  assign n37964 = ~n38304;
  assign n37954 = ~n37964 & ~n37953;
  assign n37970 = ~n38305 & ~n39549;
  assign n37962 = ~n37961;
  assign n37966 = ~n37965 & ~n37964;
  assign n37967 = ~n37966 & ~n39511;
  assign n37969 = ~n39540 & ~n38306;
  assign P2_U3145 = ~n37972 | ~n37971;
  assign n37974 = ~n38305 & ~n39240;
  assign n37973 = ~n39241 & ~n38304;
  assign n37980 = ~n37974 & ~n37973;
  assign n37978 = ~n39515 & ~n38306;
  assign n37975 = ~n38933 | ~n39244;
  assign P2_U3144 = ~n37980 | ~n37979;
  assign n37982 = ~n38305 & ~n41290;
  assign n37981 = ~n39601 & ~n38304;
  assign n37988 = ~n37982 & ~n37981;
  assign n37986 = ~n41289 & ~n38306;
  assign n37983 = ~n38933 | ~n39606;
  assign P2_U3151 = ~n37988 | ~n37987;
  assign n37990 = ~n38305 & ~n40894;
  assign n37989 = ~n39280 & ~n38304;
  assign n37996 = ~n37990 & ~n37989;
  assign n37994 = ~n40896 & ~n38306;
  assign n37991 = ~n38933 | ~n39285;
  assign P2_U3147 = ~n37996 | ~n37995;
  assign n37998 = ~n38305 & ~n40883;
  assign n37997 = ~n39153 & ~n38304;
  assign n38004 = ~n37998 & ~n37997;
  assign n38002 = ~n40882 & ~n38306;
  assign n37999 = ~n38933 | ~n39156;
  assign P2_U3149 = ~n38004 | ~n38003;
  assign n38006 = ~n38305 & ~n40906;
  assign n38005 = ~n39230 & ~n38304;
  assign n38012 = ~n38006 & ~n38005;
  assign n38010 = ~n40908 & ~n38306;
  assign n38007 = ~n38933 | ~n39233;
  assign P2_U3146 = ~n38012 | ~n38011;
  assign n38026 = n42287 & n41756;
  assign n38017 = ~BUF2_REG_18__SCAN_IN;
  assign n38022 = ~n42802 & ~n38017;
  assign n38020 = ~n42804 | ~n38018;
  assign n38019 = ~n43698 | ~P2_EAX_REG_18__SCAN_IN;
  assign n38021 = ~n38020 | ~n38019;
  assign n38024 = ~n38022 & ~n38021;
  assign n38023 = ~n43690 | ~BUF1_REG_18__SCAN_IN;
  assign n38025 = ~n38024 | ~n38023;
  assign P2_U2901 = ~n38028 | ~n38027;
  assign n38046 = ~n40421 & ~n38029;
  assign n38032 = ~n38031 | ~n38155;
  assign n38034 = ~n38033 | ~n38032;
  assign n38041 = ~n38034 | ~P3_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n38036 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN | ~n38035;
  assign n38039 = ~n38036 & ~P3_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n38038 = ~n38037 & ~n41520;
  assign n38040 = ~n38039 & ~n38038;
  assign n38042 = ~n38041 | ~n38040;
  assign n40434 = ~n41145 | ~P3_REIP_REG_19__SCAN_IN;
  assign P3_U2811 = ~n38049 | ~n38048;
  assign n38122 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n38050;
  assign n38052 = ~n34188 | ~n38122;
  assign n38051 = ~n39970 | ~n38123;
  assign n38071 = ~n38052 | ~n38051;
  assign n38055 = ~n39307 & ~n38122;
  assign n38060 = ~n38059 & ~n39953;
  assign n38067 = ~n39956 | ~n38062;
  assign n38065 = ~n38063;
  assign n38072 = ~n39978 | ~n38132;
  assign P1_U3114 = ~n38073 | ~n38072;
  assign n38075 = ~n34150 | ~n38122;
  assign n38074 = ~n40025 | ~n38123;
  assign n38079 = ~n38075 | ~n38074;
  assign n38080 = ~n40033 | ~n38132;
  assign P1_U3119 = ~n38081 | ~n38080;
  assign n38083 = ~n34135 | ~n38122;
  assign n38082 = ~n39981 | ~n38123;
  assign n38087 = ~n38083 | ~n38082;
  assign n38088 = ~n39989 | ~n38132;
  assign P1_U3117 = ~n38089 | ~n38088;
  assign n38091 = ~n34098 | ~n38122;
  assign n38090 = ~n40038 | ~n38123;
  assign n38095 = ~n38091 | ~n38090;
  assign n38096 = ~n40049 | ~n38132;
  assign P1_U3118 = ~n38097 | ~n38096;
  assign n38099 = ~n34227 | ~n38122;
  assign n38098 = ~n40003 | ~n38123;
  assign n38103 = ~n38099 | ~n38098;
  assign n38104 = ~n40011 | ~n38132;
  assign P1_U3115 = ~n38105 | ~n38104;
  assign n38107 = ~n34242 | ~n38122;
  assign n38106 = ~n39939 | ~n38123;
  assign n38111 = ~n38107 | ~n38106;
  assign n38112 = ~n39967 | ~n38132;
  assign P1_U3113 = ~n38113 | ~n38112;
  assign n38115 = ~n34165 | ~n38122;
  assign n38114 = ~n39992 | ~n38123;
  assign n38119 = ~n38115 | ~n38114;
  assign n38120 = ~n40000 | ~n38132;
  assign P1_U3116 = ~n38121 | ~n38120;
  assign n38125 = ~n34072 | ~n38122;
  assign n38124 = ~n40014 | ~n38123;
  assign n38131 = ~n38125 | ~n38124;
  assign n38133 = ~n40022 | ~n38132;
  assign P1_U3120 = ~n38134 | ~n38133;
  assign n38137 = ~n42439 | ~n43525;
  assign n38136 = n43525 | P2_EBX_REG_18__SCAN_IN;
  assign P2_U2869 = ~n38139 | ~n38138;
  assign n38180 = ~n38140 & ~n40872;
  assign n38141 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN | ~n38180;
  assign n38166 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN & ~n38141;
  assign n38145 = ~n38143;
  assign n38146 = ~n38145 | ~n38144;
  assign n38162 = ~n38154 & ~n41520;
  assign n38179 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n38158 = ~n38179 | ~n38155;
  assign n38171 = ~n38157 & ~n38156;
  assign n38159 = ~n38158 | ~n38171;
  assign n38160 = ~n38159 | ~P3_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n39803 = ~n41145 | ~P3_REIP_REG_22__SCAN_IN;
  assign n38161 = ~n38160 | ~n39803;
  assign n38163 = ~n38162 & ~n38161;
  assign P3_U2808 = ~n38170 | ~n38169;
  assign n38187 = ~n38171 & ~n38179;
  assign n40533 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN | ~n40531;
  assign n38183 = ~n41520 & ~n38178;
  assign n40540 = ~n41145 | ~P3_REIP_REG_21__SCAN_IN;
  assign n38181 = ~n38180 | ~n38179;
  assign n38182 = ~n40540 | ~n38181;
  assign n38184 = ~n38183 & ~n38182;
  assign P3_U2809 = ~n38190 | ~n38189;
  assign n38196 = ~n39280 & ~n38207;
  assign n38192 = ~n38208 & ~n40894;
  assign n38191 = ~n40896 & ~n38209;
  assign n38193 = ~n38212 | ~n39285;
  assign P2_U3115 = ~n38198 | ~n38197;
  assign n38204 = ~n39601 & ~n38207;
  assign n38200 = ~n38208 & ~n41290;
  assign n38199 = ~n41289 & ~n38209;
  assign n38201 = ~n38212 | ~n39606;
  assign P2_U3119 = ~n38206 | ~n38205;
  assign n38216 = ~n39268 & ~n38207;
  assign n38211 = ~n38208 & ~n41318;
  assign n38210 = ~n41317 & ~n38209;
  assign n38213 = ~n38212 | ~n39271;
  assign P2_U3116 = ~n38219 | ~n38218;
  assign n38234 = ~n39241 & ~n39016;
  assign n38230 = ~n39015 & ~n39240;
  assign n38225 = ~n39016;
  assign n38224 = ~n38225 & ~n38235;
  assign n38226 = ~n38237 & ~n38225;
  assign n38227 = ~n38226 & ~n39511;
  assign n39019 = ~n38228 & ~n38227;
  assign n38229 = ~n39515 & ~n39019;
  assign n38231 = ~n39021 | ~n39244;
  assign n38240 = n38236 | n38235;
  assign P2_U3064 = ~n38244 | ~n38243;
  assign n38250 = ~n39251 & ~n39016;
  assign n38246 = ~n39015 & ~n39549;
  assign n38245 = ~n39540 & ~n39019;
  assign n38247 = ~n39021 | ~n39542;
  assign P2_U3065 = ~n38252 | ~n38251;
  assign n38255 = ~n43803 | ~n38662;
  assign n38254 = ~P1_REIP_REG_12__SCAN_IN | ~n38253;
  assign n38264 = ~n38255 | ~n38254;
  assign n38257 = ~P1_REIP_REG_12__SCAN_IN & ~n38256;
  assign n38259 = ~n38257 | ~n38781;
  assign n38258 = ~n43796 | ~P1_EBX_REG_12__SCAN_IN;
  assign n38260 = ~n38259 | ~n38258;
  assign n38262 = ~n43469 & ~n38260;
  assign n38261 = ~n43797 | ~P1_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n38263 = ~n38262 | ~n38261;
  assign n38268 = ~n38264 & ~n38263;
  assign n38265 = ~n38389 & ~n42175;
  assign P1_U2828 = ~n38268 | ~n38267;
  assign n38274 = ~n39200 & ~n38304;
  assign n38270 = ~n38305 & ~n41302;
  assign n38269 = ~n41301 & ~n38306;
  assign n38271 = ~n38933 | ~n39201;
  assign P2_U3150 = ~n38276 | ~n38275;
  assign n38278 = ~n38277 & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n38617 = ~n38626;
  assign n38293 = ~n39153 & ~n39279;
  assign n39278 = ~n38615 | ~n38279;
  assign n38289 = ~n39278 & ~n40883;
  assign n38284 = ~n39279;
  assign n38283 = ~n38284 & ~n38294;
  assign n38285 = ~n38296 & ~n38284;
  assign n38286 = ~n38285 & ~n39511;
  assign n38288 = ~n40882 & ~n39283;
  assign n38290 = ~n39286 | ~n39156;
  assign n38299 = n38295 | n38294;
  assign P2_U3133 = ~n38303 | ~n38302;
  assign n38312 = ~n39268 & ~n38304;
  assign n38308 = ~n38305 & ~n41318;
  assign n38307 = ~n41317 & ~n38306;
  assign n38309 = ~n38933 | ~n39271;
  assign P2_U3148 = ~n38315 | ~n38314;
  assign n38318 = ~n39602 & ~n40906;
  assign n38332 = ~n38316 & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n38317 = ~n39230 & ~n39600;
  assign n38344 = ~n38318 & ~n38317;
  assign n38335 = ~n38324 | ~n38323;
  assign n38326 = ~n38329 & ~n38332;
  assign n38327 = ~n38326 & ~n39511;
  assign n39603 = ~n38328 & ~n38327;
  assign n38342 = ~n40908 & ~n39603;
  assign n38333 = ~n38332 & ~n38331;
  assign n38338 = ~n38334 & ~n38333;
  assign n38339 = ~n39607 | ~n39233;
  assign P2_U3082 = ~n38344 | ~n38343;
  assign n38346 = ~n39602 & ~n40894;
  assign n38345 = ~n39280 & ~n39600;
  assign n38352 = ~n38346 & ~n38345;
  assign n38350 = ~n40896 & ~n39603;
  assign n38347 = ~n39607 | ~n39285;
  assign P2_U3083 = ~n38352 | ~n38351;
  assign n38354 = ~n39602 & ~n39549;
  assign n38353 = ~n39251 & ~n39600;
  assign n38360 = ~n38354 & ~n38353;
  assign n38358 = ~n39540 & ~n39603;
  assign n38355 = ~n39607 | ~n39542;
  assign P2_U3081 = ~n38360 | ~n38359;
  assign n38362 = ~n39602 & ~n41302;
  assign n38361 = ~n39200 & ~n39600;
  assign n38368 = ~n38362 & ~n38361;
  assign n38366 = ~n41301 & ~n39603;
  assign n38363 = ~n39607 | ~n39201;
  assign P2_U3086 = ~n38368 | ~n38367;
  assign n38371 = ~n43911 & ~n40363;
  assign n39653 = ~n43880 | ~P2_REIP_REG_5__SCAN_IN;
  assign n38369 = ~n43917 | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n38370 = ~n39653 | ~n38369;
  assign n38382 = ~n38371 & ~n38370;
  assign n38375 = n38373 | n38372;
  assign n39652 = ~n38375 | ~n38374;
  assign n38380 = ~n39652 & ~n43811;
  assign n38378 = ~n43813 | ~n40368;
  assign P2_U3009 = ~n38382 | ~n38381;
  assign n38387 = ~n38384 | ~n38383;
  assign n38386 = ~n40094 & ~n38385;
  assign n38391 = ~n38388 | ~n43367;
  assign n38390 = n43713 | n38389;
  assign n38660 = ~n43469 | ~P1_REIP_REG_12__SCAN_IN;
  assign n38392 = ~n43709 | ~P1_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n38393 = ~n38660 | ~n38392;
  assign P1_U2987 = ~n38396 | ~n38395;
  assign n38468 = ~n38397 & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n38399 = ~n34150 | ~n38468;
  assign n38398 = ~n40033 | ~n38469;
  assign n38417 = ~n38399 | ~n38398;
  assign n38400 = ~n38482;
  assign n38404 = ~n38468;
  assign n38405 = ~n38404 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n38408 = ~n39310;
  assign n39957 = ~n39311 & ~n38408;
  assign n39954 = n39957 | n43722;
  assign n38413 = ~n39957 | ~n39819;
  assign n38418 = ~n40025 | ~n38478;
  assign P1_U3071 = ~n38419 | ~n38418;
  assign n38421 = ~n34135 | ~n38468;
  assign n38420 = ~n39989 | ~n38469;
  assign n38425 = ~n38421 | ~n38420;
  assign n38426 = ~n39981 | ~n38478;
  assign P1_U3069 = ~n38427 | ~n38426;
  assign n38429 = ~n34098 | ~n38468;
  assign n38428 = ~n40049 | ~n38469;
  assign n38433 = ~n38429 | ~n38428;
  assign n38434 = ~n40038 | ~n38478;
  assign P1_U3070 = ~n38435 | ~n38434;
  assign n38437 = ~n34188 | ~n38468;
  assign n38436 = ~n39978 | ~n38469;
  assign n38441 = ~n38437 | ~n38436;
  assign n38442 = ~n39970 | ~n38478;
  assign P1_U3066 = ~n38443 | ~n38442;
  assign n38445 = ~n34242 | ~n38468;
  assign n38444 = ~n39967 | ~n38469;
  assign n38449 = ~n38445 | ~n38444;
  assign n38450 = ~n39939 | ~n38478;
  assign P1_U3065 = ~n38451 | ~n38450;
  assign n38453 = ~n34072 | ~n38468;
  assign n38452 = ~n40022 | ~n38469;
  assign n38457 = ~n38453 | ~n38452;
  assign n38458 = ~n40014 | ~n38478;
  assign P1_U3072 = ~n38459 | ~n38458;
  assign n38461 = ~n34165 | ~n38468;
  assign n38460 = ~n40000 | ~n38469;
  assign n38465 = ~n38461 | ~n38460;
  assign n38466 = ~n39992 | ~n38478;
  assign P1_U3068 = ~n38467 | ~n38466;
  assign n38471 = ~n34227 | ~n38468;
  assign n38470 = ~n40011 | ~n38469;
  assign n38477 = ~n38471 | ~n38470;
  assign n38479 = ~n40003 | ~n38478;
  assign P1_U3067 = ~n38480 | ~n38479;
  assign n38483 = ~n38481 | ~n39937;
  assign n38552 = ~n38483;
  assign n38488 = ~n34072 | ~n38552;
  assign n39029 = ~n39310 & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n38486 = ~n39819 | ~n39029;
  assign n38485 = n39946 | n38492;
  assign n38487 = ~n40017 | ~n38553;
  assign n38501 = ~n38488 | ~n38487;
  assign n38496 = ~n38552 & ~n39307;
  assign n39041 = n39029 | n43722;
  assign n38498 = ~n40014 | ~n38557;
  assign n38503 = ~n38501 & ~n38500;
  assign n38502 = ~n40022 | ~n38562;
  assign P1_U3088 = ~n38503 | ~n38502;
  assign n38505 = ~n34165 | ~n38552;
  assign n38504 = ~n39995 | ~n38553;
  assign n38509 = ~n38505 | ~n38504;
  assign n38506 = ~n40000 | ~n38562;
  assign n38511 = ~n38509 & ~n38508;
  assign n38510 = ~n39992 | ~n38557;
  assign P1_U3084 = ~n38511 | ~n38510;
  assign n38513 = ~n34098 | ~n38552;
  assign n38512 = ~n40043 | ~n38553;
  assign n38517 = ~n38513 | ~n38512;
  assign n38514 = ~n40049 | ~n38562;
  assign n38519 = ~n38517 & ~n38516;
  assign n38518 = ~n40038 | ~n38557;
  assign P1_U3086 = ~n38519 | ~n38518;
  assign n38521 = ~n34188 | ~n38552;
  assign n38520 = ~n39973 | ~n38553;
  assign n38525 = ~n38521 | ~n38520;
  assign n38522 = ~n39970 | ~n38557;
  assign n38527 = ~n38525 & ~n38524;
  assign n38526 = ~n39978 | ~n38562;
  assign P1_U3082 = ~n38527 | ~n38526;
  assign n38529 = ~n34242 | ~n38552;
  assign n38528 = ~n39962 | ~n38553;
  assign n38533 = ~n38529 | ~n38528;
  assign n38530 = ~n39967 | ~n38562;
  assign n38535 = ~n38533 & ~n38532;
  assign n38534 = ~n39939 | ~n38557;
  assign P1_U3081 = ~n38535 | ~n38534;
  assign n38537 = ~n34227 | ~n38552;
  assign n38536 = ~n40006 | ~n38553;
  assign n38541 = ~n38537 | ~n38536;
  assign n38538 = ~n40003 | ~n38557;
  assign n38543 = ~n38541 & ~n38540;
  assign n38542 = ~n40011 | ~n38562;
  assign P1_U3083 = ~n38543 | ~n38542;
  assign n38545 = ~n34135 | ~n38552;
  assign n38544 = ~n39984 | ~n38553;
  assign n38549 = ~n38545 | ~n38544;
  assign n38546 = ~n39989 | ~n38562;
  assign n38551 = ~n38549 & ~n38548;
  assign n38550 = ~n39981 | ~n38557;
  assign P1_U3085 = ~n38551 | ~n38550;
  assign n38555 = ~n34150 | ~n38552;
  assign n38554 = ~n40028 | ~n38553;
  assign n38561 = ~n38555 | ~n38554;
  assign n38558 = ~n40025 | ~n38557;
  assign n38564 = ~n38561 & ~n38560;
  assign n38563 = ~n40033 | ~n38562;
  assign P1_U3087 = ~n38564 | ~n38563;
  assign n38568 = ~n39241 & ~n39600;
  assign n38566 = ~n39607 | ~n39244;
  assign n38570 = ~n39602 & ~n39240;
  assign P2_U3080 = ~n38572 | ~n38571;
  assign n38576 = ~n39153 & ~n39600;
  assign n38574 = ~n39607 | ~n39156;
  assign n38578 = ~n39602 & ~n40883;
  assign P2_U3085 = ~n38580 | ~n38579;
  assign n38584 = ~n39268 & ~n39600;
  assign n38582 = ~n39607 | ~n39271;
  assign n38586 = ~n39602 & ~n41318;
  assign P2_U3084 = ~n38588 | ~n38587;
  assign n38591 = ~n42338 & ~n38589;
  assign n38611 = ~n38591 & ~n38590;
  assign n40262 = ~n40202;
  assign n38608 = ~n40262 | ~n38592;
  assign n38606 = ~n41235 & ~n38593;
  assign n38596 = ~n38732 & ~P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n38604 = ~n38596 | ~n40167;
  assign n38601 = ~n38732 | ~n40508;
  assign n40175 = ~n38732 & ~n40384;
  assign n38600 = ~n40175 & ~n41537;
  assign n38597 = n41540 | n40168;
  assign n38599 = ~n38598 | ~n38597;
  assign n38722 = ~n38600 & ~n38599;
  assign n38602 = ~n38601 | ~n38722;
  assign n38603 = ~n38602 | ~P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n38607 = ~n38606 & ~n38605;
  assign P3_U2858 = ~n38611 | ~n38610;
  assign n38624 = ~n41290 & ~n38612;
  assign n38613 = ~n38628 | ~n39522;
  assign n38627 = ~n38626 & ~n39114;
  assign n38622 = ~P2_INSTQUEUE_REG_11__7__SCAN_IN | ~n38938;
  assign n38621 = ~n41284 | ~n38627;
  assign n38633 = ~n39278 & ~n41283;
  assign n38629 = ~n38628 & ~n38627;
  assign n38630 = ~n38629 & ~n39511;
  assign n38632 = ~n41289 & ~n38930;
  assign n38634 = ~n38633 & ~n38632;
  assign P2_U3143 = ~n38635 | ~n38634;
  assign n38637 = ~n43734 & ~n44039;
  assign n38639 = ~n40436 | ~n42942;
  assign P1_U2892 = ~n38640 | ~n38639;
  assign n38646 = ~n38642 & ~n38641;
  assign n38644 = ~n39557 | ~n38646;
  assign n38658 = ~n38644 | ~n38643;
  assign n38656 = ~n38645 & ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n38647 = ~n38646;
  assign n38649 = ~n38648 & ~n38647;
  assign n38651 = ~n38649 & ~n41976;
  assign n38654 = ~n38651 & ~n38650;
  assign n38653 = ~n41979 | ~n38652;
  assign n38655 = ~n38654 | ~n38653;
  assign n39641 = ~n38656 & ~n38655;
  assign n38657 = ~n39641 | ~P1_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n38666 = ~n38658 | ~n38657;
  assign n38663 = n43344 & n38662;
  assign P1_U3019 = ~n38666 | ~n38665;
  assign n38668 = ~n39278 & ~n40895;
  assign n38667 = ~n39280 & ~n38929;
  assign n38675 = ~n38668 & ~n38667;
  assign n38673 = ~n40896 & ~n38930;
  assign n38671 = ~P2_INSTQUEUE_REG_11__3__SCAN_IN | ~n38938;
  assign n38670 = ~n38933 | ~n38669;
  assign P2_U3139 = ~n38675 | ~n38674;
  assign n38677 = ~n39278 & ~n41308;
  assign n38676 = ~n39268 & ~n38929;
  assign n38684 = ~n38677 & ~n38676;
  assign n38682 = ~n41317 & ~n38930;
  assign n38680 = ~P2_INSTQUEUE_REG_11__4__SCAN_IN | ~n38938;
  assign n38679 = ~n38933 | ~n38678;
  assign P2_U3140 = ~n38684 | ~n38683;
  assign n38686 = ~n39278 & ~n40881;
  assign n38685 = ~n39153 & ~n38929;
  assign n38693 = ~n38686 & ~n38685;
  assign n38691 = ~n40882 & ~n38930;
  assign n38689 = ~P2_INSTQUEUE_REG_11__5__SCAN_IN | ~n38938;
  assign n38688 = ~n38933 | ~n38687;
  assign P2_U3141 = ~n38693 | ~n38692;
  assign n38695 = ~n39278 & ~n41295;
  assign n38694 = ~n39200 & ~n38929;
  assign n38702 = ~n38695 & ~n38694;
  assign n38700 = ~n41301 & ~n38930;
  assign n38698 = ~P2_INSTQUEUE_REG_11__6__SCAN_IN | ~n38938;
  assign n38697 = ~n38933 | ~n38696;
  assign P2_U3142 = ~n38702 | ~n38701;
  assign n38705 = ~n39278 & ~n38703;
  assign n38704 = ~n39251 & ~n38929;
  assign n38712 = ~n38705 & ~n38704;
  assign n38710 = ~n39540 & ~n38930;
  assign n38708 = ~P2_INSTQUEUE_REG_11__1__SCAN_IN | ~n38938;
  assign n38707 = ~n38933 | ~n38706;
  assign P2_U3137 = ~n38712 | ~n38711;
  assign n38714 = ~n39278 & ~n40907;
  assign n38713 = ~n39230 & ~n38929;
  assign n38721 = ~n38714 & ~n38713;
  assign n38719 = ~n40908 & ~n38930;
  assign n38717 = ~P2_INSTQUEUE_REG_11__2__SCAN_IN | ~n38938;
  assign n38716 = ~n38933 | ~n38715;
  assign P2_U3138 = ~n38721 | ~n38720;
  assign n38730 = ~n38722 & ~n38732;
  assign n38726 = ~n41235 & ~n38723;
  assign n38725 = ~n40202 & ~n38724;
  assign n38728 = ~n38726 & ~n38725;
  assign n38727 = ~n38732 | ~n40167;
  assign n38729 = ~n38728 | ~n38727;
  assign n38734 = ~n42336 & ~n38731;
  assign n38733 = ~n42338 & ~n38732;
  assign n38736 = ~n38734 & ~n38733;
  assign P3_U2859 = ~n38736 | ~n38735;
  assign n38742 = ~n39280 & ~n38769;
  assign n38738 = ~n41307 & ~n40894;
  assign n38737 = ~n40896 & ~n38770;
  assign n38739 = ~n38773 | ~n39285;
  assign P2_U3163 = ~n38744 | ~n38743;
  assign n38750 = ~n39230 & ~n38769;
  assign n38746 = ~n41307 & ~n40906;
  assign n38745 = ~n40908 & ~n38770;
  assign n38747 = ~n38773 | ~n39233;
  assign P2_U3162 = ~n38752 | ~n38751;
  assign n38758 = ~n39200 & ~n38769;
  assign n38754 = ~n41307 & ~n41302;
  assign n38753 = ~n41301 & ~n38770;
  assign n38755 = ~n38773 | ~n39201;
  assign P2_U3166 = ~n38760 | ~n38759;
  assign n38766 = ~n39601 & ~n38769;
  assign n38762 = ~n41307 & ~n41290;
  assign n38761 = ~n41289 & ~n38770;
  assign n38763 = ~n38773 | ~n39606;
  assign P2_U3167 = ~n38768 | ~n38767;
  assign n38777 = ~n39268 & ~n38769;
  assign n38772 = ~n41307 & ~n41318;
  assign n38771 = ~n41317 & ~n38770;
  assign n38774 = ~n38773 | ~n39271;
  assign P2_U3164 = ~n38780 | ~n38779;
  assign n38782 = ~P1_REIP_REG_10__SCAN_IN | ~n38781;
  assign n38789 = ~n38782 & ~P1_REIP_REG_11__SCAN_IN;
  assign n38784 = ~n39646 | ~n43803;
  assign n38783 = ~n43796 | ~P1_EBX_REG_11__SCAN_IN;
  assign n38785 = ~n38784 | ~n38783;
  assign n38787 = ~n43469 & ~n38785;
  assign n38786 = ~n43797 | ~P1_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n38788 = ~n38787 | ~n38786;
  assign n38797 = ~n38789 & ~n38788;
  assign n38795 = ~n38791 & ~n38790;
  assign n38793 = ~n39592 | ~n43559;
  assign P1_U2829 = ~n38797 | ~n38796;
  assign n38800 = ~n38799 | ~n43462;
  assign n39558 = ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n38805 = ~n43713 & ~n38804;
  assign n38811 = n43469 & P1_REIP_REG_10__SCAN_IN;
  assign n38809 = ~n43709 | ~P1_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign P1_U2989 = ~n38813 | ~n38812;
  assign n38819 = ~n38814 & ~n40350;
  assign n38817 = ~P2_PHYADDRPOINTER_REG_3__SCAN_IN | ~n41921;
  assign n38816 = ~n38815 | ~n40602;
  assign n38818 = ~n38817 | ~n38816;
  assign n38827 = ~n38819 & ~n38818;
  assign n38825 = ~n38820 & ~n41888;
  assign n38823 = ~n38821 | ~n41934;
  assign n38822 = ~n41935 | ~P2_EBX_REG_3__SCAN_IN;
  assign n38824 = ~n38823 | ~n38822;
  assign n38826 = ~n38825 & ~n38824;
  assign n38830 = ~n41204 & ~n38828;
  assign n38831 = n38830 ^ n38829;
  assign n38832 = ~n38831 & ~n41919;
  assign n38834 = ~n23700 | ~n40579;
  assign P2_U2852 = ~n38835 | ~n38834;
  assign n38837 = ~n34135 | ~n38884;
  assign n38836 = ~n39984 | ~n38885;
  assign n38841 = ~n38837 | ~n38836;
  assign n38838 = ~n39981 | ~n38894;
  assign n38842 = ~n39989 | ~n38889;
  assign P1_U3149 = ~n38843 | ~n38842;
  assign n38845 = ~n34165 | ~n38884;
  assign n38844 = ~n39995 | ~n38885;
  assign n38849 = ~n38845 | ~n38844;
  assign n38846 = ~n39992 | ~n38894;
  assign n38850 = ~n40000 | ~n38889;
  assign P1_U3148 = ~n38851 | ~n38850;
  assign n38853 = ~n34188 | ~n38884;
  assign n38852 = ~n39973 | ~n38885;
  assign n38857 = ~n38853 | ~n38852;
  assign n38854 = ~n39978 | ~n38889;
  assign n38858 = ~n39970 | ~n38894;
  assign P1_U3146 = ~n38859 | ~n38858;
  assign n38861 = ~n34227 | ~n38884;
  assign n38860 = ~n40006 | ~n38885;
  assign n38865 = ~n38861 | ~n38860;
  assign n38862 = ~n40011 | ~n38889;
  assign n38866 = ~n40003 | ~n38894;
  assign P1_U3147 = ~n38867 | ~n38866;
  assign n38869 = ~n34072 | ~n38884;
  assign n38868 = ~n40017 | ~n38885;
  assign n38873 = ~n38869 | ~n38868;
  assign n38870 = ~n40022 | ~n38889;
  assign n38874 = ~n40014 | ~n38894;
  assign P1_U3152 = ~n38875 | ~n38874;
  assign n38877 = ~n34150 | ~n38884;
  assign n38876 = ~n40028 | ~n38885;
  assign n38881 = ~n38877 | ~n38876;
  assign n38878 = ~n40033 | ~n38889;
  assign n38882 = ~n40025 | ~n38894;
  assign P1_U3151 = ~n38883 | ~n38882;
  assign n38887 = ~n34098 | ~n38884;
  assign n38886 = ~n40043 | ~n38885;
  assign n38893 = ~n38887 | ~n38886;
  assign n38890 = ~n40049 | ~n38889;
  assign n38895 = ~n40038 | ~n38894;
  assign P1_U3150 = ~n38896 | ~n38895;
  assign n38900 = ~n38898 & ~n35967;
  assign n38899 = ~n43525 & ~P2_EBX_REG_19__SCAN_IN;
  assign P2_U2868 = n38902 | n38901;
  assign n38908 = n40750 | n38903;
  assign n38912 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN & ~P3_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n39427 = ~n38909 & ~n40872;
  assign n38911 = ~n39427 | ~n38910;
  assign n38916 = ~n38912 & ~n38911;
  assign n38914 = ~n38913 | ~n41400;
  assign n40845 = ~n41145 | ~P3_REIP_REG_25__SCAN_IN;
  assign n38915 = ~n38914 | ~n40845;
  assign n38920 = ~n38916 & ~n38915;
  assign n39428 = ~n38918 | ~n38917;
  assign n38919 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN | ~n39428;
  assign n38921 = ~n38920 | ~n38919;
  assign n38926 = ~n41408 & ~n40815;
  assign P3_U2805 = ~n38928 | ~n38927;
  assign n38937 = ~n39241 & ~n38929;
  assign n38932 = ~n39278 & ~n39535;
  assign n38931 = ~n39515 & ~n38930;
  assign n38935 = ~n38932 & ~n38931;
  assign n38934 = ~n38933 | ~n39517;
  assign P2_U3136 = ~n38940 | ~n38939;
  assign n38942 = ~n41176 | ~n38941;
  assign n38943 = ~n41869 | ~n38942;
  assign n38957 = ~n39471 & ~n38943;
  assign n38953 = ~n41172 & ~n41888;
  assign n38944 = ~P2_REIP_REG_8__SCAN_IN | ~n41920;
  assign n38949 = ~n40668 | ~n38944;
  assign n38947 = ~n38945 | ~n41934;
  assign n38946 = ~n39732 | ~n41176;
  assign n38948 = ~n38947 | ~n38946;
  assign n38951 = ~n38949 & ~n38948;
  assign n38950 = ~P2_PHYADDRPOINTER_REG_8__SCAN_IN | ~n41921;
  assign n38952 = ~n38951 | ~n38950;
  assign n38955 = ~n38953 & ~n38952;
  assign n38954 = ~P2_EBX_REG_8__SCAN_IN | ~n41935;
  assign n38958 = ~n41081 | ~n40602;
  assign P2_U2847 = ~n38959 | ~n38958;
  assign n38963 = ~n39280 & ~n39016;
  assign n38961 = ~n39021 | ~n39285;
  assign n38965 = ~n39015 & ~n40894;
  assign n38964 = ~n40896 & ~n39019;
  assign P2_U3067 = ~n38967 | ~n38966;
  assign n38971 = ~BUF2_REG_20__SCAN_IN;
  assign n38976 = ~n42802 & ~n38971;
  assign n38974 = ~n42804 | ~n38972;
  assign n38973 = ~n43698 | ~P2_EAX_REG_20__SCAN_IN;
  assign n38975 = ~n38974 | ~n38973;
  assign n38978 = ~n38976 & ~n38975;
  assign n38977 = ~n43690 | ~BUF1_REG_20__SCAN_IN;
  assign n38979 = ~n38978 | ~n38977;
  assign P2_U2899 = ~n38982 | ~n38981;
  assign n38986 = ~n39268 & ~n39016;
  assign n38984 = ~n39021 | ~n39271;
  assign n38988 = ~n39015 & ~n41318;
  assign n38987 = ~n41317 & ~n39019;
  assign P2_U3068 = ~n38990 | ~n38989;
  assign n38992 = ~n39015 & ~n41290;
  assign n38991 = ~n39601 & ~n39016;
  assign n38998 = ~n38992 & ~n38991;
  assign n38996 = ~n41289 & ~n39019;
  assign n38993 = ~n39021 | ~n39606;
  assign P2_U3071 = ~n38998 | ~n38997;
  assign n39000 = ~n39015 & ~n40883;
  assign n38999 = ~n39153 & ~n39016;
  assign n39006 = ~n39000 & ~n38999;
  assign n39004 = ~n40882 & ~n39019;
  assign n39001 = ~n39021 | ~n39156;
  assign P2_U3069 = ~n39006 | ~n39005;
  assign n39008 = ~n39015 & ~n41302;
  assign n39007 = ~n39200 & ~n39016;
  assign n39014 = ~n39008 & ~n39007;
  assign n39012 = ~n41301 & ~n39019;
  assign n39009 = ~n39021 | ~n39201;
  assign P2_U3070 = ~n39014 | ~n39013;
  assign n39018 = ~n39015 & ~n40906;
  assign n39017 = ~n39230 & ~n39016;
  assign n39027 = ~n39018 & ~n39017;
  assign n39025 = ~n40908 & ~n39019;
  assign n39022 = ~n39021 | ~n39233;
  assign P2_U3066 = ~n39027 | ~n39026;
  assign n39034 = ~n34165 | ~n39097;
  assign n39032 = ~n39956 | ~n39029;
  assign n39031 = ~n39315 | ~n39036;
  assign n39033 = ~n39995 | ~n39098;
  assign n39046 = ~n39034 | ~n39033;
  assign n39043 = ~n39992 | ~n39102;
  assign n39047 = ~n40000 | ~n39107;
  assign P1_U3052 = ~n39048 | ~n39047;
  assign n39050 = ~n34135 | ~n39097;
  assign n39049 = ~n39984 | ~n39098;
  assign n39054 = ~n39050 | ~n39049;
  assign n39051 = ~n39989 | ~n39107;
  assign n39055 = ~n39981 | ~n39102;
  assign P1_U3053 = ~n39056 | ~n39055;
  assign n39058 = ~n34098 | ~n39097;
  assign n39057 = ~n40043 | ~n39098;
  assign n39062 = ~n39058 | ~n39057;
  assign n39059 = ~n40049 | ~n39107;
  assign n39063 = ~n40038 | ~n39102;
  assign P1_U3054 = ~n39064 | ~n39063;
  assign n39066 = ~n34188 | ~n39097;
  assign n39065 = ~n39973 | ~n39098;
  assign n39070 = ~n39066 | ~n39065;
  assign n39067 = ~n39970 | ~n39102;
  assign n39071 = ~n39978 | ~n39107;
  assign P1_U3050 = ~n39072 | ~n39071;
  assign n39074 = ~n34242 | ~n39097;
  assign n39073 = ~n39962 | ~n39098;
  assign n39078 = ~n39074 | ~n39073;
  assign n39075 = ~n39939 | ~n39102;
  assign n39079 = ~n39967 | ~n39107;
  assign P1_U3049 = ~n39080 | ~n39079;
  assign n39082 = ~n34227 | ~n39097;
  assign n39081 = ~n40006 | ~n39098;
  assign n39086 = ~n39082 | ~n39081;
  assign n39083 = ~n40003 | ~n39102;
  assign n39087 = ~n40011 | ~n39107;
  assign P1_U3051 = ~n39088 | ~n39087;
  assign n39090 = ~n34072 | ~n39097;
  assign n39089 = ~n40017 | ~n39098;
  assign n39094 = ~n39090 | ~n39089;
  assign n39091 = ~n40022 | ~n39107;
  assign n39095 = ~n40014 | ~n39102;
  assign P1_U3056 = ~n39096 | ~n39095;
  assign n39100 = ~n34150 | ~n39097;
  assign n39099 = ~n40028 | ~n39098;
  assign n39106 = ~n39100 | ~n39099;
  assign n39103 = ~n40025 | ~n39102;
  assign n39108 = ~n40033 | ~n39107;
  assign P1_U3055 = ~n39109 | ~n39108;
  assign n39115 = ~n39113;
  assign n39117 = ~n39188;
  assign n39116 = ~n39117 & ~n39123;
  assign n39118 = ~n39125 & ~n39117;
  assign n39191 = ~n39120 & ~n39119;
  assign n39122 = ~n39187 & ~n39240;
  assign n39121 = ~n39241 & ~n39188;
  assign n39132 = ~n39122 & ~n39121;
  assign n39128 = n39124 | n39123;
  assign n39131 = ~P2_INSTQUEUE_REG_6__0__SCAN_IN | ~n39192;
  assign n39135 = ~n39193 | ~n39244;
  assign P2_U3096 = ~n39136 | ~n39135;
  assign n39138 = ~n39187 & ~n41318;
  assign n39137 = ~n39268 & ~n39188;
  assign n39144 = ~n39138 & ~n39137;
  assign n39140 = ~P2_INSTQUEUE_REG_6__4__SCAN_IN | ~n39192;
  assign P2_U3100 = ~n39144 | ~n39143;
  assign n39146 = ~n39187 & ~n39549;
  assign n39145 = ~n39251 & ~n39188;
  assign n39152 = ~n39146 & ~n39145;
  assign n39148 = ~P2_INSTQUEUE_REG_6__1__SCAN_IN | ~n39192;
  assign P2_U3097 = ~n39152 | ~n39151;
  assign n39155 = ~n39187 & ~n40883;
  assign n39154 = ~n39153 & ~n39188;
  assign n39162 = ~n39155 & ~n39154;
  assign n39160 = ~n40882 & ~n39191;
  assign n39158 = ~P2_INSTQUEUE_REG_6__5__SCAN_IN | ~n39192;
  assign P2_U3101 = ~n39162 | ~n39161;
  assign n39164 = ~n39187 & ~n40894;
  assign n39163 = ~n39280 & ~n39188;
  assign n39170 = ~n39164 & ~n39163;
  assign n39166 = ~P2_INSTQUEUE_REG_6__3__SCAN_IN | ~n39192;
  assign P2_U3099 = ~n39170 | ~n39169;
  assign n39172 = ~n39187 & ~n40906;
  assign n39171 = ~n39230 & ~n39188;
  assign n39178 = ~n39172 & ~n39171;
  assign n39174 = ~P2_INSTQUEUE_REG_6__2__SCAN_IN | ~n39192;
  assign P2_U3098 = ~n39178 | ~n39177;
  assign n39180 = ~n39187 & ~n41302;
  assign n39179 = ~n39200 & ~n39188;
  assign n39186 = ~n39180 & ~n39179;
  assign n39182 = ~P2_INSTQUEUE_REG_6__6__SCAN_IN | ~n39192;
  assign P2_U3102 = ~n39186 | ~n39185;
  assign n39190 = ~n39187 & ~n41290;
  assign n39189 = ~n39601 & ~n39188;
  assign n39199 = ~n39190 & ~n39189;
  assign n39195 = ~P2_INSTQUEUE_REG_6__7__SCAN_IN | ~n39192;
  assign P2_U3103 = ~n39199 | ~n39198;
  assign n39205 = ~n39200 & ~n39279;
  assign n39207 = ~n39278 & ~n41302;
  assign n39206 = ~n41301 & ~n39283;
  assign P2_U3134 = ~n39209 | ~n39208;
  assign n39213 = ~n42256 | ~n41934;
  assign n39212 = ~n41935 | ~P2_EBX_REG_17__SCAN_IN;
  assign n39215 = ~n39213 | ~n39212;
  assign n39214 = ~n42260 & ~n41926;
  assign n39216 = ~n39215 & ~n39214;
  assign n39220 = ~n39216 | ~n40668;
  assign n39218 = ~n41920 | ~P2_REIP_REG_17__SCAN_IN;
  assign n39217 = ~n41921 | ~P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n39219 = ~n39218 | ~n39217;
  assign n39229 = ~n39220 & ~n39219;
  assign n39227 = ~n42612 & ~n41931;
  assign n39225 = ~n42616 | ~n41942;
  assign n39221 = ~n42260 & ~n40624;
  assign n39223 = ~n39221 & ~n40669;
  assign n39224 = ~n39223 | ~n39222;
  assign n39226 = ~n39225 | ~n39224;
  assign P2_U2838 = ~n39229 | ~n39228;
  assign n39232 = ~n39278 & ~n40906;
  assign n39231 = ~n39230 & ~n39279;
  assign n39239 = ~n39232 & ~n39231;
  assign n39237 = ~n40908 & ~n39283;
  assign n39234 = ~n39286 | ~n39233;
  assign P2_U3130 = ~n39239 | ~n39238;
  assign n39243 = ~n39278 & ~n39240;
  assign n39242 = ~n39241 & ~n39279;
  assign n39250 = ~n39243 & ~n39242;
  assign n39248 = ~n39515 & ~n39283;
  assign n39245 = ~n39286 | ~n39244;
  assign P2_U3128 = ~n39250 | ~n39249;
  assign n39253 = ~n39278 & ~n39549;
  assign n39252 = ~n39251 & ~n39279;
  assign n39259 = ~n39253 & ~n39252;
  assign n39257 = ~n39540 & ~n39283;
  assign n39254 = ~n39286 | ~n39542;
  assign P2_U3129 = ~n39259 | ~n39258;
  assign n39261 = ~n39278 & ~n41290;
  assign n39260 = ~n39601 & ~n39279;
  assign n39267 = ~n39261 & ~n39260;
  assign n39265 = ~n41289 & ~n39283;
  assign n39262 = ~n39286 | ~n39606;
  assign P2_U3135 = ~n39267 | ~n39266;
  assign n39270 = ~n39278 & ~n41318;
  assign n39269 = ~n39268 & ~n39279;
  assign n39277 = ~n39270 & ~n39269;
  assign n39275 = ~n41317 & ~n39283;
  assign n39272 = ~n39286 | ~n39271;
  assign P2_U3132 = ~n39277 | ~n39276;
  assign n39282 = ~n39278 & ~n40894;
  assign n39281 = ~n39280 & ~n39279;
  assign n39292 = ~n39282 & ~n39281;
  assign n39290 = ~n40896 & ~n39283;
  assign n39287 = ~n39286 | ~n39285;
  assign P2_U3131 = ~n39292 | ~n39291;
  assign n39294 = n43525 | P2_EBX_REG_20__SCAN_IN;
  assign P2_U2867 = ~n39297 | ~n39296;
  assign n39373 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n39298;
  assign n39300 = ~n34072 | ~n39373;
  assign n39299 = ~n40014 | ~n39374;
  assign n39322 = ~n39300 | ~n39299;
  assign n39306 = ~n39302 & ~n39301;
  assign n39305 = n39946 | n39304;
  assign n39308 = ~n39307 & ~n39373;
  assign n39314 = ~n39311 | ~n39310;
  assign n39816 = n39314 & P1_STATE2_REG_2__SCAN_IN;
  assign n39312 = ~n39816 & ~n39953;
  assign n39820 = ~n39314;
  assign n39318 = ~n39820 | ~n39956;
  assign n39317 = ~n39316 | ~n39958;
  assign n39319 = ~n40017 | ~n39378;
  assign n39323 = ~n40022 | ~n39383;
  assign P1_U3104 = ~n39324 | ~n39323;
  assign n39326 = ~n34242 | ~n39373;
  assign n39325 = ~n39939 | ~n39374;
  assign n39330 = ~n39326 | ~n39325;
  assign n39327 = ~n39962 | ~n39378;
  assign n39331 = ~n39967 | ~n39383;
  assign P1_U3097 = ~n39332 | ~n39331;
  assign n39334 = ~n34165 | ~n39373;
  assign n39333 = ~n39992 | ~n39374;
  assign n39338 = ~n39334 | ~n39333;
  assign n39335 = ~n39995 | ~n39378;
  assign n39339 = ~n40000 | ~n39383;
  assign P1_U3100 = ~n39340 | ~n39339;
  assign n39342 = ~n34227 | ~n39373;
  assign n39341 = ~n40003 | ~n39374;
  assign n39346 = ~n39342 | ~n39341;
  assign n39343 = ~n40006 | ~n39378;
  assign n39347 = ~n40011 | ~n39383;
  assign P1_U3099 = ~n39348 | ~n39347;
  assign n39350 = ~n34135 | ~n39373;
  assign n39349 = ~n39981 | ~n39374;
  assign n39354 = ~n39350 | ~n39349;
  assign n39351 = ~n39984 | ~n39378;
  assign n39355 = ~n39989 | ~n39383;
  assign P1_U3101 = ~n39356 | ~n39355;
  assign n39358 = ~n34188 | ~n39373;
  assign n39357 = ~n39970 | ~n39374;
  assign n39362 = ~n39358 | ~n39357;
  assign n39359 = ~n39973 | ~n39378;
  assign n39363 = ~n39978 | ~n39383;
  assign P1_U3098 = ~n39364 | ~n39363;
  assign n39366 = ~n34098 | ~n39373;
  assign n39365 = ~n40038 | ~n39374;
  assign n39370 = ~n39366 | ~n39365;
  assign n39367 = ~n40043 | ~n39378;
  assign n39371 = ~n40049 | ~n39383;
  assign P1_U3102 = ~n39372 | ~n39371;
  assign n39376 = ~n34150 | ~n39373;
  assign n39375 = ~n40025 | ~n39374;
  assign n39382 = ~n39376 | ~n39375;
  assign n39379 = ~n40028 | ~n39378;
  assign n39384 = ~n40033 | ~n39383;
  assign P1_U3103 = ~n39385 | ~n39384;
  assign n40222 = ~n40132 & ~n39386;
  assign n40212 = ~n40422 | ~n40222;
  assign n39391 = ~n40339 & ~n40212;
  assign n39403 = ~n39440 & ~n40415;
  assign n39402 = ~n39394 & ~n41240;
  assign n39406 = n40221 & P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n39397 = ~n42322 & ~n39406;
  assign n39396 = ~n41235 & ~n39395;
  assign n39400 = ~n39397 & ~n39396;
  assign n40126 = ~n41540 & ~n39405;
  assign n39399 = ~n40418 & ~n39398;
  assign n40124 = ~n39399 & ~n41537;
  assign n40226 = ~n40126 & ~n40124;
  assign n39407 = ~n40210 | ~n39406;
  assign n39408 = ~n39440 | ~n39407;
  assign n39416 = ~n42338 & ~n39440;
  assign P3_U2845 = ~n39419 | ~n39418;
  assign n41017 = ~n41145 | ~P3_REIP_REG_24__SCAN_IN;
  assign n39436 = ~n41017;
  assign n39421 = ~n41149 ^ P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n39432 = ~n39425 & ~n41520;
  assign n39430 = ~n39427 | ~n39426;
  assign n39429 = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN | ~n39428;
  assign n39431 = ~n39430 | ~n39429;
  assign n39433 = ~n39432 & ~n39431;
  assign P3_U2806 = ~n39439 | ~n39438;
  assign n39458 = ~n42338 & ~n40421;
  assign n39441 = n39440 | n40415;
  assign n39443 = ~n39441 | ~n41005;
  assign P3_U2844 = ~n39460 | ~n39459;
  assign n39463 = n39461 | n39482;
  assign n39462 = ~n41935 | ~P2_EBX_REG_9__SCAN_IN;
  assign n39465 = ~n39463 | ~n39462;
  assign n39464 = ~n41504 & ~n41926;
  assign n39466 = ~n39465 & ~n39464;
  assign n39468 = ~n41920 | ~P2_REIP_REG_9__SCAN_IN;
  assign n39467 = ~n41921 | ~P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n39469 = ~n39468 | ~n39467;
  assign n39479 = ~n39470 & ~n39469;
  assign n39477 = ~n41703 & ~n41931;
  assign n39475 = ~n41707 | ~n41942;
  assign n39472 = ~n41504 & ~n39471;
  assign n39473 = ~n39472 & ~n40669;
  assign n39474 = ~n39473 | ~n40293;
  assign n39476 = ~n39475 | ~n39474;
  assign n39478 = ~n39477 & ~n39476;
  assign P2_U2846 = ~n39479 | ~n39478;
  assign n39484 = n42066 | n39482;
  assign n39483 = ~n41935 | ~P2_EBX_REG_11__SCAN_IN;
  assign n39486 = ~n39484 | ~n39483;
  assign n39485 = ~n42061 & ~n41926;
  assign n39487 = ~n39486 & ~n39485;
  assign n39489 = ~n41920 | ~P2_REIP_REG_11__SCAN_IN;
  assign n39488 = ~n41921 | ~P2_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n39490 = ~n39489 | ~n39488;
  assign n39499 = ~n39491 & ~n39490;
  assign n39497 = ~n42568 & ~n41931;
  assign n39495 = ~n42565 | ~n41942;
  assign n39492 = ~n42061 & ~n40296;
  assign n39493 = ~n39492 & ~n40669;
  assign n39494 = ~n39493 | ~n40647;
  assign n39496 = ~n39495 | ~n39494;
  assign n39498 = ~n39497 & ~n39496;
  assign P2_U2844 = ~n39499 | ~n39498;
  assign n39506 = ~n42135 | ~n39500;
  assign n39501 = ~P3_EBX_REG_22__SCAN_IN | ~n43930;
  assign P3_U2681 = ~n39506 | ~n39505;
  assign n39512 = ~n39523 & ~n41310;
  assign n39513 = ~n39512 & ~n39511;
  assign n39521 = ~n39515 & ~n41316;
  assign n39519 = ~n39516 | ~n41310;
  assign n39518 = ~n39548 | ~n39517;
  assign n39520 = ~n39519 | ~n39518;
  assign n39539 = ~n39521 & ~n39520;
  assign n39533 = ~n41310 & ~n39526;
  assign n39537 = ~n40891 & ~n39534;
  assign n39536 = ~n39535 & ~n41307;
  assign n39538 = ~n39537 & ~n39536;
  assign P2_U3168 = ~n39539 | ~n39538;
  assign n39547 = ~n39540 & ~n41316;
  assign n39545 = ~n39541 | ~n41310;
  assign n39544 = ~n39543 | ~n39542;
  assign n39546 = ~n39545 | ~n39544;
  assign n39553 = ~n39547 & ~n39546;
  assign n39551 = ~n40891 & ~n41578;
  assign n39550 = ~n39549 & ~n41319;
  assign n39552 = ~n39551 & ~n39550;
  assign P2_U3169 = ~n39553 | ~n39552;
  assign n39554 = ~P1_INSTADDRPOINTER_REG_10__SCAN_IN & ~P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n39556 = ~n39555 & ~n39554;
  assign n39568 = ~n39557 | ~n39556;
  assign n39566 = ~n39559 & ~n39558;
  assign n39561 = ~n43469 | ~P1_REIP_REG_10__SCAN_IN;
  assign P1_U3021 = ~n39568 | ~n39567;
  assign n39570 = ~n39569;
  assign n39582 = ~n39571 & ~n39570;
  assign n39572 = ~P2_REIP_REG_31__SCAN_IN;
  assign n39577 = ~n28361 & ~n39572;
  assign n39575 = ~n39573 | ~P2_EBX_REG_31__SCAN_IN;
  assign n39574 = ~P2_PHYADDRPOINTER_REG_31__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n39576 = ~n39575 | ~n39574;
  assign n39580 = ~n39577 & ~n39576;
  assign n39579 = ~n39578 | ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n39581 = ~n39580 | ~n39579;
  assign n39584 = ~n35967 | ~P2_EBX_REG_31__SCAN_IN;
  assign P2_U2856 = ~n39585 | ~n39584;
  assign n39644 = ~n43469 | ~P1_REIP_REG_11__SCAN_IN;
  assign n39591 = ~n43709 | ~P1_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n39597 = ~n39644 | ~n39591;
  assign n39595 = ~n43362 | ~n39592;
  assign P1_U2988 = ~n39599 | ~n39598;
  assign n39611 = ~n39601 & ~n39600;
  assign n39605 = ~n39602 & ~n41290;
  assign n39604 = ~n41289 & ~n39603;
  assign n39608 = ~n39607 | ~n39606;
  assign P2_U3087 = ~n39614 | ~n39613;
  assign n39637 = ~n42338 & ~n39620;
  assign n39617 = ~n39616 ^ n39615;
  assign n39634 = ~n39617 & ~n40202;
  assign n39632 = ~n41542 | ~n39618;
  assign n39619 = ~n39624;
  assign n39621 = ~n39619 | ~n40167;
  assign n39630 = ~n39621 | ~n39620;
  assign n39623 = ~n39622 | ~n40170;
  assign n39628 = ~n39623 | ~n40422;
  assign n39625 = ~n39624 & ~n40384;
  assign n40444 = ~n39625 & ~n41537;
  assign n40267 = ~n40444 & ~n40260;
  assign n39626 = ~n40125 & ~n40267;
  assign n40505 = ~n40968 | ~n40389;
  assign n40446 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN | ~n40505;
  assign n39627 = ~n39626 & ~n40446;
  assign n39629 = ~n39628 | ~n39627;
  assign n39639 = ~n39637 & ~n39636;
  assign P3_U2854 = ~n39639 | ~n39638;
  assign n39642 = ~n39640 & ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n39650 = n39642 | n39641;
  assign n39647 = n43344 & n39646;
  assign P1_U3020 = ~n39650 | ~n39649;
  assign n39666 = ~n40770 & ~n39651;
  assign n39662 = ~n39652 & ~n43755;
  assign n39655 = ~n43877 & ~n40354;
  assign n39654 = ~n39653;
  assign n39660 = ~n39655 & ~n39654;
  assign n39657 = ~P2_INSTADDRPOINTER_REG_5__SCAN_IN & ~n39656;
  assign n39659 = ~n39658 | ~n39657;
  assign n39661 = ~n39660 | ~n39659;
  assign n39664 = ~n39662 & ~n39661;
  assign n39663 = ~n43767 | ~n40368;
  assign P2_U3041 = ~n39669 | ~n39668;
  assign n39674 = ~BUF2_REG_21__SCAN_IN;
  assign n39679 = ~n42802 & ~n39674;
  assign n39677 = ~n42804 | ~n39675;
  assign n39676 = ~n43698 | ~P2_EAX_REG_21__SCAN_IN;
  assign n39678 = ~n39677 | ~n39676;
  assign n39681 = ~n39679 & ~n39678;
  assign n39680 = ~n43690 | ~BUF1_REG_21__SCAN_IN;
  assign n39682 = ~n39681 | ~n39680;
  assign P2_U2898 = ~n39685 | ~n39684;
  assign n39687 = ~n40436 | ~n43121;
  assign n39686 = ~P1_EAX_REG_13__SCAN_IN | ~n43732;
  assign n39690 = n39687 & n39686;
  assign P1_U2891 = ~n39690 | ~n39689;
  assign n39692 = ~n41920 | ~P2_REIP_REG_22__SCAN_IN;
  assign n39691 = ~n41921 | ~P2_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n39697 = ~n39692 | ~n39691;
  assign n39694 = ~n39693 | ~n41718;
  assign n39695 = n39694 ^ n43000;
  assign n39696 = ~n39695 & ~n41919;
  assign n39699 = ~n39697 & ~n39696;
  assign n39698 = ~P2_EBX_REG_22__SCAN_IN | ~n41935;
  assign n39706 = ~n43016 | ~n40602;
  assign n39705 = ~n39704 | ~n41942;
  assign n39711 = ~n42899 | ~n41934;
  assign P2_U2833 = ~n39712 | ~n39711;
  assign n39714 = n43525 | P2_EBX_REG_21__SCAN_IN;
  assign P2_U2866 = ~n39717 | ~n39716;
  assign n39720 = ~n40350 & ~n26537;
  assign n39718 = ~P2_PHYADDRPOINTER_REG_6__SCAN_IN | ~n41921;
  assign n39719 = ~n39718 | ~n40668;
  assign n39726 = ~n39720 & ~n39719;
  assign n39724 = ~n39721 & ~n40669;
  assign n39723 = ~n40157 | ~n39722;
  assign n39725 = ~n39724 | ~n39723;
  assign n39729 = ~n39726 | ~n39725;
  assign n39728 = n39727 & n41934;
  assign n39731 = ~n39729 & ~n39728;
  assign n39730 = ~P2_EBX_REG_6__SCAN_IN | ~n41935;
  assign n39736 = ~n39731 | ~n39730;
  assign n39734 = ~n39732 | ~n40157;
  assign n39733 = ~n40154 | ~n41942;
  assign n39735 = ~n39734 | ~n39733;
  assign n39739 = ~n39736 & ~n39735;
  assign n39738 = n39737 | n41931;
  assign P2_U2849 = ~n39739 | ~n39738;
  assign n39746 = ~n42135 | ~n39740;
  assign n39742 = ~P3_EBX_REG_23__SCAN_IN | ~n43930;
  assign P3_U2680 = ~n39746 | ~n39745;
  assign n39748 = ~n41920 | ~P2_REIP_REG_24__SCAN_IN;
  assign n39747 = ~n41921 | ~P2_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n39755 = ~n39748 | ~n39747;
  assign n39750 = ~n39749 | ~n41718;
  assign n39751 = ~n39750 ^ n43217;
  assign n39753 = ~n39751 | ~n41206;
  assign n39752 = ~P2_EBX_REG_24__SCAN_IN | ~n41935;
  assign n39760 = ~n39759;
  assign n43225 = ~n39910 & ~n39762;
  assign n39766 = ~n43225 | ~n40602;
  assign P2_U2831 = ~n39770 | ~n39769;
  assign n39778 = ~n39775 | ~n40823;
  assign n39777 = ~n39776 | ~n42320;
  assign n39779 = ~n39778 | ~n39777;
  assign n40240 = n40999 | n39779;
  assign n40523 = n41540 | n39780;
  assign n39781 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN | ~n40523;
  assign n39784 = ~n39781 | ~n40508;
  assign n40821 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~n40243;
  assign n39782 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~n41537;
  assign n39783 = ~n40821 | ~n39782;
  assign n39793 = ~n39784 | ~n39783;
  assign n39787 = ~n40422 | ~n39786;
  assign n39791 = ~n41546 | ~n39790;
  assign n39800 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n39801 = ~n42338 & ~n39800;
  assign P3_U2840 = ~n39804 | ~n39803;
  assign n39878 = n39805 & n39937;
  assign n39807 = ~n34135 | ~n39878;
  assign n39806 = ~n39989 | ~n39879;
  assign n39827 = ~n39807 | ~n39806;
  assign n39812 = ~n39878;
  assign n39813 = ~n39812 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n39823 = ~n39820 | ~n39819;
  assign n39822 = ~n39821 | ~n39958;
  assign n39824 = ~n39984 | ~n39883;
  assign n39828 = ~n39981 | ~n39888;
  assign P1_U3133 = ~n39829 | ~n39828;
  assign n39831 = ~n34227 | ~n39878;
  assign n39830 = ~n40011 | ~n39879;
  assign n39835 = ~n39831 | ~n39830;
  assign n39832 = ~n40006 | ~n39883;
  assign n39836 = ~n40003 | ~n39888;
  assign P1_U3131 = ~n39837 | ~n39836;
  assign n39839 = ~n34072 | ~n39878;
  assign n39838 = ~n40022 | ~n39879;
  assign n39843 = ~n39839 | ~n39838;
  assign n39840 = ~n40017 | ~n39883;
  assign n39844 = ~n40014 | ~n39888;
  assign P1_U3136 = ~n39845 | ~n39844;
  assign n39847 = ~n34098 | ~n39878;
  assign n39846 = ~n40049 | ~n39879;
  assign n39851 = ~n39847 | ~n39846;
  assign n39848 = ~n40043 | ~n39883;
  assign n39852 = ~n40038 | ~n39888;
  assign P1_U3134 = ~n39853 | ~n39852;
  assign n39855 = ~n34150 | ~n39878;
  assign n39854 = ~n40033 | ~n39879;
  assign n39859 = ~n39855 | ~n39854;
  assign n39856 = ~n40028 | ~n39883;
  assign n39860 = ~n40025 | ~n39888;
  assign P1_U3135 = ~n39861 | ~n39860;
  assign n39863 = ~n34188 | ~n39878;
  assign n39862 = ~n39978 | ~n39879;
  assign n39867 = ~n39863 | ~n39862;
  assign n39864 = ~n39973 | ~n39883;
  assign n39868 = ~n39970 | ~n39888;
  assign P1_U3130 = ~n39869 | ~n39868;
  assign n39871 = ~n34242 | ~n39878;
  assign n39870 = ~n39967 | ~n39879;
  assign n39875 = ~n39871 | ~n39870;
  assign n39872 = ~n39962 | ~n39883;
  assign n39876 = ~n39939 | ~n39888;
  assign P1_U3129 = ~n39877 | ~n39876;
  assign n39881 = ~n34165 | ~n39878;
  assign n39880 = ~n40000 | ~n39879;
  assign n39887 = ~n39881 | ~n39880;
  assign n39884 = ~n39995 | ~n39883;
  assign n39889 = ~n39992 | ~n39888;
  assign P1_U3132 = ~n39890 | ~n39889;
  assign n39893 = ~n39892 & ~n39891;
  assign n39899 = ~n43306 | ~n39894;
  assign n39900 = ~n39895;
  assign n39897 = ~n39896 & ~n39900;
  assign n39898 = ~n43737 | ~BUF1_REG_16__SCAN_IN;
  assign n39906 = ~n39899 | ~n39898;
  assign n39902 = ~n39901 & ~n39900;
  assign n39904 = ~n43738 | ~DATAI_16_;
  assign n39903 = ~n43732 | ~P1_EAX_REG_16__SCAN_IN;
  assign n39905 = ~n39904 | ~n39903;
  assign n39908 = ~n39906 & ~n39905;
  assign P1_U2888 = ~n39908 | ~n39907;
  assign n39912 = ~n41920 | ~P2_REIP_REG_25__SCAN_IN;
  assign n39911 = ~n41921 | ~P2_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n39919 = ~n39912 | ~n39911;
  assign n39914 = ~n41204 & ~n39913;
  assign n39915 = ~n39914 ^ n43546;
  assign n39917 = ~n39915 | ~n41206;
  assign n39916 = ~P2_EBX_REG_25__SCAN_IN | ~n41935;
  assign n39918 = ~n39917 | ~n39916;
  assign n39924 = ~n39919 & ~n39918;
  assign n39923 = ~n39922 | ~n41942;
  assign P2_U2830 = ~n39930 | ~n39929;
  assign n39933 = ~n40436 | ~n39931;
  assign n39932 = ~n43732 | ~P1_EAX_REG_15__SCAN_IN;
  assign P1_U2889 = n39936 | n39935;
  assign n39949 = ~n39938 | ~n39937;
  assign n40036 = ~n39949;
  assign n39941 = ~n34242 | ~n40036;
  assign n39940 = ~n39939 | ~n40037;
  assign n39966 = ~n39941 | ~n39940;
  assign n39950 = ~n39949 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n39961 = ~n39957 | ~n39956;
  assign n39960 = ~n39959 | ~n39958;
  assign n39963 = ~n39962 | ~n40042;
  assign n39968 = ~n39967 | ~n40048;
  assign P1_U3033 = ~n39969 | ~n39968;
  assign n39972 = ~n34188 | ~n40036;
  assign n39971 = ~n39970 | ~n40037;
  assign n39977 = ~n39972 | ~n39971;
  assign n39974 = ~n39973 | ~n40042;
  assign n39979 = ~n39978 | ~n40048;
  assign P1_U3034 = ~n39980 | ~n39979;
  assign n39983 = ~n34135 | ~n40036;
  assign n39982 = ~n39981 | ~n40037;
  assign n39988 = ~n39983 | ~n39982;
  assign n39985 = ~n39984 | ~n40042;
  assign n39990 = ~n39989 | ~n40048;
  assign P1_U3037 = ~n39991 | ~n39990;
  assign n39994 = ~n34165 | ~n40036;
  assign n39993 = ~n39992 | ~n40037;
  assign n39999 = ~n39994 | ~n39993;
  assign n39996 = ~n39995 | ~n40042;
  assign n40001 = ~n40000 | ~n40048;
  assign P1_U3036 = ~n40002 | ~n40001;
  assign n40005 = ~n34227 | ~n40036;
  assign n40004 = ~n40003 | ~n40037;
  assign n40010 = ~n40005 | ~n40004;
  assign n40007 = ~n40006 | ~n40042;
  assign n40012 = ~n40011 | ~n40048;
  assign P1_U3035 = ~n40013 | ~n40012;
  assign n40016 = ~n34072 | ~n40036;
  assign n40015 = ~n40014 | ~n40037;
  assign n40021 = ~n40016 | ~n40015;
  assign n40018 = ~n40017 | ~n40042;
  assign n40023 = ~n40022 | ~n40048;
  assign P1_U3040 = ~n40024 | ~n40023;
  assign n40027 = ~n34150 | ~n40036;
  assign n40026 = ~n40025 | ~n40037;
  assign n40032 = ~n40027 | ~n40026;
  assign n40029 = ~n40028 | ~n40042;
  assign n40034 = ~n40033 | ~n40048;
  assign P1_U3039 = ~n40035 | ~n40034;
  assign n40040 = ~n34098 | ~n40036;
  assign n40039 = ~n40038 | ~n40037;
  assign n40047 = ~n40040 | ~n40039;
  assign n40044 = ~n40043 | ~n40042;
  assign n40050 = ~n40049 | ~n40048;
  assign P1_U3038 = ~n40051 | ~n40050;
  assign n40060 = ~n42802 & ~n40055;
  assign n40058 = ~n42804 | ~n40056;
  assign n40057 = ~n43698 | ~P2_EAX_REG_22__SCAN_IN;
  assign n40059 = ~n40058 | ~n40057;
  assign n40062 = ~n40060 & ~n40059;
  assign n40061 = ~n43690 | ~BUF1_REG_22__SCAN_IN;
  assign n40063 = ~n40062 | ~n40061;
  assign P2_U2897 = ~n40066 | ~n40065;
  assign n40068 = n43525 | P2_EBX_REG_22__SCAN_IN;
  assign P2_U2865 = ~n40071 | ~n40070;
  assign n40087 = ~P1_EBX_REG_31__SCAN_IN | ~n44023;
  assign n40077 = ~n42979 & ~n40072;
  assign n40075 = ~n40080 | ~P1_EBX_REG_30__SCAN_IN;
  assign n40074 = ~n40081 | ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n42982 = ~n40075 | ~n40074;
  assign n40076 = ~n42982;
  assign n40083 = ~n40080 | ~P1_EBX_REG_31__SCAN_IN;
  assign n40082 = ~n40081 | ~P1_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n40084 = ~n40083 | ~n40082;
  assign P1_U2841 = ~n40087 | ~n40086;
  assign n40090 = ~P1_INSTADDRPOINTER_REG_13__SCAN_IN & ~n40088;
  assign n40487 = ~n43033 & ~n40089;
  assign n40104 = ~n40090 & ~n40487;
  assign n40102 = ~n40092 & ~n40091;
  assign n40095 = ~n40093;
  assign P1_U3018 = ~n40104 | ~n40103;
  assign n40106 = ~n41920 | ~P2_REIP_REG_23__SCAN_IN;
  assign n40105 = ~n41921 | ~P2_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n40111 = ~n40106 | ~n40105;
  assign n40108 = ~n41204 & ~n40107;
  assign n40109 = n40108 ^ n42960;
  assign n40110 = ~n40109 & ~n41919;
  assign n40113 = ~n40111 & ~n40110;
  assign n40112 = ~P2_EBX_REG_23__SCAN_IN | ~n41935;
  assign n40117 = ~n42909 | ~n40602;
  assign n40116 = ~n41265 | ~n41942;
  assign n40122 = ~n42904 | ~n41934;
  assign P2_U2832 = ~n40123 | ~n40122;
  assign n40149 = ~n42338 & ~n40132;
  assign n40965 = ~n40962 & ~n40124;
  assign n40131 = ~n40965 & ~n40125;
  assign n40967 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN & ~n40442;
  assign n40129 = ~n40126 & ~n40967;
  assign n40128 = ~n40127 | ~n40443;
  assign n40393 = ~n40422 | ~n40128;
  assign n40130 = ~n40129 | ~n40393;
  assign n40133 = ~n40131 & ~n40130;
  assign n40139 = ~n40133 & ~n40132;
  assign n40137 = ~n40134 | ~n40980;
  assign n40136 = ~n40135 | ~n41542;
  assign n40138 = ~n40137 | ~n40136;
  assign n40143 = ~n40139 & ~n40138;
  assign n40140 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN & ~n40373;
  assign n40145 = ~n40144 & ~n41240;
  assign P3_U2848 = ~n40151 | ~n40150;
  assign n40165 = ~n40152 & ~n43924;
  assign n40163 = ~n40153 | ~n43913;
  assign n40156 = ~n43813 | ~n40154;
  assign n40155 = ~n43917 | ~P2_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n40161 = ~n40156 | ~n40155;
  assign n40158 = ~n43896 | ~n40157;
  assign n40160 = ~n40159 | ~n40158;
  assign n40162 = ~n40161 & ~n40160;
  assign P2_U3008 = n40165 | n40164;
  assign n40188 = ~n42338 & ~n40191;
  assign n40171 = ~n40166;
  assign n40169 = ~n40171 | ~n40168;
  assign n40174 = ~n40169 | ~n40968;
  assign n40172 = ~n40171 | ~n40170;
  assign n40173 = ~n40422 | ~n40172;
  assign n40178 = ~n40191 & ~n40269;
  assign n40176 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN | ~n40175;
  assign n40177 = ~n40176 | ~n42320;
  assign n40181 = ~n41542 | ~n40180;
  assign n40184 = ~n40202 & ~n40183;
  assign n40187 = ~n42336 & ~n40186;
  assign n40190 = ~n40188 & ~n40187;
  assign P3_U2857 = ~n40190 | ~n40189;
  assign n40207 = ~n42338 & ~n40196;
  assign n40192 = ~n40270 & ~n40191;
  assign n40198 = ~n41235 & ~n40193;
  assign n40195 = ~n41005 | ~n40194;
  assign n40197 = ~n40196 & ~n40195;
  assign n40199 = ~n40198 & ~n40197;
  assign n40203 = ~n40202 & ~n40201;
  assign n40206 = ~n42336 & ~n40205;
  assign n40209 = ~n40207 & ~n40206;
  assign P3_U2856 = ~n40209 | ~n40208;
  assign n40338 = n40212 & n40211;
  assign n40220 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN & ~n40338;
  assign n40329 = ~n40213 & ~n41240;
  assign n40218 = ~n40329 | ~n40214;
  assign n40330 = ~n40215 & ~n41235;
  assign n40217 = ~n40330 | ~n40216;
  assign n40219 = ~n40218 | ~n40217;
  assign n40228 = ~n40220 & ~n40219;
  assign n40224 = ~n40221 & ~n42322;
  assign n40223 = ~n40442 & ~n40222;
  assign n40225 = ~n40224 & ~n40223;
  assign n40227 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN | ~n40331;
  assign n40230 = ~n40229 & ~n42318;
  assign n40233 = ~n42338 & ~n40339;
  assign P3_U2847 = ~n40236 | ~n40235;
  assign n40238 = ~n40820 & ~n42338;
  assign n40259 = ~n40238 & ~n40237;
  assign n40250 = ~n40242 & ~n41240;
  assign n40246 = ~n40243 & ~n42322;
  assign n40832 = ~n40422 | ~n40251;
  assign n41004 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~n40832;
  assign n40252 = ~n41004;
  assign P3_U2839 = ~n40259 | ~n40258;
  assign n40279 = ~n42338 & ~n40260;
  assign n40265 = ~n40261 | ~n41542;
  assign n40264 = ~n40263 | ~n40262;
  assign n40276 = ~n40265 | ~n40264;
  assign n40266 = ~n40508 | ~n40271;
  assign n40268 = ~n40267 | ~n40266;
  assign n40274 = ~n40269 & ~n40268;
  assign n40272 = ~n40271 & ~n40270;
  assign n40273 = ~n40272 & ~P3_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n40281 = ~n40279 & ~n40278;
  assign P3_U2855 = ~n40281 | ~n40280;
  assign n40284 = ~n40282 | ~n41934;
  assign n40283 = ~n41935 | ~P2_EBX_REG_10__SCAN_IN;
  assign n40287 = ~n40284 | ~n40283;
  assign n40286 = ~n40285 & ~n41926;
  assign n40288 = ~n40287 & ~n40286;
  assign n40292 = ~n40288 | ~n40668;
  assign n40290 = ~n41920 | ~P2_REIP_REG_10__SCAN_IN;
  assign n40289 = ~n41921 | ~P2_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n40291 = ~n40290 | ~n40289;
  assign n40305 = ~n40292 & ~n40291;
  assign n40295 = ~n40294 | ~n40293;
  assign n40297 = ~n41869 | ~n40295;
  assign n40303 = ~n40297 & ~n40296;
  assign n40301 = n40298 | n41931;
  assign n40300 = ~n40299 | ~n41942;
  assign n40302 = ~n40301 | ~n40300;
  assign n40304 = ~n40303 & ~n40302;
  assign P2_U2845 = ~n40305 | ~n40304;
  assign n40310 = ~n23636 & ~n40350;
  assign n40308 = ~n40306 | ~n41942;
  assign n40307 = ~P2_PHYADDRPOINTER_REG_2__SCAN_IN | ~n41921;
  assign n40309 = ~n40308 | ~n40307;
  assign n40318 = ~n40310 & ~n40309;
  assign n40316 = ~n40311 & ~n41931;
  assign n40314 = ~n40312 | ~n41934;
  assign n40313 = ~n41935 | ~P2_EBX_REG_2__SCAN_IN;
  assign n40315 = ~n40314 | ~n40313;
  assign n40317 = ~n40316 & ~n40315;
  assign n40321 = ~n40319 | ~n41718;
  assign n40322 = n40321 ^ n40320;
  assign n40323 = ~n40322 & ~n41919;
  assign n40326 = ~n40325 | ~n40579;
  assign P2_U2853 = ~n40327 | ~n40326;
  assign n40328 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN & ~n40442;
  assign n40333 = ~n40329 & ~n40328;
  assign n40332 = ~n40331 & ~n40330;
  assign n40334 = ~n40333 | ~n40332;
  assign n40337 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN | ~n40334;
  assign n40336 = ~n40980 | ~n40335;
  assign n40340 = ~n40339 & ~n40338;
  assign n40342 = ~n40341 & ~n40340;
  assign n40343 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN & ~n40342;
  assign n40346 = n40529 & P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign P3_U2846 = ~n40349 | ~n40348;
  assign n40353 = ~n40350 & ~n26530;
  assign n40351 = ~P2_PHYADDRPOINTER_REG_5__SCAN_IN | ~n41921;
  assign n40352 = ~n40351 | ~n40668;
  assign n40361 = ~n40353 & ~n40352;
  assign n40359 = ~n40354 & ~n41931;
  assign n40357 = ~n40355 | ~n41934;
  assign n40356 = ~n41935 | ~P2_EBX_REG_5__SCAN_IN;
  assign n40358 = ~n40357 | ~n40356;
  assign n40360 = ~n40359 & ~n40358;
  assign n40364 = ~n41204 & ~n40362;
  assign n40365 = n40364 ^ n40363;
  assign n40366 = ~n40365 & ~n41919;
  assign n40370 = ~n40367 & ~n40366;
  assign n40369 = ~n40368 | ~n41942;
  assign P2_U2850 = ~n40370 | ~n40369;
  assign n40380 = ~n40377 & ~n40960;
  assign n40379 = ~n42318 & ~n40378;
  assign n40381 = ~n40380 & ~n40379;
  assign n40399 = ~n41537 & ~P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n40386 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN & ~n42322;
  assign n40383 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN | ~n40382;
  assign n40385 = ~n40384 & ~n40383;
  assign n40499 = ~n40385 & ~n41537;
  assign n40397 = ~n40386 & ~n40499;
  assign n40396 = ~n40387 & ~n41240;
  assign n40392 = ~n40388 & ~n41235;
  assign n40390 = ~n40959 & ~n40389;
  assign n40391 = ~n40390 & ~n41540;
  assign n40394 = ~n40392 & ~n40391;
  assign P3_U2850 = ~n40407 | ~n40406;
  assign n40413 = ~n41546 | ~n40410;
  assign n40416 = ~n40968 | ~n40417;
  assign n40419 = ~n40418 & ~n40417;
  assign n40420 = ~n40419 & ~n41537;
  assign n40424 = ~n40420 & ~n40431;
  assign n40423 = ~n40422 | ~n40421;
  assign n40473 = ~n40424 | ~n40423;
  assign n40426 = ~n40425 & ~n40473;
  assign n40432 = ~n42338 & ~n40431;
  assign P3_U2843 = ~n40435 | ~n40434;
  assign n40438 = ~n40436 | ~n43305;
  assign n40437 = ~n43732 | ~P1_EAX_REG_14__SCAN_IN;
  assign n40440 = n40438 & n40437;
  assign n40439 = ~n32242 | ~n41130;
  assign P1_U2890 = ~n40440 | ~n40439;
  assign n40450 = ~n41235 & ~n40441;
  assign n40498 = ~n40443 & ~n40442;
  assign n40448 = ~n40444 & ~n40498;
  assign n40447 = ~n40446 | ~n40445;
  assign n40449 = ~n40448 | ~n40447;
  assign n40453 = ~n40450 & ~n40449;
  assign n40452 = ~n40451 | ~n41546;
  assign n40454 = ~n40453 | ~n40452;
  assign n40457 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN | ~n40454;
  assign n40456 = ~n40980 | ~n40455;
  assign n40458 = ~n40960 & ~P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n40461 = ~n42338 & ~n27696;
  assign P3_U2853 = ~n40464 | ~n40463;
  assign n40472 = n40471 & n40470;
  assign n40477 = ~n40472 & ~n41540;
  assign n40474 = ~n41535 | ~n40473;
  assign P3_U2842 = ~n40485 | ~n40484;
  assign n40489 = ~n40487;
  assign n40488 = ~n43709 | ~P1_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n40492 = n40489 & n40488;
  assign n40491 = ~n43362 | ~n40490;
  assign n40495 = ~n40492 | ~n40491;
  assign P1_U2986 = ~n40497 | ~n40496;
  assign n40518 = ~n42338 & ~n27697;
  assign n40502 = ~n40499 & ~n40498;
  assign n40501 = ~n41542 | ~n40500;
  assign n40507 = ~n40502 | ~n40501;
  assign n40504 = ~n41546 | ~n40503;
  assign n40506 = ~n40505 | ~n40504;
  assign n40990 = ~n40507 & ~n40506;
  assign n40988 = ~n27696 | ~n40508;
  assign n40509 = ~n40990 | ~n40988;
  assign n40512 = ~n40509 | ~P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n40511 = ~n40980 | ~n40510;
  assign n40514 = ~n40960 & ~n40513;
  assign P3_U2852 = ~n40520 | ~n40519;
  assign n40522 = ~n42320 | ~n40521;
  assign n40525 = ~n40523 | ~n40522;
  assign P3_U2841 = ~n40541 | ~n40540;
  assign n40548 = ~n42135 | ~n40542;
  assign n40543 = ~P3_EBX_REG_24__SCAN_IN | ~n43930;
  assign n41058 = ~n40545 & ~n40544;
  assign P3_U2679 = ~n40548 | ~n40547;
  assign n40552 = ~n43306 | ~n40550;
  assign n40551 = ~n43737 | ~BUF1_REG_17__SCAN_IN;
  assign n40556 = ~n40552 | ~n40551;
  assign n40554 = ~n43738 | ~DATAI_17_;
  assign n40553 = ~n43732 | ~P1_EAX_REG_17__SCAN_IN;
  assign n40555 = ~n40554 | ~n40553;
  assign n40557 = ~n40556 & ~n40555;
  assign P1_U2887 = ~n40558 | ~n40557;
  assign n40563 = ~n40559 & ~n41931;
  assign n40561 = ~n41920 | ~P2_REIP_REG_4__SCAN_IN;
  assign n40560 = ~n41921 | ~P2_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n40562 = ~n40561 | ~n40560;
  assign n40564 = ~n40563 & ~n40562;
  assign n40569 = ~n40564 | ~n40668;
  assign n40567 = ~n40565 | ~n41942;
  assign n40566 = ~P2_EBX_REG_4__SCAN_IN | ~n41935;
  assign n40568 = ~n40567 | ~n40566;
  assign n40571 = ~n40570 | ~n41934;
  assign n40575 = ~n40573 | ~n41718;
  assign n40576 = n40575 ^ n40574;
  assign n40577 = ~n40576 & ~n41919;
  assign n40581 = ~n40580 | ~n40579;
  assign P2_U2851 = ~n40582 | ~n40581;
  assign n40599 = n42219 & n40602;
  assign n40595 = ~n42429 & ~n41926;
  assign n40583 = ~P2_REIP_REG_15__SCAN_IN | ~n41920;
  assign n40591 = ~n40668 | ~n40583;
  assign n40584 = ~n42429 & ~n40670;
  assign n40585 = ~n40584 & ~n40669;
  assign n40589 = ~n40585 | ~n40625;
  assign n40588 = ~n42209 | ~n41934;
  assign n40590 = ~n40589 | ~n40588;
  assign n40593 = ~n40591 & ~n40590;
  assign n40592 = ~P2_PHYADDRPOINTER_REG_15__SCAN_IN | ~n41921;
  assign n40594 = ~n40593 | ~n40592;
  assign n40597 = ~n40595 & ~n40594;
  assign n40596 = ~P2_EBX_REG_15__SCAN_IN | ~n41935;
  assign n40600 = ~n42424 | ~n41942;
  assign P2_U2840 = ~n40601 | ~n40600;
  assign n40619 = n42117 & n40602;
  assign n40615 = ~n42145 & ~n41926;
  assign n40603 = ~P2_REIP_REG_13__SCAN_IN | ~n41920;
  assign n40611 = ~n40668 | ~n40603;
  assign n40604 = ~n42145 & ~n40646;
  assign n40605 = ~n40604 & ~n40669;
  assign n40609 = ~n40605 | ~n40671;
  assign n40608 = ~n42099 | ~n41934;
  assign n40610 = ~n40609 | ~n40608;
  assign n40613 = ~n40611 & ~n40610;
  assign n40612 = ~P2_PHYADDRPOINTER_REG_13__SCAN_IN | ~n41921;
  assign n40614 = ~n40613 | ~n40612;
  assign n40617 = ~n40615 & ~n40614;
  assign n40616 = ~P2_EBX_REG_13__SCAN_IN | ~n41935;
  assign n40621 = ~n40620 | ~n41942;
  assign P2_U2842 = ~n40622 | ~n40621;
  assign n40642 = ~n42633 & ~n41931;
  assign n40638 = ~n42393 & ~n41926;
  assign n40623 = ~P2_REIP_REG_16__SCAN_IN | ~n41920;
  assign n40634 = ~n40668 | ~n40623;
  assign n40628 = ~n40624 & ~n40669;
  assign n40627 = ~n40626 | ~n40625;
  assign n40632 = ~n40628 | ~n40627;
  assign n40631 = ~n42243 | ~n41934;
  assign n40633 = ~n40632 | ~n40631;
  assign n40636 = ~n40634 & ~n40633;
  assign n40635 = ~P2_PHYADDRPOINTER_REG_16__SCAN_IN | ~n41921;
  assign n40637 = ~n40636 | ~n40635;
  assign n40640 = ~n40638 & ~n40637;
  assign n40639 = ~P2_EBX_REG_16__SCAN_IN | ~n41935;
  assign n40643 = ~n42637 | ~n41942;
  assign P2_U2839 = ~n40644 | ~n40643;
  assign n40664 = ~n42309 & ~n41931;
  assign n40660 = ~n42457 & ~n41926;
  assign n40645 = ~P2_REIP_REG_12__SCAN_IN | ~n41920;
  assign n40656 = ~n40668 | ~n40645;
  assign n40650 = ~n40646 & ~n40669;
  assign n40649 = ~n40648 | ~n40647;
  assign n40654 = ~n40650 | ~n40649;
  assign n40653 = ~n42094 | ~n41934;
  assign n40655 = ~n40654 | ~n40653;
  assign n40658 = ~n40656 & ~n40655;
  assign n40657 = ~P2_PHYADDRPOINTER_REG_12__SCAN_IN | ~n41921;
  assign n40659 = ~n40658 | ~n40657;
  assign n40662 = ~n40660 & ~n40659;
  assign n40661 = ~P2_EBX_REG_12__SCAN_IN | ~n41935;
  assign n40665 = ~n42452 | ~n41942;
  assign P2_U2843 = ~n40666 | ~n40665;
  assign n40688 = n42665 & n40602;
  assign n40684 = ~n42847 & ~n41926;
  assign n40667 = ~P2_REIP_REG_14__SCAN_IN | ~n41920;
  assign n40680 = ~n40668 | ~n40667;
  assign n40674 = ~n40670 & ~n40669;
  assign n40673 = ~n40672 | ~n40671;
  assign n40678 = ~n40674 | ~n40673;
  assign n40677 = ~n42204 | ~n41934;
  assign n40679 = ~n40678 | ~n40677;
  assign n40682 = ~n40680 & ~n40679;
  assign n40681 = ~P2_PHYADDRPOINTER_REG_14__SCAN_IN | ~n41921;
  assign n40683 = ~n40682 | ~n40681;
  assign n40686 = ~n40684 & ~n40683;
  assign n40685 = ~P2_EBX_REG_14__SCAN_IN | ~n41935;
  assign n40689 = ~n42842;
  assign n40690 = ~n40689 | ~n41942;
  assign P2_U2841 = ~n40691 | ~n40690;
  assign n40701 = n40692 | n43358;
  assign n40699 = ~n40707 & ~n43729;
  assign n40694 = ~n40693 & ~n40709;
  assign n40697 = ~n40695 & ~n40694;
  assign n40696 = ~n43362 | ~n40708;
  assign n40698 = ~n40697 | ~n40696;
  assign P1_U2984 = ~n40701 | ~n40700;
  assign n40702 = ~n42400 & ~n40703;
  assign n40722 = ~P1_REIP_REG_15__SCAN_IN | ~n41124;
  assign n40705 = ~n42185 & ~n40703;
  assign n40720 = n40705 & n40704;
  assign n40714 = ~n40708 | ~n43559;
  assign n40712 = ~n43796 | ~P1_EBX_REG_15__SCAN_IN;
  assign n40710 = ~n40709 & ~n41129;
  assign n40711 = ~n43469 & ~n40710;
  assign n40713 = n40712 & n40711;
  assign P1_U2825 = ~n40722 | ~n40721;
  assign n40730 = ~n41560;
  assign n40728 = ~n40724;
  assign n40870 = ~n40726 | ~n40725;
  assign n40727 = ~n41520 | ~n40870;
  assign n40729 = ~n40728 | ~n40727;
  assign n40742 = ~n40730 | ~n40729;
  assign n40737 = ~n40732 & ~n40731;
  assign n40735 = ~n41100 | ~n40733;
  assign n40736 = ~n40735 | ~n40734;
  assign n40871 = ~n40737 & ~n40736;
  assign n40739 = n41095 & n40738;
  assign n40740 = ~n40739 & ~P3_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n40741 = ~n40871 & ~n40740;
  assign n40756 = ~n40742 & ~n40741;
  assign n40749 = n41233 & n40847;
  assign P3_U2804 = ~n40756 | ~n40755;
  assign n40764 = ~n42242 | ~n40760;
  assign n40761 = ~n41078;
  assign n40763 = n40762 & n41078;
  assign n40942 = n40766 | n40765;
  assign n40944 = ~n43880 | ~P2_REIP_REG_7__SCAN_IN;
  assign n40774 = ~n40944;
  assign n40768 = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN | ~n40767;
  assign n41069 = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN & ~n40768;
  assign n40772 = ~n41069;
  assign n41068 = ~n40770 | ~n40769;
  assign n40771 = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN | ~n41068;
  assign n40773 = ~n40772 | ~n40771;
  assign n40777 = ~n40774 & ~n40773;
  assign n40776 = ~n43583 | ~n40775;
  assign n40779 = ~n40777 | ~n40776;
  assign n40778 = ~n43886 & ~n40943;
  assign n40780 = n40779 | n40778;
  assign P2_U3039 = ~n40783 | ~n40782;
  assign n40792 = ~n40784 & ~n43358;
  assign n40785 = ~n43709 | ~P1_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n40788 = ~n40786 | ~n40785;
  assign n40787 = ~n43713 & ~n41131;
  assign n40790 = ~n40788 & ~n40787;
  assign n40789 = ~n41130 | ~n43367;
  assign P1_U2985 = n40792 | n40791;
  assign n40794 = ~n40793 & ~n40798;
  assign n40801 = ~n40795 | ~n40794;
  assign n40799 = ~n40797 | ~n40796;
  assign n40800 = ~n40799 | ~n40798;
  assign n40808 = ~n40801 | ~n40800;
  assign P1_U3015 = ~n40808 | ~n40807;
  assign n40814 = ~n42135 | ~n40809;
  assign n40811 = ~P3_EBX_REG_25__SCAN_IN | ~n43930;
  assign n41390 = ~n41058 | ~P3_EBX_REG_25__SCAN_IN;
  assign P3_U2678 = ~n40814 | ~n40813;
  assign n40822 = ~n40821 & ~n40820;
  assign n40826 = ~n40822 | ~n42320;
  assign n40825 = ~n40824 | ~n40823;
  assign n40827 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~n40997;
  assign n40837 = ~n42321 | ~n40827;
  assign n40828 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~n41537;
  assign n40829 = ~n41005 | ~n40828;
  assign n40834 = ~n41538 & ~n40829;
  assign n40831 = ~n40968 | ~n40830;
  assign n40833 = ~n40832 | ~n40831;
  assign n40835 = ~n40834 & ~n40833;
  assign P3_U2837 = ~n40846 | ~n40845;
  assign n40849 = ~n40848 & ~n41259;
  assign n40867 = ~n40864 | ~n41400;
  assign n41260 = ~n40865 & ~n35543;
  assign n40866 = ~n41260;
  assign n40868 = ~n40867 | ~n40866;
  assign n40878 = n40869 | n40868;
  assign n41157 = ~n40871 | ~n40870;
  assign n40874 = ~P3_PHYADDRPOINTER_REG_28__SCAN_IN | ~n41157;
  assign n41159 = ~n41093 & ~n40872;
  assign n40873 = ~n41159 | ~n41092;
  assign n40876 = n40874 & n40873;
  assign n40875 = ~P3_PHYADDRPOINTER_REG_28__SCAN_IN & ~P3_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n40877 = ~n40876 & ~n40875;
  assign P3_U2802 = ~n40880 | ~n40879;
  assign n40890 = ~n40881 & ~n41307;
  assign n40885 = ~n40882 & ~n41316;
  assign n40884 = ~n41319 & ~n40883;
  assign n40888 = ~n40885 & ~n40884;
  assign n40887 = ~n40886 | ~n41310;
  assign P2_U3173 = ~n40893 | ~n40892;
  assign n40903 = ~n40894 & ~n41319;
  assign n40898 = ~n41307 & ~n40895;
  assign n40897 = ~n40896 & ~n41316;
  assign n40901 = ~n40898 & ~n40897;
  assign n40900 = ~n40899 | ~n41310;
  assign n40905 = ~n40903 & ~n40902;
  assign P2_U3171 = ~n40905 | ~n40904;
  assign n40915 = ~n40906 & ~n41319;
  assign n40910 = ~n41307 & ~n40907;
  assign n40909 = ~n40908 & ~n41316;
  assign n40913 = ~n40910 & ~n40909;
  assign n40912 = ~n40911 | ~n41310;
  assign n40917 = ~n40915 & ~n40914;
  assign P2_U3170 = ~n40917 | ~n40916;
  assign n40919 = ~n40918 | ~n41718;
  assign n40920 = ~n40919 ^ n43326;
  assign n40940 = ~n40920 | ~n41206;
  assign n40922 = ~n40921;
  assign n40924 = ~n40923 | ~n40922;
  assign n43196 = ~n41209 | ~n40924;
  assign n40930 = n41935 & P2_EBX_REG_26__SCAN_IN;
  assign n40928 = ~n41920 | ~P2_REIP_REG_26__SCAN_IN;
  assign n40927 = ~n41921 | ~P2_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n40929 = ~n40928 | ~n40927;
  assign n40931 = ~n40930 & ~n40929;
  assign n40938 = n40934 | n40933;
  assign P2_U2829 = ~n40940 | ~n40939;
  assign n40947 = ~n43915 & ~n40943;
  assign n40945 = ~n43917 | ~P2_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n40946 = ~n40945 | ~n40944;
  assign n40951 = ~n40947 & ~n40946;
  assign n40949 = ~n40948;
  assign n40950 = ~n43896 | ~n40949;
  assign n40952 = ~n40951 | ~n40950;
  assign P2_U3007 = ~n40955 | ~n40954;
  assign n40957 = ~n42338 & ~n40962;
  assign n40978 = ~n40957 & ~n40956;
  assign n40975 = ~n40958 | ~n40980;
  assign n40966 = ~n40965 | ~n40964;
  assign n40971 = ~n40967 & ~n40966;
  assign n40970 = ~n40969 | ~n40968;
  assign P3_U2849 = ~n40978 | ~n40977;
  assign n40984 = ~n40980 | ~n40979;
  assign n40996 = n40987 & n40986;
  assign n40989 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN | ~n40988;
  assign n40991 = ~n40989 | ~n41005;
  assign n40995 = ~n40994 | ~P3_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign P3_U2851 = ~n40996 | ~n40995;
  assign n41001 = ~n40997;
  assign n41000 = ~n40998;
  assign n41007 = ~n41005 | ~n41004;
  assign P3_U2838 = ~n41018 | ~n41017;
  assign n41038 = ~n41019 | ~P1_REIP_REG_16__SCAN_IN;
  assign n41021 = ~n42185 & ~P1_REIP_REG_16__SCAN_IN;
  assign n41036 = n41021 & n41020;
  assign n41032 = ~n41129 & ~n41023;
  assign n41028 = ~n43796 | ~P1_EBX_REG_16__SCAN_IN;
  assign n41026 = ~n42175 & ~n41025;
  assign n41027 = ~n41026 & ~n43469;
  assign n41029 = n41028 & n41027;
  assign P1_U2824 = ~n41038 | ~n41037;
  assign n41042 = ~n43306 | ~n41040;
  assign n41041 = ~n43737 | ~BUF1_REG_19__SCAN_IN;
  assign n41046 = ~n41042 | ~n41041;
  assign n41044 = ~n43738 | ~DATAI_19_;
  assign n41043 = ~n43732 | ~P1_EAX_REG_19__SCAN_IN;
  assign n41045 = ~n41044 | ~n41043;
  assign n41047 = ~n41046 & ~n41045;
  assign P1_U2885 = ~n41048 | ~n41047;
  assign n41057 = ~n41454 | ~n32242;
  assign n41051 = ~n43306 | ~n41049;
  assign n41050 = ~n43737 | ~BUF1_REG_18__SCAN_IN;
  assign n41055 = ~n41051 | ~n41050;
  assign n41053 = ~n43738 | ~DATAI_18_;
  assign n41052 = ~n43732 | ~P1_EAX_REG_18__SCAN_IN;
  assign n41054 = ~n41053 | ~n41052;
  assign n41056 = ~n41055 & ~n41054;
  assign P1_U2886 = ~n41057 | ~n41056;
  assign n41061 = ~n42135 & ~n41058;
  assign n41060 = ~n41059 & ~P3_EBX_REG_25__SCAN_IN;
  assign n41062 = ~n41061 & ~n41060;
  assign n41066 = ~n42135 | ~n41065;
  assign P3_U2677 = ~n41067 | ~n41066;
  assign n41071 = ~n41068;
  assign n41070 = ~n41069 & ~n41072;
  assign n41075 = ~n41071 | ~n41070;
  assign n41074 = ~n41073 | ~n41072;
  assign n41090 = ~n41075 | ~n41074;
  assign n41080 = ~n41491 ^ P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n41086 = ~n41171 | ~n43876;
  assign n41082 = ~n43583 | ~n41081;
  assign n41178 = ~n43880 | ~P2_REIP_REG_8__SCAN_IN;
  assign n41084 = ~n41082 | ~n41178;
  assign n41083 = ~n43886 & ~n41172;
  assign n41085 = ~n41084 & ~n41083;
  assign P2_U3038 = ~n41090 | ~n41089;
  assign n41094 = ~n41093 & ~n41092;
  assign n41097 = ~n41095 | ~n41094;
  assign n41103 = ~n41097 | ~n41096;
  assign n41404 = ~n41097 & ~n41096;
  assign n41102 = n41098 | n41404;
  assign n41101 = ~n41100 | ~n41099;
  assign n41417 = ~n41102 | ~n41101;
  assign n41110 = ~n41103 | ~n41417;
  assign n41108 = ~n41104;
  assign n41418 = ~P3_PHYADDRPOINTER_REG_29__SCAN_IN & ~n41403;
  assign n41106 = ~n41418 & ~n41400;
  assign n41107 = ~n41106 & ~n41105;
  assign n41109 = ~n41108 & ~n41107;
  assign n41116 = ~n41408 & ~n41113;
  assign P3_U2801 = ~n41123 | ~n41122;
  assign n41144 = ~n41124 | ~P1_REIP_REG_14__SCAN_IN;
  assign n41126 = ~n42185 & ~P1_REIP_REG_14__SCAN_IN;
  assign n41142 = n41126 & n41125;
  assign n41138 = ~n41129 & ~n41128;
  assign n41134 = ~n43796 | ~P1_EBX_REG_14__SCAN_IN;
  assign n41132 = ~n42175 & ~n41131;
  assign n41133 = ~n41132 & ~n43469;
  assign n41135 = n41134 & n41133;
  assign P1_U2826 = ~n41144 | ~n41143;
  assign n42341 = ~n41145 | ~P3_REIP_REG_27__SCAN_IN;
  assign n41163 = ~n41520 & ~n41156;
  assign n41161 = ~P3_PHYADDRPOINTER_REG_27__SCAN_IN | ~n41157;
  assign n41160 = ~n41159 | ~n41158;
  assign n41162 = ~n41161 | ~n41160;
  assign n41164 = ~n41163 & ~n41162;
  assign P3_U2803 = ~n41169 | ~n41168;
  assign n41184 = ~n41170 & ~n43924;
  assign n41175 = ~n43813 | ~n41173;
  assign n41174 = ~n43917 | ~P2_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n41180 = ~n41175 | ~n41174;
  assign n41177 = ~n43896 | ~n41176;
  assign n41179 = ~n41178 | ~n41177;
  assign n41181 = ~n41180 & ~n41179;
  assign P2_U3006 = n41184 | n41183;
  assign n41188 = ~n41185;
  assign n41193 = ~n41186 | ~n41188;
  assign n41189 = ~n41187;
  assign n41190 = ~n41189 | ~n41188;
  assign n41192 = ~n41191 | ~n41190;
  assign n41202 = n41275 | n43358;
  assign n41277 = ~n43469 | ~P1_REIP_REG_17__SCAN_IN;
  assign n41195 = ~n43709 | ~P1_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n41198 = n41277 & n41195;
  assign n41197 = ~n43362 | ~n41196;
  assign n41199 = ~n41198 | ~n41197;
  assign P1_U2982 = ~n41202 | ~n41201;
  assign n41205 = ~n41204 & ~n41203;
  assign n41207 = ~n41205 ^ n43654;
  assign n41228 = ~n41207 | ~n41206;
  assign n41210 = ~n41209 | ~n41208;
  assign n41220 = ~n43607 | ~n41934;
  assign n41218 = ~n41214 & ~n41213;
  assign n41216 = ~n41920 | ~P2_REIP_REG_27__SCAN_IN;
  assign n41215 = ~n41921 | ~P2_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n41217 = ~n41216 | ~n41215;
  assign n41219 = ~n41218 & ~n41217;
  assign n41226 = n41222 | n41221;
  assign P2_U2828 = ~n41228 | ~n41227;
  assign n41247 = n41236 | n41235;
  assign n41241 = ~n41240 & ~n41239;
  assign n41251 = ~n41250;
  assign n41261 = ~n42338 & ~n41259;
  assign n41262 = ~n41261 & ~n41260;
  assign P3_U2834 = ~n41263 | ~n41262;
  assign n41267 = ~n41265 & ~n35967;
  assign n41266 = ~n43525 & ~P2_EBX_REG_23__SCAN_IN;
  assign P2_U2864 = n41269 | n41268;
  assign n41274 = ~n42364 | ~n41272;
  assign n41270 = ~n43330 | ~n41979;
  assign n41273 = n41965 | n41272;
  assign n41282 = ~n41274 | ~n41273;
  assign P1_U3014 = ~n41282 | ~n41281;
  assign n41288 = ~n41283 & ~n41307;
  assign n41285 = ~n41284 | ~n41310;
  assign n41292 = ~n41289 & ~n41316;
  assign n41291 = ~n41319 & ~n41290;
  assign n41293 = ~n41292 & ~n41291;
  assign P2_U3175 = ~n41294 | ~n41293;
  assign n41300 = ~n41295 & ~n41307;
  assign n41297 = ~n41296 | ~n41310;
  assign n41304 = ~n41301 & ~n41316;
  assign n41303 = ~n41319 & ~n41302;
  assign n41305 = ~n41304 & ~n41303;
  assign P2_U3174 = ~n41306 | ~n41305;
  assign n41315 = ~n41308 & ~n41307;
  assign n41313 = ~P2_INSTQUEUE_REG_15__4__SCAN_IN | ~n41309;
  assign n41312 = ~n41311 | ~n41310;
  assign n41323 = ~n41315 & ~n41314;
  assign n41321 = ~n41317 & ~n41316;
  assign n41320 = ~n41319 & ~n41318;
  assign n41322 = ~n41321 & ~n41320;
  assign P2_U3172 = ~n41323 | ~n41322;
  assign n41379 = ~n41325 | ~n41324;
  assign n41328 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~n41331;
  assign n41353 = n41333 | n41332;
  assign n41334 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n41343 = ~n41345 | ~n41341;
  assign n41346 = ~n41345 & ~n41344;
  assign n41347 = ~n41346 & ~n41371;
  assign n41360 = ~P3_MORE_REG_SCAN_IN & ~P3_FLUSH_REG_SCAN_IN;
  assign n41361 = ~n41360 & ~n41359;
  assign n41364 = ~n41362 & ~n41361;
  assign n41366 = ~n41364 | ~n41363;
  assign n41367 = ~n41366 & ~n41365;
  assign n41377 = n41374 | n42024;
  assign n41376 = ~n41375 | ~n32190;
  assign n41383 = ~n41382 | ~n42016;
  assign n41385 = ~n41384 & ~n41383;
  assign P3_U2997 = ~n41387 | ~n41386;
  assign n41396 = ~n42135 | ~n41388;
  assign n41392 = ~P3_EBX_REG_27__SCAN_IN | ~n43930;
  assign P3_U2676 = ~n41396 | ~n41395;
  assign n41405 = ~n41403 & ~n41402;
  assign n41419 = ~n41405 & ~n41404;
  assign n41406 = ~n41419 & ~P3_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n41412 = ~n41406 | ~P3_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n41409 = n41408 | n41407;
  assign n41517 = ~n41418 & ~n41417;
  assign n41523 = P3_PHYADDRPOINTER_REG_30__SCAN_IN | n41419;
  assign n41420 = ~n41517 | ~n41523;
  assign P3_U2799 = n41424 | n41423;
  assign n41428 = ~n43306 | ~n41426;
  assign n41427 = ~n43737 | ~BUF1_REG_21__SCAN_IN;
  assign n41432 = ~n41428 | ~n41427;
  assign n41430 = ~n43738 | ~DATAI_21_;
  assign n41429 = ~n43732 | ~P1_EAX_REG_21__SCAN_IN;
  assign n41431 = ~n41430 | ~n41429;
  assign n41433 = ~n41432 & ~n41431;
  assign P1_U2883 = ~n41434 | ~n41433;
  assign n41440 = ~n44023 | ~P1_EBX_REG_20__SCAN_IN;
  assign P1_U2852 = ~n41443 | ~n41442;
  assign n41446 = ~n43796 | ~P1_EBX_REG_18__SCAN_IN;
  assign n41445 = ~n43559 | ~n41444;
  assign n41449 = ~n41446 | ~n41445;
  assign n41447 = ~P1_PHYADDRPOINTER_REG_18__SCAN_IN | ~n43797;
  assign n41448 = ~n43033 | ~n41447;
  assign n41460 = ~n41449 & ~n41448;
  assign n41452 = ~P1_REIP_REG_18__SCAN_IN & ~n41450;
  assign P1_U2822 = ~n41460 | ~n41459;
  assign n41464 = ~n43306 | ~n41462;
  assign n41463 = ~n43737 | ~BUF1_REG_20__SCAN_IN;
  assign n41468 = ~n41464 | ~n41463;
  assign n41466 = ~n43738 | ~DATAI_20_;
  assign n41465 = ~n43732 | ~P1_EAX_REG_20__SCAN_IN;
  assign n41467 = ~n41466 | ~n41465;
  assign n41469 = ~n41468 & ~n41467;
  assign P1_U2884 = ~n41470 | ~n41469;
  assign n41930 = ~n41471;
  assign n41480 = ~n41930 & ~n41472;
  assign n41478 = n41473 & P2_REIP_REG_31__SCAN_IN;
  assign n41476 = ~n41474 | ~P2_EAX_REG_31__SCAN_IN;
  assign n41475 = ~n28191 | ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n41477 = ~n41476 | ~n41475;
  assign n41479 = ~n41478 & ~n41477;
  assign n43847 = n41480 ^ n41479;
  assign n41487 = n43847 | n43695;
  assign n41485 = ~n42802 & ~n41481;
  assign n41483 = ~n43690 | ~BUF1_REG_31__SCAN_IN;
  assign n41482 = ~n43698 | ~P2_EAX_REG_31__SCAN_IN;
  assign n41484 = ~n41483 | ~n41482;
  assign n41486 = ~n41485 & ~n41484;
  assign P2_U2888 = ~n41487 | ~n41486;
  assign n41489 = ~n41699 & ~n43924;
  assign n41700 = n41488 | P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n41494 = n41490 | P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n41497 = n41495 & P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n41498 = ~n41497 & ~n41496;
  assign n41500 = ~n41707;
  assign n41503 = ~n43915 & ~n41500;
  assign n41501 = ~n43917 | ~P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n41704 = ~n43880 | ~P2_REIP_REG_9__SCAN_IN;
  assign n41502 = ~n41501 | ~n41704;
  assign n41507 = ~n41503 & ~n41502;
  assign n41505 = ~n41504;
  assign n41506 = ~n43896 | ~n41505;
  assign n41508 = ~n41507 | ~n41506;
  assign P2_U3005 = ~n41511 | ~n41510;
  assign n41522 = ~n41518 & ~n41517;
  assign n41521 = ~n41520 & ~n41519;
  assign n41524 = ~n41522 & ~n41521;
  assign n41525 = ~n41524 | ~n41523;
  assign n41533 = n41532 | n41531;
  assign P3_U2800 = ~n41534 | ~n41533;
  assign n41551 = ~n41536 | ~n41535;
  assign n41550 = ~n41538 & ~n41537;
  assign n41544 = ~n41540 & ~n41539;
  assign P3_U2836 = ~n41563 | ~n41562;
  assign n41570 = ~n41569;
  assign n41617 = ~n41789 & ~n41570;
  assign n41572 = ~n43499 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n41571 = ~n43496 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n41576 = ~n41572 | ~n41571;
  assign n41574 = ~n43500 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n41573 = ~n43503 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n41575 = ~n41574 | ~n41573;
  assign n41582 = ~n41576 & ~n41575;
  assign n41577 = ~n43495 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n41580 = ~n41577 | ~n43509;
  assign n41579 = ~n22927 & ~n41578;
  assign n41581 = ~n41580 & ~n41579;
  assign n41586 = ~n41582 | ~n41581;
  assign n41584 = ~n22911 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n41583 = ~n43484 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n41585 = ~n41584 | ~n41583;
  assign n41610 = ~n41586 & ~n41585;
  assign n41587 = ~n43495 | ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n41590 = ~n41587 | ~n43490;
  assign n41589 = ~n43514 & ~n41588;
  assign n41596 = ~n41590 & ~n41589;
  assign n41594 = ~n43098 & ~n41591;
  assign n41593 = ~n43100 & ~n41592;
  assign n41595 = ~n41594 & ~n41593;
  assign n41608 = ~n41596 | ~n41595;
  assign n41600 = ~n43092 & ~n41597;
  assign n41599 = ~n22927 & ~n41598;
  assign n41606 = ~n41600 & ~n41599;
  assign n41604 = ~n43094 & ~n41601;
  assign n41603 = ~n43408 & ~n41602;
  assign n41605 = ~n41604 & ~n41603;
  assign n41607 = ~n41606 | ~n41605;
  assign n41609 = ~n41608 & ~n41607;
  assign n41787 = ~n41610 & ~n41609;
  assign n41612 = ~n43525 & ~P2_EBX_REG_24__SCAN_IN;
  assign P2_U2863 = n41615 | n41614;
  assign n41616 = ~n41783;
  assign n41618 = ~n41617 | ~n41787;
  assign n41621 = ~n43495 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n41620 = ~n43499 | ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n41630 = ~n41621 | ~n41620;
  assign n41623 = ~n43496 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n41622 = ~n43503 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n41627 = ~n41623 | ~n41622;
  assign n41625 = ~n22911 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n41624 = ~n43483 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n41626 = ~n41625 | ~n41624;
  assign n41628 = ~n41627 & ~n41626;
  assign n41629 = ~n43509 | ~n41628;
  assign n41636 = ~n41630 & ~n41629;
  assign n41634 = ~n43408 & ~n41631;
  assign n41632 = ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n41633 = ~n43514 & ~n41632;
  assign n41635 = ~n41634 & ~n41633;
  assign n41655 = ~n41636 | ~n41635;
  assign n41638 = ~n43495 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n41637 = ~n43499 | ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n41647 = ~n41638 | ~n41637;
  assign n41640 = ~n22911 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n41639 = ~n43484 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n41644 = ~n41640 | ~n41639;
  assign n41642 = ~n43496 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n41641 = ~n43483 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n41643 = ~n41642 | ~n41641;
  assign n41645 = ~n41644 & ~n41643;
  assign n41646 = ~n43490 | ~n41645;
  assign n41653 = ~n41647 & ~n41646;
  assign n41651 = ~n43408 & ~n41648;
  assign n41649 = ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n41650 = ~n43100 & ~n41649;
  assign n41652 = ~n41651 & ~n41650;
  assign n41654 = ~n41653 | ~n41652;
  assign n41782 = ~n41655 | ~n41654;
  assign n41786 = ~n41782;
  assign n41658 = ~BUF2_REG_25__SCAN_IN;
  assign n41663 = ~n42802 & ~n41658;
  assign n41661 = ~n42804 | ~n41659;
  assign n41660 = ~n43698 | ~P2_EAX_REG_25__SCAN_IN;
  assign n41662 = ~n41661 | ~n41660;
  assign n41665 = ~n41663 & ~n41662;
  assign n41664 = ~n43690 | ~BUF1_REG_25__SCAN_IN;
  assign n41666 = ~n41665 | ~n41664;
  assign P2_U2894 = ~n41669 | ~n41668;
  assign n41674 = n43992 | n42017;
  assign n41673 = ~n41672;
  assign P3_U3282 = ~n41674 | ~n41673;
  assign n41676 = n43525 | P2_EBX_REG_25__SCAN_IN;
  assign P2_U2862 = ~n41679 | ~n41678;
  assign n41686 = ~n42135 | ~n41680;
  assign P3_U2675 = ~n41686 | ~n41685;
  assign n41690 = ~n43306 | ~n41688;
  assign n41689 = ~n43737 | ~BUF1_REG_23__SCAN_IN;
  assign n41694 = ~n41690 | ~n41689;
  assign n41692 = ~n43738 | ~DATAI_23_;
  assign n41691 = ~n43732 | ~P1_EAX_REG_23__SCAN_IN;
  assign n41693 = ~n41692 | ~n41691;
  assign n41695 = ~n41694 & ~n41693;
  assign P1_U2881 = ~n41696 | ~n41695;
  assign n41717 = ~n42558 | ~n41697;
  assign n41715 = ~n41698 & ~n41697;
  assign n41701 = ~n41699 & ~n43893;
  assign n41706 = ~n43877 & ~n41703;
  assign n41705 = ~n41704;
  assign n41709 = ~n41706 & ~n41705;
  assign n41708 = ~n43767 | ~n41707;
  assign n41710 = ~n41709 | ~n41708;
  assign P2_U3037 = ~n41717 | ~n41716;
  assign n41720 = ~n41719 | ~n41718;
  assign n41721 = n41720 ^ n43774;
  assign n41739 = ~n41721 & ~n41919;
  assign n41723 = ~n41920 | ~P2_REIP_REG_28__SCAN_IN;
  assign n41722 = ~n41921 | ~P2_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n41729 = ~n43668 | ~n41934;
  assign n41738 = n41737 | n41736;
  assign P2_U2827 = n41739 | n41738;
  assign n41740 = ~P1_INSTADDRPOINTER_REG_18__SCAN_IN & ~P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n41741 = ~n41740 & ~n42364;
  assign n41751 = n41741 & n41962;
  assign P1_U3013 = n41751 | n41750;
  assign n41753 = ~BUF2_REG_24__SCAN_IN | ~n43689;
  assign n41752 = ~BUF1_REG_24__SCAN_IN | ~n43690;
  assign n41767 = ~n41753 | ~n41752;
  assign n41761 = ~n43697 & ~n41757;
  assign n41760 = ~n41759 & ~n41758;
  assign n41762 = ~n41761 & ~n41760;
  assign n41766 = n41765 | n41764;
  assign P2_U2895 = n41767 | n41766;
  assign n41768 = ~n44023 | ~P1_EBX_REG_22__SCAN_IN;
  assign P1_U2850 = ~n41771 | ~n41770;
  assign n41775 = ~n43306 | ~n41773;
  assign n41774 = ~n43737 | ~BUF1_REG_22__SCAN_IN;
  assign n41779 = ~n41775 | ~n41774;
  assign n41777 = ~n43738 | ~DATAI_22_;
  assign n41776 = ~n43732 | ~P1_EAX_REG_22__SCAN_IN;
  assign n41778 = ~n41777 | ~n41776;
  assign n41780 = ~n41779 & ~n41778;
  assign P1_U2882 = ~n41781 | ~n41780;
  assign n41788 = ~n41787 | ~n41786;
  assign n41792 = ~n41789 & ~n41788;
  assign n41791 = ~n41790;
  assign n42755 = n41792 & n41791;
  assign n41794 = ~n43500 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n41793 = ~n43499 | ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n41803 = ~n41794 | ~n41793;
  assign n41796 = ~n43495 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n41795 = ~n43483 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n41800 = ~n41796 | ~n41795;
  assign n41798 = ~n43496 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n41797 = ~n22911 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n41799 = ~n41798 | ~n41797;
  assign n41801 = ~n41800 & ~n41799;
  assign n41802 = ~n43509 | ~n41801;
  assign n41809 = ~n41803 & ~n41802;
  assign n41807 = ~n43514 & ~n41804;
  assign n41806 = ~n43100 & ~n41805;
  assign n41808 = ~n41807 & ~n41806;
  assign n41828 = ~n41809 | ~n41808;
  assign n41811 = ~n43503 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n41810 = ~n43499 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n41820 = ~n41811 | ~n41810;
  assign n41813 = ~n43483 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n41812 = ~n43484 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n41817 = ~n41813 | ~n41812;
  assign n41815 = ~n43496 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n41814 = ~n43495 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n41816 = ~n41815 | ~n41814;
  assign n41818 = ~n41817 & ~n41816;
  assign n41819 = ~n43490 | ~n41818;
  assign n41826 = ~n41820 & ~n41819;
  assign n41824 = ~n43098 & ~n41821;
  assign n41823 = ~n43408 & ~n41822;
  assign n41825 = ~n41824 & ~n41823;
  assign n41827 = ~n41826 | ~n41825;
  assign n42753 = ~n41828 | ~n41827;
  assign n41829 = ~n42755 ^ n42753;
  assign n41830 = ~BUF2_REG_26__SCAN_IN;
  assign n41835 = ~n42802 & ~n41830;
  assign n41833 = ~n42804 | ~n41831;
  assign n41832 = ~n43698 | ~P2_EAX_REG_26__SCAN_IN;
  assign n41834 = ~n41833 | ~n41832;
  assign n41837 = ~n41835 & ~n41834;
  assign n41836 = ~n43690 | ~BUF1_REG_26__SCAN_IN;
  assign n41838 = ~n41837 | ~n41836;
  assign P2_U2893 = ~n41841 | ~n41840;
  assign n41843 = n43525 | P2_EBX_REG_26__SCAN_IN;
  assign P2_U2861 = ~n41846 | ~n41845;
  assign n41847 = ~n42400 & ~n42184;
  assign n41861 = ~n42171 | ~P1_REIP_REG_21__SCAN_IN;
  assign n41897 = ~n42185 & ~n41848;
  assign n41849 = ~P1_REIP_REG_20__SCAN_IN | ~n41897;
  assign n41853 = ~n42507 | ~n43559;
  assign n41851 = ~n43796 | ~P1_EBX_REG_21__SCAN_IN;
  assign n41850 = ~n43797 | ~P1_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n41852 = n41851 & n41850;
  assign P1_U2819 = ~n41861 | ~n41860;
  assign n41868 = ~n42135 | ~n41862;
  assign P3_U2674 = ~n41868 | ~n41867;
  assign n41870 = ~n43897 & ~n41916;
  assign n41892 = ~n41870 | ~n41869;
  assign n41887 = ~n43847 & ~n41931;
  assign n41871 = ~n41873 & ~P2_EBX_REG_30__SCAN_IN;
  assign n41885 = ~n43836 | ~n41934;
  assign n41878 = ~n41877 | ~P2_EBX_REG_31__SCAN_IN;
  assign n41883 = ~n41879 & ~n41878;
  assign n41881 = ~n41920 | ~P2_REIP_REG_31__SCAN_IN;
  assign n41880 = ~n41921 | ~P2_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n41882 = ~n41881 | ~n41880;
  assign n41884 = ~n41883 & ~n41882;
  assign n41890 = n41887 | n41886;
  assign P2_U2824 = ~n41892 | ~n41891;
  assign n41895 = ~n41894 | ~n41893;
  assign n41911 = ~n41895 | ~P1_REIP_REG_20__SCAN_IN;
  assign n41909 = ~n41897 | ~n41896;
  assign n41903 = ~n43796 | ~P1_EBX_REG_20__SCAN_IN;
  assign n41901 = n43797 & P1_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n41900 = ~n42175 & ~n41899;
  assign P1_U2820 = ~n41911 | ~n41910;
  assign n41915 = ~n41912 | ~n43808;
  assign n41914 = ~n41913;
  assign n41917 = ~n41915 | ~n41914;
  assign n41918 = ~n41917 | ~n41916;
  assign n41925 = ~n41919 & ~n41918;
  assign n41923 = ~n41920 | ~P2_REIP_REG_29__SCAN_IN;
  assign n41922 = ~n41921 | ~P2_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n41924 = ~n41923 | ~n41922;
  assign n41948 = ~n41925 & ~n41924;
  assign n41929 = ~n41928 | ~n41927;
  assign n43756 = ~n41930 | ~n41929;
  assign n41937 = ~n43753 | ~n41934;
  assign P2_U2826 = ~n41948 | ~n41947;
  assign n41950 = ~n42501 & ~n43462;
  assign n41961 = n41968 | n43358;
  assign n41970 = ~n43469 | ~P1_REIP_REG_19__SCAN_IN;
  assign n41954 = ~n43709 | ~P1_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n41957 = n41970 & n41954;
  assign n41956 = ~n43362 | ~n41955;
  assign P1_U2980 = ~n41961 | ~n41960;
  assign n42582 = ~n42364 & ~n41962;
  assign n41967 = n42582 | P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n42967 = ~n42539;
  assign n41964 = ~n41963 & ~n42967;
  assign n41966 = ~n42584 | ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n41975 = ~n41967 | ~n41966;
  assign n41971 = ~n43344 | ~n41969;
  assign P1_U3012 = ~n41975 | ~n41974;
  assign n42825 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN | ~n42365;
  assign n43337 = ~n42828 & ~n42825;
  assign n41978 = ~n41976 & ~n43337;
  assign n43350 = ~n43337 | ~n42919;
  assign n41982 = ~n41979 | ~n43350;
  assign n41980 = ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n41981 = ~n43351 & ~n41980;
  assign n41983 = ~n41982 | ~n41981;
  assign n41984 = ~n41983 | ~n42539;
  assign n41985 = ~n42538;
  assign n41987 = ~n41985 | ~P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n42544 = ~P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n42921 = ~P1_INSTADDRPOINTER_REG_25__SCAN_IN | ~n43337;
  assign n41986 = ~n42544 | ~n42537;
  assign n42010 = ~n41987 | ~n41986;
  assign n41993 = ~n41989 & ~n41988;
  assign n41991 = ~P1_INSTADDRPOINTER_REG_18__SCAN_IN | ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n41992 = ~n41991 & ~n41990;
  assign n41994 = ~n41993 | ~n41992;
  assign n41997 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN & ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n41996 = ~P1_INSTADDRPOINTER_REG_24__SCAN_IN & ~P1_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n41998 = ~n41997 | ~n41996;
  assign n42000 = ~n41999 & ~n41998;
  assign n42001 = n43462 | n42000;
  assign n42548 = ~n42546 | ~n42004;
  assign n42005 = ~n43462 ^ P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign P1_U3004 = ~n42010 | ~n42009;
  assign n42014 = ~n42012 & ~n42011;
  assign P3_U2996 = ~n42027 | ~n42026;
  assign n42031 = ~n43306 | ~n42029;
  assign n42030 = ~n43737 | ~BUF1_REG_25__SCAN_IN;
  assign n42035 = ~n42031 | ~n42030;
  assign n42033 = ~n43738 | ~DATAI_25_;
  assign n42032 = ~n43732 | ~P1_EAX_REG_25__SCAN_IN;
  assign n42034 = ~n42033 | ~n42032;
  assign n42036 = ~n42035 & ~n42034;
  assign P1_U2879 = ~n42037 | ~n42036;
  assign n42039 = ~n42833 | ~n44021;
  assign n42038 = ~n44023 | ~P1_EBX_REG_24__SCAN_IN;
  assign P1_U2848 = ~n42041 | ~n42040;
  assign n42045 = ~n43306 | ~n42043;
  assign n42044 = ~n43737 | ~BUF1_REG_24__SCAN_IN;
  assign n42049 = ~n42045 | ~n42044;
  assign n42047 = ~n43738 | ~DATAI_24_;
  assign n42046 = ~n43732 | ~P1_EAX_REG_24__SCAN_IN;
  assign n42048 = ~n42047 | ~n42046;
  assign n42050 = ~n42049 & ~n42048;
  assign P1_U2880 = ~n42051 | ~n42050;
  assign n42053 = ~n42052 | ~n42130;
  assign P3_U2672 = ~n42057 | ~n42056;
  assign n42060 = ~n42561 | ~n43809;
  assign n42080 = n42060 | n42562;
  assign n42078 = ~n43911 & ~n42061;
  assign n42065 = n42062 | P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n42067 = n42089 & P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n42068 = ~n42067 & ~n42085;
  assign n42072 = ~n43813 | ~n42565;
  assign n42071 = n43540 | n42070;
  assign n42074 = ~n42072 | ~n42071;
  assign n42566 = ~n43880 | ~P2_REIP_REG_11__SCAN_IN;
  assign n42073 = ~n42566;
  assign n42075 = ~n42074 & ~n42073;
  assign P2_U3003 = ~n42080 | ~n42079;
  assign n42087 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n42082 = ~n42081 | ~n42087;
  assign n42088 = ~n42104 | ~n42087;
  assign n42101 = n42201 | n42100;
  assign n42102 = ~n42101 | ~n42198;
  assign n42116 = ~n43886 & ~n42140;
  assign n42141 = ~n43880 | ~P2_REIP_REG_13__SCAN_IN;
  assign n42108 = ~n42557 & ~n42104;
  assign n42702 = n42105 & n42108;
  assign n42106 = ~n42702;
  assign n42107 = ~n42106 & ~n42303;
  assign n42112 = ~n43159 & ~n42107;
  assign n43150 = ~n42109 | ~n42108;
  assign n42300 = ~n42112 & ~n42700;
  assign n42113 = ~n43158 | ~n42303;
  assign n42650 = ~n42300 | ~n42113;
  assign n42114 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN | ~n42650;
  assign n42115 = ~n42141 | ~n42114;
  assign n42119 = ~n42116 & ~n42115;
  assign n42118 = ~n43583 | ~n42117;
  assign n42124 = n42119 & n42118;
  assign n42120 = ~n43150;
  assign n42123 = ~n42303 & ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n42648 = ~n42727 | ~n42123;
  assign P2_U3033 = ~n42128 | ~n42127;
  assign n42136 = ~n42135 | ~n42134;
  assign P3_U2673 = ~n42137 | ~n42136;
  assign n42144 = ~n43915 & ~n42140;
  assign n42142 = ~n43917 | ~P2_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n42143 = ~n42142 | ~n42141;
  assign n42148 = ~n42144 & ~n42143;
  assign n42146 = ~n42145;
  assign n42147 = ~n43896 | ~n42146;
  assign P2_U3001 = ~n42152 | ~n42151;
  assign n42170 = ~n43803 | ~n43343;
  assign n42159 = ~n43796 | ~P1_EBX_REG_25__SCAN_IN;
  assign n42154 = ~n43797 | ~P1_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n42153 = ~n42400 | ~P1_REIP_REG_25__SCAN_IN;
  assign n42157 = ~n42154 | ~n42153;
  assign n42155 = ~n43035;
  assign n42156 = ~n42175 & ~n42155;
  assign n42158 = ~n42157 & ~n42156;
  assign n42163 = ~n42160;
  assign n42162 = ~n42161 & ~P1_REIP_REG_25__SCAN_IN;
  assign n42164 = n42163 | n42162;
  assign n42165 = ~n42185 & ~n42164;
  assign n42167 = n42166 | n42165;
  assign P1_U2815 = ~n42170 | ~n42169;
  assign n42179 = ~n43796 | ~P1_EBX_REG_22__SCAN_IN;
  assign n42177 = n43797 & P1_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n42176 = ~n42175 & ~n42174;
  assign n42187 = ~n42185 & ~n42184;
  assign n42188 = ~n42187 | ~n42186;
  assign P1_U2818 = ~n42191 | ~n42190;
  assign n42651 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n42192 = ~n42214;
  assign n42193 = ~n42192 & ~n42700;
  assign n42195 = ~n42193 & ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n42194 = ~n42699 & ~n42626;
  assign n42597 = ~n42700 & ~n42194;
  assign n42230 = n42195 | n42597;
  assign n42200 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN & ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n42210 = ~n42240;
  assign n42211 = ~n42210 | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n42216 = ~n42702 | ~n42214;
  assign n42217 = ~n42216 | ~n42215;
  assign n42595 = ~n42702 | ~n42626;
  assign n42218 = n42217 & n42595;
  assign n42221 = ~n43148 | ~n42218;
  assign n42220 = ~n43583 | ~n42219;
  assign n42222 = ~n43767 | ~n42424;
  assign n42425 = ~n43880 | ~P2_REIP_REG_15__SCAN_IN;
  assign n42223 = ~n42222 | ~n42425;
  assign P2_U3031 = ~n42230 | ~n42229;
  assign n42601 = ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n42231 = ~n42601 & ~n42628;
  assign n42291 = ~n42626 | ~n42231;
  assign n42232 = ~n42291;
  assign n42271 = n42234 | n42233;
  assign n42381 = ~n42238 | ~n42237;
  assign n42239 = ~P2_INSTADDRPOINTER_REG_15__SCAN_IN & ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n42241 = ~n42381 & ~n42385;
  assign n42251 = ~n42242 | ~n42241;
  assign n42261 = ~n42260;
  assign n42267 = ~n42261 | ~n43896;
  assign n42262 = ~n42616;
  assign n42265 = ~n42262 & ~n43915;
  assign n42263 = ~n43917 | ~P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n42613 = ~n43880 | ~P2_REIP_REG_17__SCAN_IN;
  assign n42264 = ~n42263 | ~n42613;
  assign n42266 = ~n42265 & ~n42264;
  assign P2_U2997 = ~n42271 | ~n42270;
  assign n42272 = ~n42524 | ~n42702;
  assign n42274 = ~n43148 | ~n42272;
  assign n42273 = ~n43158 | ~n42291;
  assign n42275 = ~n42274 | ~n42273;
  assign n42299 = n42527 | n42282;
  assign n42286 = ~n42348 | ~n42347;
  assign n42290 = ~n42439 & ~n43886;
  assign n42440 = ~n43880 | ~P2_REIP_REG_18__SCAN_IN;
  assign n42292 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN & ~n42291;
  assign P2_U3028 = ~n42299 | ~n42298;
  assign n42302 = ~n42300 | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n42301 = ~n42652 | ~n42303;
  assign n42317 = ~n42302 | ~n42301;
  assign n42306 = ~n42305 ^ P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n42313 = ~n42451 | ~n43876;
  assign n42308 = ~n43767 | ~n42452;
  assign n42453 = ~n43880 | ~P2_REIP_REG_12__SCAN_IN;
  assign n42311 = ~n42308 | ~n42453;
  assign n42310 = ~n43877 & ~n42309;
  assign n42312 = ~n42311 & ~n42310;
  assign P2_U3034 = ~n42317 | ~n42316;
  assign n42328 = ~n42321 | ~n42320;
  assign n42326 = ~n42322 & ~P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign P3_U2835 = ~n42342 | ~n42341;
  assign n42350 = ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n42698 = ~n42524 | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n42363 = n42869 | n43924;
  assign n42361 = ~n43911 & ~n42345;
  assign n42349 = ~n42347 | ~n42346;
  assign n42357 = ~n42871 & ~n43915;
  assign n42355 = n43540 | n42354;
  assign n42873 = ~n43880 | ~P2_REIP_REG_19__SCAN_IN;
  assign n42356 = ~n42355 | ~n42873;
  assign P2_U2995 = ~n42363 | ~n42362;
  assign n42366 = ~n42364 & ~n43335;
  assign n42368 = ~n42366 | ~n42365;
  assign n42370 = ~n42368 | ~n42367;
  assign n42369 = ~n42825 | ~n42539;
  assign n42377 = ~n42370 | ~n42829;
  assign P1_U3008 = ~n42377 | ~n42376;
  assign n42399 = n42380 | n42604;
  assign n42384 = ~n42382 & ~n42381;
  assign n42389 = ~n42637;
  assign n42392 = ~n42389 & ~n43915;
  assign n42390 = ~n43917 | ~P2_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n42634 = ~n43880 | ~P2_REIP_REG_16__SCAN_IN;
  assign n42391 = ~n42390 | ~n42634;
  assign n42395 = ~n42392 & ~n42391;
  assign n42394 = n43911 | n42393;
  assign P2_U2998 = ~n42399 | ~n42398;
  assign n42402 = ~n42400 | ~P1_REIP_REG_23__SCAN_IN;
  assign n42401 = ~n43796 | ~P1_EBX_REG_23__SCAN_IN;
  assign n42421 = ~n42402 | ~n42401;
  assign n42407 = ~n42403 & ~P1_REIP_REG_23__SCAN_IN;
  assign n42406 = ~n42405 | ~n42404;
  assign n42419 = ~n42407 & ~n42406;
  assign n42413 = ~n43797 | ~P1_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n42411 = ~n42410;
  assign n42420 = n42419 | n42418;
  assign P1_U2817 = n42421 | n42420;
  assign n42428 = ~n43813 | ~n42424;
  assign n42426 = ~n43917 | ~P2_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n42427 = n42426 & n42425;
  assign n42430 = ~n43911 & ~n42429;
  assign P2_U2999 = n42435 | n42434;
  assign n42445 = ~n42438 | ~n43896;
  assign n42443 = ~n42439 & ~n43915;
  assign n42441 = ~n43917 | ~P2_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n42442 = ~n42441 | ~n42440;
  assign n42444 = ~n42443 & ~n42442;
  assign P2_U2996 = n42449 | n42448;
  assign n42456 = ~n43813 | ~n42452;
  assign n42454 = ~n43917 | ~P2_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n42455 = n42454 & n42453;
  assign n42459 = ~n42456 | ~n42455;
  assign n42458 = ~n43911 & ~n42457;
  assign n42460 = ~n42459 & ~n42458;
  assign P2_U3002 = n42463 | n42462;
  assign n42478 = ~n42473 | ~n43896;
  assign n42476 = ~n42516 & ~n43915;
  assign n42474 = ~n43917 | ~P2_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n42518 = ~n43880 | ~P2_REIP_REG_20__SCAN_IN;
  assign n42475 = ~n42474 | ~n42518;
  assign P2_U2994 = ~n42482 | ~n42481;
  assign n42497 = ~n42538 | ~P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n42484 = ~n22933 | ~n42544;
  assign n42485 = ~n42546 & ~n42484;
  assign n43043 = ~n43033 & ~n42488;
  assign n42489 = n42544 ^ P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n42490 = ~n42489 & ~n42537;
  assign n42493 = ~n43043 & ~n42490;
  assign P1_U3003 = ~n42497 | ~n42496;
  assign n42502 = ~n42501 & ~n42500;
  assign n42513 = n42679 | n43358;
  assign n42681 = ~n43469 | ~P1_REIP_REG_21__SCAN_IN;
  assign n42506 = ~n43709 | ~P1_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n42509 = n42681 & n42506;
  assign n42508 = ~n42507 | ~n43362;
  assign P1_U2978 = ~n42513 | ~n42512;
  assign n42521 = ~n42516 & ~n43886;
  assign n42523 = ~n42727 | ~n42522;
  assign n42530 = ~n42523 | ~n42697;
  assign n42525 = ~n42524 | ~n42727;
  assign n42884 = ~P2_INSTADDRPOINTER_REG_19__SCAN_IN & ~n42525;
  assign n42528 = ~n42884 & ~n42868;
  assign n42529 = ~P2_INSTADDRPOINTER_REG_20__SCAN_IN | ~n42528;
  assign n42531 = ~n42530 | ~n42529;
  assign P2_U3026 = ~n42536 | ~n42535;
  assign n42542 = P1_INSTADDRPOINTER_REG_29__SCAN_IN | n42965;
  assign n43463 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n42541 = ~n43463 & ~n42538;
  assign n42540 = ~n42539 | ~n42547;
  assign n42543 = ~P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n42545 = ~n42544 | ~n42543;
  assign n42972 = ~n42546 & ~n42545;
  assign n43449 = ~n42549 & ~n42971;
  assign n42550 = ~n43462 & ~n43463;
  assign P1_U3002 = ~n42556 | ~n42555;
  assign n42559 = ~n42557 & ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n42578 = ~n42559 | ~n42558;
  assign n42576 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN | ~n42560;
  assign n42567 = ~n43767 | ~n42565;
  assign n42570 = ~n42567 | ~n42566;
  assign n42569 = ~n43877 & ~n42568;
  assign n42571 = ~n42570 & ~n42569;
  assign P2_U3035 = ~n42578 | ~n42577;
  assign n42581 = ~n42580 & ~n42579;
  assign n42594 = ~n42582 | ~n42581;
  assign n42583 = ~P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n42591 = n42590 | n42589;
  assign P1_U3011 = ~n42594 | ~n42593;
  assign n42596 = ~n43148 | ~n42595;
  assign n42602 = ~n42600 & ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n42603 = ~n42602 & ~n42601;
  assign n42605 = ~n42626 | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n42606 = ~n42652 & ~n42605;
  assign n42607 = ~n42606 & ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n42615 = ~n43877 & ~n42612;
  assign n42614 = ~n42613;
  assign n42618 = ~n42615 & ~n42614;
  assign n42617 = ~n43767 | ~n42616;
  assign P2_U3029 = ~n42622 | ~n42621;
  assign n42636 = ~n43877 & ~n42633;
  assign n42635 = ~n42634;
  assign n42639 = ~n42636 & ~n42635;
  assign n42638 = ~n43767 | ~n42637;
  assign P2_U3030 = ~n42643 | ~n42642;
  assign n42644 = ~n44023 | ~P1_EBX_REG_26__SCAN_IN;
  assign P1_U2846 = ~n42647 | ~n42646;
  assign n42649 = ~n42648 | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n42655 = ~n42650 & ~n42649;
  assign n42653 = ~n42652 & ~n42651;
  assign n42654 = ~n42653 & ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n42674 = n42655 | n42654;
  assign n42663 = ~n42662 ^ P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n42666 = ~n43583 | ~n42665;
  assign n42843 = ~n43880 | ~P2_REIP_REG_14__SCAN_IN;
  assign n42667 = ~n43886 & ~n42842;
  assign P2_U3032 = ~n42674 | ~n42673;
  assign n42678 = ~n42826 | ~n42675;
  assign n42677 = ~n42676 | ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n42686 = ~n42678 | ~n42677;
  assign P1_U3010 = ~n42686 | ~n42685;
  assign n42690 = ~n43306 | ~n42688;
  assign n42689 = ~n43737 | ~BUF1_REG_26__SCAN_IN;
  assign n42694 = ~n42690 | ~n42689;
  assign n42692 = ~n43738 | ~DATAI_26_;
  assign n42691 = ~n43732 | ~P1_EAX_REG_26__SCAN_IN;
  assign n42693 = ~n42692 | ~n42691;
  assign n42695 = ~n42694 & ~n42693;
  assign P1_U2878 = ~n42696 | ~n42695;
  assign n43152 = ~n42698 & ~n42697;
  assign n42701 = ~n43152 & ~n42699;
  assign n42704 = ~n42701 & ~n42700;
  assign n43147 = ~n43152 | ~n42702;
  assign n42703 = ~n43148 | ~n43147;
  assign n42735 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN | ~n42894;
  assign n42993 = ~n42720 & ~n42719;
  assign n42726 = ~n42857 & ~n43886;
  assign n42724 = ~n42723 | ~n43583;
  assign n42858 = ~n43880 | ~P2_REIP_REG_21__SCAN_IN;
  assign n42729 = n42726 | n42725;
  assign n42728 = ~n42892 & ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign P2_U3025 = ~n42735 | ~n42734;
  assign n42738 = ~n43306 | ~n42736;
  assign n42737 = ~n43737 | ~BUF1_REG_27__SCAN_IN;
  assign n42742 = ~n42738 | ~n42737;
  assign n42740 = ~n43738 | ~DATAI_27_;
  assign n42739 = ~n43732 | ~P1_EAX_REG_27__SCAN_IN;
  assign n42741 = ~n42740 | ~n42739;
  assign n42743 = ~n42742 & ~n42741;
  assign P1_U2877 = ~n42744 | ~n42743;
  assign n42752 = ~n42746 | ~n42745;
  assign n42751 = ~n42750 | ~n42749;
  assign n43059 = ~n42755 | ~n42754;
  assign n42757 = ~n43500 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n42756 = ~n43483 | ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n42761 = ~n42757 | ~n42756;
  assign n42759 = ~n22911 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n42758 = ~n43495 | ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n42760 = ~n42759 | ~n42758;
  assign n42767 = ~n42761 & ~n42760;
  assign n42762 = ~n43499 | ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n42765 = ~n42762 | ~n43509;
  assign n42763 = ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n42764 = ~n43514 & ~n42763;
  assign n42766 = ~n42765 & ~n42764;
  assign n42771 = ~n42767 | ~n42766;
  assign n42769 = ~n43503 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n42768 = ~n43496 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n42770 = ~n42769 | ~n42768;
  assign n42795 = ~n42771 & ~n42770;
  assign n42772 = ~n43495 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n42775 = ~n42772 | ~n43490;
  assign n42773 = ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n42774 = ~n43514 & ~n42773;
  assign n42781 = ~n42775 & ~n42774;
  assign n42776 = ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n42779 = ~n43408 & ~n42776;
  assign n42777 = ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n42778 = ~n22927 & ~n42777;
  assign n42780 = ~n42779 & ~n42778;
  assign n42793 = ~n42781 | ~n42780;
  assign n42785 = ~n43092 & ~n42782;
  assign n42784 = ~n43094 & ~n42783;
  assign n42791 = ~n42785 & ~n42784;
  assign n42789 = ~n43098 & ~n42786;
  assign n42788 = ~n43100 & ~n42787;
  assign n42790 = ~n42789 & ~n42788;
  assign n42792 = ~n42791 | ~n42790;
  assign n42794 = ~n42793 & ~n42792;
  assign n43060 = ~n42795 & ~n42794;
  assign n42797 = ~n43059 ^ n43060;
  assign n42798 = ~n43060 | ~n43061;
  assign n43058 = ~n42799 & ~n42798;
  assign n42808 = ~n42802 & ~n42801;
  assign n42806 = ~n42804 | ~n42803;
  assign n42805 = ~n43698 | ~P2_EAX_REG_27__SCAN_IN;
  assign n42807 = ~n42806 | ~n42805;
  assign n42810 = ~n42808 & ~n42807;
  assign n42809 = ~n43690 | ~BUF1_REG_27__SCAN_IN;
  assign n42811 = ~n42810 | ~n42809;
  assign P2_U2892 = ~n42814 | ~n42813;
  assign n42816 = ~n43709 | ~P1_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n42819 = n42817 & n42816;
  assign n42818 = ~n43362 | ~n43378;
  assign P1_U2972 = ~n42824 | ~n42823;
  assign n42827 = ~n42826 & ~n42825;
  assign n42831 = ~n42827 & ~P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n42830 = ~n42829 & ~n42828;
  assign n42839 = n42831 | n42830;
  assign P1_U3007 = ~n42839 | ~n42838;
  assign n42846 = ~n43915 & ~n42842;
  assign n42844 = ~n43917 | ~P2_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n42845 = ~n42844 | ~n42843;
  assign n42849 = n42846 | n42845;
  assign n42848 = ~n43911 & ~n42847;
  assign P2_U3000 = n42853 | n42852;
  assign n42863 = ~n42856 & ~n43911;
  assign n42861 = ~n42857 & ~n43915;
  assign n42859 = ~n43917 | ~P2_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n42860 = ~n42859 | ~n42858;
  assign n42862 = n42861 | n42860;
  assign P2_U2993 = n42867 | n42866;
  assign P2_U3027 = n42884 | n42883;
  assign n42886 = n43525 | P2_EBX_REG_27__SCAN_IN;
  assign P2_U2860 = ~n42889 | ~n42888;
  assign n43010 = ~n42992 & ~n42892;
  assign n42890 = ~n43010 | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n42896 = ~n42906 | ~n42890;
  assign n42996 = ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n42891 = ~n42992 & ~n42996;
  assign n42893 = ~n42892 & ~n42891;
  assign n42895 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN | ~n43012;
  assign n42918 = ~n42896 | ~n42895;
  assign n42903 = ~n42993 & ~n43173;
  assign n42902 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN & ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n43206 = ~n42903 & ~n43182;
  assign n42912 = ~n42953 & ~n43886;
  assign n42910 = ~n42909 | ~n43583;
  assign n42954 = ~n43880 | ~P2_REIP_REG_23__SCAN_IN;
  assign P2_U3023 = ~n42918 | ~n42917;
  assign n42920 = ~n42919;
  assign n42923 = ~n42921 & ~n42920;
  assign n43352 = ~n42923 & ~n42922;
  assign n42925 = ~n42924 | ~n43350;
  assign n42926 = ~n43352 & ~n43329;
  assign n42929 = ~n42926 | ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n42928 = ~n42927 & ~P1_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n42932 = ~n42929 & ~n42928;
  assign n42931 = ~n42930 & ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n42940 = n42932 | n42931;
  assign P1_U3005 = ~n42940 | ~n42939;
  assign n42944 = ~n43306 | ~n42942;
  assign n42943 = ~n43737 | ~BUF1_REG_28__SCAN_IN;
  assign n42948 = ~n42944 | ~n42943;
  assign n42946 = ~n43738 | ~DATAI_28_;
  assign n42945 = ~n43732 | ~P1_EAX_REG_28__SCAN_IN;
  assign n42947 = ~n42946 | ~n42945;
  assign n42949 = ~n42948 & ~n42947;
  assign P1_U2876 = ~n42950 | ~n42949;
  assign n42964 = n42951 | n43924;
  assign n42957 = ~n42953 & ~n43915;
  assign n42955 = ~n43917 | ~P2_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n42956 = ~n42955 | ~n42954;
  assign n42961 = ~n42960 & ~n43911;
  assign P2_U2991 = ~n42964 | ~n42963;
  assign n43461 = ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n42970 = ~n43447 | ~n43461;
  assign n43438 = ~n42967 | ~n42966;
  assign n42968 = ~n43437 | ~n43438;
  assign n42969 = ~n42968 | ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n42984 = n43441 | n43569;
  assign P1_U3001 = ~n42988 | ~n42987;
  assign n42991 = ~n43181 | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n42994 = ~n42993 | ~n42992;
  assign n43005 = ~n43000 | ~n43896;
  assign n43003 = ~n43015 & ~n43915;
  assign n43001 = ~n43917 | ~P2_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n43017 = ~n43880 | ~P2_REIP_REG_22__SCAN_IN;
  assign n43002 = ~n43001 | ~n43017;
  assign P2_U2992 = n43009 | n43008;
  assign n43011 = ~n43010 & ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n43026 = n43012 | n43011;
  assign n43020 = ~n43015 & ~n43886;
  assign P2_U3024 = ~n43026 | ~n43025;
  assign n43041 = n43342 | n43358;
  assign n43034 = n43709 & P1_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n43345 = ~n43033 & ~n43032;
  assign n43037 = ~n43034 & ~n43345;
  assign n43036 = ~n43362 | ~n43035;
  assign P1_U2974 = ~n43041 | ~n43040;
  assign n43045 = ~n43043;
  assign n43044 = ~n43709 | ~P1_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n43048 = ~n43045 | ~n43044;
  assign n43047 = ~n43713 & ~n43046;
  assign n43049 = n43048 | n43047;
  assign P1_U2971 = ~n43053 | ~n43052;
  assign n43064 = ~n43059;
  assign n43062 = ~n43060;
  assign n43063 = ~n43062 & ~n43061;
  assign n43393 = ~n43064 | ~n43063;
  assign n43066 = ~n43483 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n43065 = ~n43496 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n43070 = ~n43066 | ~n43065;
  assign n43068 = ~n43503 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n43067 = ~n43499 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n43069 = ~n43068 | ~n43067;
  assign n43076 = ~n43070 & ~n43069;
  assign n43071 = ~n22911 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n43074 = ~n43071 | ~n43509;
  assign n43073 = ~n43408 & ~n43072;
  assign n43075 = ~n43074 & ~n43073;
  assign n43080 = ~n43076 | ~n43075;
  assign n43078 = ~n43484 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n43077 = ~n43495 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n43079 = ~n43078 | ~n43077;
  assign n43108 = ~n43080 & ~n43079;
  assign n43081 = ~n43495 | ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n43084 = ~n43081 | ~n43490;
  assign n43083 = ~n43514 & ~n43082;
  assign n43090 = ~n43084 & ~n43083;
  assign n43088 = ~n43408 & ~n43085;
  assign n43087 = ~n22927 & ~n43086;
  assign n43089 = ~n43088 & ~n43087;
  assign n43106 = ~n43090 | ~n43089;
  assign n43096 = ~n43092 & ~n43091;
  assign n43095 = ~n43094 & ~n43093;
  assign n43104 = ~n43096 & ~n43095;
  assign n43102 = ~n43098 & ~n43097;
  assign n43101 = ~n43100 & ~n43099;
  assign n43103 = ~n43102 & ~n43101;
  assign n43105 = ~n43104 | ~n43103;
  assign n43107 = ~n43106 & ~n43105;
  assign n43391 = ~n43108 & ~n43107;
  assign n43110 = ~n43689 | ~BUF2_REG_28__SCAN_IN;
  assign n43109 = ~n43690 | ~BUF1_REG_28__SCAN_IN;
  assign n43115 = ~n43110 | ~n43109;
  assign n43113 = n43697 | n43111;
  assign n43112 = ~n43698 | ~P2_EAX_REG_28__SCAN_IN;
  assign n43114 = ~n43113 | ~n43112;
  assign n43116 = n43115 | n43114;
  assign P2_U2891 = ~n43119 | ~n43118;
  assign n43123 = ~n43306 | ~n43121;
  assign n43122 = ~n43737 | ~BUF1_REG_29__SCAN_IN;
  assign n43127 = ~n43123 | ~n43122;
  assign n43125 = ~n43738 | ~DATAI_29_;
  assign n43124 = ~n43732 | ~P1_EAX_REG_29__SCAN_IN;
  assign n43126 = ~n43125 | ~n43124;
  assign n43128 = ~n43127 & ~n43126;
  assign P1_U2875 = ~n43129 | ~n43128;
  assign n43131 = n43525 | P2_EBX_REG_28__SCAN_IN;
  assign P2_U2859 = ~n43134 | ~n43133;
  assign n43136 = ~n43709 | ~P1_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n43140 = n43137 & n43136;
  assign n43139 = ~n43362 | ~n43138;
  assign P1_U2970 = ~n43145 | ~n43144;
  assign n43187 = ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n43149 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN | ~n43146;
  assign n43160 = ~n43149 & ~n43147;
  assign n43151 = ~n43150 & ~n43149;
  assign n43157 = ~n43152 | ~n43151;
  assign n43153 = ~n43157;
  assign n43163 = ~n43158 | ~n43157;
  assign n43161 = ~n43160 & ~n43159;
  assign n43162 = ~n43164 & ~n43161;
  assign n43226 = ~n43613 & ~n43549;
  assign n43757 = ~n43165 & ~n43164;
  assign n43166 = ~n43226 & ~n43757;
  assign n43580 = ~n43578 & ~n43166;
  assign n43169 = ~n43580 | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n43167 = ~n43617 | ~n43612;
  assign n43168 = ~n43167 | ~n43599;
  assign n43205 = ~n43169 | ~n43168;
  assign n43191 = ~n43181 | ~n43180;
  assign n43197 = n43196 | n43877;
  assign n43318 = ~n43880 | ~P2_REIP_REG_26__SCAN_IN;
  assign P2_U3020 = ~n43205 | ~n43204;
  assign n43532 = ~n43210 | ~n43209;
  assign n43214 = ~n43224 & ~n43915;
  assign n43212 = ~n43917 | ~P2_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n43228 = ~n43880 | ~P2_REIP_REG_24__SCAN_IN;
  assign n43213 = ~n43212 | ~n43228;
  assign n43218 = n43217 & n43896;
  assign P2_U2990 = ~n43221 | ~n43220;
  assign n43234 = ~n43224 & ~n43886;
  assign n43232 = ~n43225 | ~n43583;
  assign n43227 = ~n43617 & ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n43230 = ~n43227 & ~n43226;
  assign n43229 = ~n43228;
  assign n43231 = ~n43230 & ~n43229;
  assign P2_U3022 = n43238 | n43237;
  assign n43285 = ~n43240 & ~n43239;
  assign n43244 = ~n43241 | ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n43243 = ~n43242 | ~P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n43250 = ~n43244 | ~n43243;
  assign n43248 = ~n43245 | ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n43247 = ~n43246 | ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n43249 = ~n43248 | ~n43247;
  assign n43259 = ~n43250 & ~n43249;
  assign n43253 = ~n22907 | ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n43252 = ~n43251 | ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n43257 = ~n43253 | ~n43252;
  assign n43255 = ~n22908 | ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n43254 = ~n22915 | ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n43256 = ~n43255 | ~n43254;
  assign n43258 = ~n43257 & ~n43256;
  assign n43283 = ~n43259 | ~n43258;
  assign n43263 = ~n43260 | ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n43262 = ~n43261 | ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n43269 = ~n43263 | ~n43262;
  assign n43267 = ~n43264 | ~P1_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n43266 = ~n43265 | ~P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n43268 = ~n43267 | ~n43266;
  assign n43281 = ~n43269 & ~n43268;
  assign n43273 = ~n43270 | ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n43272 = ~n43271 | ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n43279 = ~n43273 | ~n43272;
  assign n43277 = ~n43274 | ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n43276 = ~n43275 | ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n43278 = ~n43277 | ~n43276;
  assign n43280 = ~n43279 & ~n43278;
  assign n43282 = ~n43281 | ~n43280;
  assign n43284 = ~n43283 & ~n43282;
  assign n43287 = n43285 ^ n43284;
  assign n43292 = n43287 | n43286;
  assign n43289 = ~n43721 | ~P1_EAX_REG_30__SCAN_IN;
  assign n43288 = ~P1_PHYADDRPOINTER_REG_30__SCAN_IN | ~n43722;
  assign n43290 = ~n43289 | ~n43288;
  assign n43291 = ~n43290 & ~n43294;
  assign n43296 = ~n43292 | ~n43291;
  assign n43299 = ~P1_EBX_REG_30__SCAN_IN;
  assign n43301 = ~n43300 & ~n43299;
  assign P1_U2842 = ~n43304 | ~n43303;
  assign n43308 = ~n43306 | ~n43305;
  assign n43307 = ~n43737 | ~BUF1_REG_30__SCAN_IN;
  assign n43312 = ~n43308 | ~n43307;
  assign n43310 = ~n43738 | ~DATAI_30_;
  assign n43309 = ~n43732 | ~P1_EAX_REG_30__SCAN_IN;
  assign n43311 = ~n43310 | ~n43309;
  assign n43313 = ~n43312 & ~n43311;
  assign P1_U2874 = ~n43314 | ~n43313;
  assign n43319 = ~n43917 | ~P2_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n43320 = ~n43319 | ~n43318;
  assign n43327 = ~n43326 | ~n43896;
  assign P2_U2988 = ~n43328 | ~n43327;
  assign n43340 = n43329 | n43351;
  assign n43332 = ~n43331 & ~n43330;
  assign n43334 = ~n43333 & ~n43332;
  assign n43336 = ~n43335 & ~n43334;
  assign n43338 = ~n43337 | ~n43336;
  assign n43339 = ~n43338 | ~n43351;
  assign n43357 = ~n43340 | ~n43339;
  assign n43349 = ~n43342 & ~n43341;
  assign n43346 = ~n43345;
  assign n43355 = ~n43349 & ~n43348;
  assign n43353 = ~n43351 | ~n43350;
  assign n43354 = ~n43353 | ~n43352;
  assign n43356 = n43355 & n43354;
  assign P1_U3006 = ~n43357 | ~n43356;
  assign n43360 = ~n43709 | ~P1_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n43364 = n43361 & n43360;
  assign n43363 = ~n43362 | ~n43558;
  assign P1_U2969 = ~n43370 | ~n43369;
  assign n43388 = ~n43371 | ~P1_REIP_REG_27__SCAN_IN;
  assign n43373 = ~P1_REIP_REG_26__SCAN_IN | ~n43372;
  assign n43375 = ~n43796 | ~P1_EBX_REG_27__SCAN_IN;
  assign n43381 = ~n43380 & ~n43379;
  assign n43385 = n43384 | n43383;
  assign P1_U2813 = ~n43388 | ~n43387;
  assign n43395 = ~n43390 & ~n43389;
  assign n43392 = ~n43391;
  assign n43397 = ~n22911 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n43396 = ~n43495 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n43406 = ~n43397 | ~n43396;
  assign n43399 = ~n43496 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n43398 = ~n43499 | ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n43403 = ~n43399 | ~n43398;
  assign n43401 = ~n43503 | ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n43400 = ~n43484 | ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n43402 = ~n43401 | ~n43400;
  assign n43404 = ~n43403 & ~n43402;
  assign n43405 = ~n43490 | ~n43404;
  assign n43413 = ~n43406 & ~n43405;
  assign n43411 = ~n43408 & ~n43407;
  assign n43410 = ~n22927 & ~n43409;
  assign n43412 = ~n43411 & ~n43410;
  assign n43432 = ~n43413 | ~n43412;
  assign n43415 = ~n43503 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n43414 = ~n43495 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n43424 = ~n43415 | ~n43414;
  assign n43417 = ~n43496 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n43416 = ~n43500 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n43421 = ~n43417 | ~n43416;
  assign n43419 = ~n43499 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n43418 = ~n22911 | ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n43420 = ~n43419 | ~n43418;
  assign n43422 = ~n43421 & ~n43420;
  assign n43423 = ~n43509 | ~n43422;
  assign n43430 = ~n43424 & ~n43423;
  assign n43428 = ~n22927 & ~n43425;
  assign n43427 = ~n43514 & ~n43426;
  assign n43429 = ~n43428 & ~n43427;
  assign n43431 = ~n43430 | ~n43429;
  assign n43433 = ~n43525 & ~P2_EBX_REG_29__SCAN_IN;
  assign n43435 = n43434 | n43433;
  assign P2_U2858 = ~n43436 | ~n43435;
  assign n43440 = ~n43461 & ~n43437;
  assign n43439 = ~P1_INSTADDRPOINTER_REG_31__SCAN_IN | ~n43438;
  assign n43445 = ~P1_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n43446 = ~P1_INSTADDRPOINTER_REG_30__SCAN_IN | ~n43445;
  assign n43450 = ~P1_INSTADDRPOINTER_REG_30__SCAN_IN & ~P1_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n43451 = ~n43462 & ~n43450;
  assign n43452 = ~n43453 & ~n43451;
  assign n43460 = ~n43452 & ~n43456;
  assign n43454 = ~n22933 & ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n43458 = ~n43455 & ~n43454;
  assign n43457 = ~n43456;
  assign n43459 = ~n43458 & ~n43457;
  assign n43468 = ~n43460 & ~n43459;
  assign n43465 = ~n43462 & ~n43461;
  assign n43464 = ~n43463 & ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n43466 = ~n43465 & ~n43464;
  assign n43467 = ~n43466 & ~P1_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n43708 = ~n43468 & ~n43467;
  assign n43470 = ~n43708 | ~n36906;
  assign n43471 = ~n43470 | ~n43711;
  assign n43473 = ~n43472 & ~n43471;
  assign P1_U3000 = ~n43474 | ~n43473;
  assign n43478 = ~n22911 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n43477 = ~n43503 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n43494 = n43478 & n43477;
  assign n43480 = ~n43495 | ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n43479 = ~n43496 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n43492 = ~n43480 | ~n43479;
  assign n43482 = ~n43499 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n43481 = ~n43500 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n43488 = ~n43482 | ~n43481;
  assign n43486 = ~n43483 | ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n43485 = ~n43484 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n43487 = ~n43486 | ~n43485;
  assign n43489 = ~n43488 & ~n43487;
  assign n43491 = ~n43490 | ~n43489;
  assign n43493 = ~n43492 & ~n43491;
  assign n43520 = ~n43494 | ~n43493;
  assign n43498 = ~n43495 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n43497 = ~n43496 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n43511 = ~n43498 | ~n43497;
  assign n43502 = ~n43499 | ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n43501 = ~n43500 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n43507 = ~n43502 | ~n43501;
  assign n43505 = ~n22911 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n43504 = ~n43503 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n43506 = ~n43505 | ~n43504;
  assign n43508 = ~n43507 & ~n43506;
  assign n43510 = ~n43509 | ~n43508;
  assign n43518 = ~n43511 & ~n43510;
  assign n43516 = ~n22927 & ~n43512;
  assign n43513 = ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n43515 = ~n43514 & ~n43513;
  assign n43517 = ~n43516 & ~n43515;
  assign n43519 = ~n43518 | ~n43517;
  assign n43521 = ~n43520 | ~n43519;
  assign n43526 = n43525 | P2_EBX_REG_30__SCAN_IN;
  assign P2_U2857 = ~n43529 | ~n43528;
  assign n43541 = n43540 | n43539;
  assign n43585 = ~n43880 | ~P2_REIP_REG_25__SCAN_IN;
  assign n43542 = ~n43541 | ~n43585;
  assign n43553 = n43552 | n43591;
  assign P2_U2989 = ~n43554 | ~n43553;
  assign n43556 = ~n43796 | ~P1_EBX_REG_30__SCAN_IN;
  assign n43555 = ~n43797 | ~P1_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n43563 = ~n43556 | ~n43555;
  assign n43557 = ~P1_REIP_REG_30__SCAN_IN & ~n43564;
  assign n43561 = ~n43557 | ~n43788;
  assign n43560 = ~n43559 | ~n43558;
  assign n43562 = ~n43561 | ~n43560;
  assign n43789 = ~n43565 & ~n43564;
  assign n43568 = n43566 | n43789;
  assign n43574 = ~n43573 & ~n43572;
  assign n43576 = n43575 & n43574;
  assign P1_U2810 = ~n43577 | ~n43576;
  assign n43579 = ~n43578 & ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n43596 = n43580 | n43579;
  assign n43588 = ~n43582 & ~n43886;
  assign P2_U3021 = ~n43596 | ~n43595;
  assign n43601 = ~n43597;
  assign n43600 = ~n43661 & ~n43599;
  assign n43746 = ~n43601 | ~n43600;
  assign n43658 = ~n43605 | ~n43604;
  assign n43608 = ~n43658 | ~n43606;
  assign n43665 = ~n43658 | ~n43657;
  assign n43610 = ~n43609 | ~n43665;
  assign n43624 = n43611 | n43877;
  assign n43615 = ~n43612 | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n43614 = ~n43613 & ~n43615;
  assign n43759 = ~n43614 & ~n43757;
  assign n43620 = ~n43759 & ~n43661;
  assign n43616 = ~n43615;
  assign n43618 = ~n43853;
  assign n43619 = ~n43618 & ~P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n43622 = ~n43620 & ~n43619;
  assign n43646 = ~n43880 | ~P2_REIP_REG_27__SCAN_IN;
  assign n43621 = ~n43646;
  assign n43623 = ~n43622 & ~n43621;
  assign P2_U3019 = n43630 | n43629;
  assign n43632 = ~BUF2_REG_29__SCAN_IN | ~n43689;
  assign n43631 = ~n43690 | ~BUF1_REG_29__SCAN_IN;
  assign n43642 = ~n43632 | ~n43631;
  assign n43636 = n43697 | n43634;
  assign n43635 = ~n43698 | ~P2_EAX_REG_29__SCAN_IN;
  assign n43637 = ~n43636 | ~n43635;
  assign P2_U2890 = n43642 | n43641;
  assign n43647 = ~n43917 | ~P2_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n43648 = ~n43647 | ~n43646;
  assign n43655 = n43654 | n43911;
  assign P2_U2987 = ~n43656 | ~n43655;
  assign n43688 = n43775 | n43893;
  assign n43664 = ~n43658 & ~n43657;
  assign n43666 = ~n43665;
  assign n43760 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n43674 = ~n43760;
  assign n43673 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN & ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n43675 = n43674 | n43673;
  assign n43677 = ~n43853 & ~n43675;
  assign n43778 = ~n43880 | ~P2_REIP_REG_28__SCAN_IN;
  assign n43676 = ~n43778;
  assign n43679 = ~n43677 & ~n43676;
  assign n43678 = ~n43759 | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n43680 = ~n43679 | ~n43678;
  assign n43683 = ~n43682 | ~n43767;
  assign P2_U3018 = ~n43688 | ~n43687;
  assign n43692 = ~n43689 | ~BUF2_REG_30__SCAN_IN;
  assign n43691 = ~n43690 | ~BUF1_REG_30__SCAN_IN;
  assign n43706 = ~n43692 | ~n43691;
  assign n43704 = ~n43694 | ~n43693;
  assign n43700 = n43697 | n43696;
  assign n43699 = ~n43698 | ~P2_EAX_REG_30__SCAN_IN;
  assign n43701 = ~n43700 | ~n43699;
  assign P2_U2889 = n43706 | n43705;
  assign n43710 = ~n43709 | ~P1_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n43715 = ~n43711 | ~n43710;
  assign n43714 = ~n43713 & ~n43712;
  assign n43724 = ~n43721 | ~P1_EAX_REG_31__SCAN_IN;
  assign n43723 = ~P1_PHYADDRPOINTER_REG_31__SCAN_IN | ~n43722;
  assign n43726 = ~n43724 | ~n43723;
  assign n43730 = ~n43795 & ~n43729;
  assign P1_U2968 = n43731 | n43730;
  assign n43733 = ~n43795 & ~n32238;
  assign n43736 = ~n43733 & ~n43732;
  assign n43742 = ~n43736 & ~n43735;
  assign n43740 = ~n43737 | ~BUF1_REG_31__SCAN_IN;
  assign n43739 = ~n43738 | ~DATAI_31_;
  assign P1_U2873 = n43742 | n43741;
  assign n43745 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n43892 = ~n43746 & ~n43745;
  assign n43810 = ~n43747 & ~n43892;
  assign n43752 = ~n43750 | ~n43749;
  assign n43827 = ~n43752 | ~n43751;
  assign n43825 = ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n43851 = ~n43825 & ~n43760;
  assign n43758 = ~n43757 & ~n43851;
  assign n43879 = ~n43759 & ~n43758;
  assign n43761 = ~n43853 & ~n43760;
  assign n43762 = ~n43761 & ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n43764 = ~n43879 & ~n43762;
  assign n43815 = ~n43880 | ~P2_REIP_REG_29__SCAN_IN;
  assign n43763 = ~n43815;
  assign n43765 = n43764 | n43763;
  assign n43768 = ~n43814 | ~n43767;
  assign P2_U3017 = ~n43773 | ~n43772;
  assign n43787 = ~n43774 | ~n43896;
  assign n43779 = ~n43917 | ~P2_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n43780 = ~n43779 | ~n43778;
  assign P2_U2986 = ~n43787 | ~n43786;
  assign n43790 = ~n43789 | ~n43788;
  assign n43793 = n43790 & n29669;
  assign n43792 = ~n43791 & ~n29669;
  assign n43801 = ~n43795 & ~n43794;
  assign n43799 = ~n43796 | ~P1_EBX_REG_31__SCAN_IN;
  assign n43798 = ~n43797 | ~P1_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n43805 = ~n43801 & ~n43800;
  assign P1_U2809 = n43807 | n43806;
  assign n43824 = ~n43808 & ~n43911;
  assign n43816 = ~n43917 | ~P2_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n43817 = n43816 & n43815;
  assign P2_U2985 = n43824 | n43823;
  assign n43831 = ~n43827 & ~n43826;
  assign n43873 = ~n43831 & ~n43830;
  assign n43839 = ~n43873 | ~n43870;
  assign n43846 = ~n43839 | ~n43838;
  assign n43841 = ~n43873;
  assign n43869 = ~n43841 | ~n43871;
  assign n43845 = ~n43869 | ~n43844;
  assign n43860 = n43847 | n43877;
  assign n43848 = ~n43891 | ~n43851;
  assign n43881 = n43853 | n43848;
  assign n43849 = ~n43881 | ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n43856 = ~n43850 & ~n43849;
  assign n43852 = ~P2_INSTADDRPOINTER_REG_30__SCAN_IN | ~n43851;
  assign n43854 = ~n43853 & ~n43852;
  assign n43855 = ~n43854 & ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n43858 = ~n43856 & ~n43855;
  assign n43918 = ~n43880 | ~P2_REIP_REG_31__SCAN_IN;
  assign n43857 = ~n43918;
  assign n43859 = ~n43858 & ~n43857;
  assign n43862 = ~n43860 | ~n43859;
  assign n43863 = ~n43862 & ~n43861;
  assign n43865 = ~n43892 | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign P2_U3015 = n43867 | n43866;
  assign n43875 = n43869 | n43868;
  assign n43874 = ~n43873 | ~n43872;
  assign n43890 = ~n43898 | ~n43876;
  assign n43885 = n43878 | n43877;
  assign n43883 = ~n43879 & ~n43891;
  assign n43900 = ~n43880 | ~P2_REIP_REG_30__SCAN_IN;
  assign n43882 = ~n43881 | ~n43900;
  assign n43884 = ~n43883 & ~n43882;
  assign n43906 = n43892 ^ n43891;
  assign P2_U3016 = n43895 | n43894;
  assign n43910 = ~n43897 | ~n43896;
  assign n43901 = ~n43917 | ~P2_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n43902 = ~n43901 | ~n43900;
  assign n43908 = ~n43905 | ~n43904;
  assign P2_U2984 = ~n43910 | ~n43909;
  assign n43929 = n43912 | n43911;
  assign n43923 = ~n43914 | ~n43913;
  assign n43919 = ~n43917 | ~P2_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n43920 = ~n43919 | ~n43918;
  assign n43926 = ~n43925 & ~n43924;
  assign n43928 = ~n43927 & ~n43926;
  assign P2_U2983 = ~n43929 | ~n43928;
  assign n43936 = ~n43931 & ~n43930;
  assign n43934 = ~P3_EBX_REG_2__SCAN_IN & ~n43932;
  assign n43935 = ~n43934 & ~n43933;
  assign P3_U2701 = n43936 | n43935;
  assign n43941 = ~n43937 & ~n43982;
  assign n43939 = ~P3_DATAO_REG_29__SCAN_IN | ~n43984;
  assign n43938 = ~P3_UWORD_REG_13__SCAN_IN | ~n32190;
  assign n43940 = ~n43939 | ~n43938;
  assign P3_U2738 = n43941 | n43940;
  assign n43946 = ~n43942 & ~n43982;
  assign n43944 = ~P3_DATAO_REG_27__SCAN_IN | ~n43984;
  assign n43943 = ~P3_UWORD_REG_11__SCAN_IN | ~n32190;
  assign n43945 = ~n43944 | ~n43943;
  assign P3_U2740 = n43946 | n43945;
  assign n43951 = ~n43947 & ~n43982;
  assign n43949 = ~P3_DATAO_REG_25__SCAN_IN | ~n43984;
  assign n43948 = ~P3_UWORD_REG_9__SCAN_IN | ~n32190;
  assign n43950 = ~n43949 | ~n43948;
  assign P3_U2742 = n43951 | n43950;
  assign n43956 = ~n43952 & ~n43982;
  assign n43954 = ~P3_DATAO_REG_24__SCAN_IN | ~n43984;
  assign n43953 = ~P3_UWORD_REG_8__SCAN_IN | ~n32190;
  assign n43955 = ~n43954 | ~n43953;
  assign P3_U2743 = n43956 | n43955;
  assign n43961 = ~n43957 & ~n43982;
  assign n43959 = ~P3_DATAO_REG_23__SCAN_IN | ~n43984;
  assign n43958 = ~P3_UWORD_REG_7__SCAN_IN | ~n32190;
  assign n43960 = ~n43959 | ~n43958;
  assign P3_U2744 = n43961 | n43960;
  assign n43966 = ~n43962 & ~n43982;
  assign n43964 = ~P3_DATAO_REG_22__SCAN_IN | ~n43984;
  assign n43963 = ~P3_UWORD_REG_6__SCAN_IN | ~n32190;
  assign n43965 = ~n43964 | ~n43963;
  assign P3_U2745 = n43966 | n43965;
  assign n43971 = ~n43967 & ~n43982;
  assign n43969 = ~P3_DATAO_REG_21__SCAN_IN | ~n43984;
  assign n43968 = ~P3_UWORD_REG_5__SCAN_IN | ~n32190;
  assign n43970 = ~n43969 | ~n43968;
  assign P3_U2746 = n43971 | n43970;
  assign n43976 = ~n43972 & ~n43982;
  assign n43974 = ~P3_DATAO_REG_20__SCAN_IN | ~n43984;
  assign n43973 = ~P3_UWORD_REG_4__SCAN_IN | ~n32190;
  assign n43975 = ~n43974 | ~n43973;
  assign P3_U2747 = n43976 | n43975;
  assign n43981 = ~n43977 & ~n43982;
  assign n43979 = ~P3_DATAO_REG_18__SCAN_IN | ~n43984;
  assign n43978 = ~P3_UWORD_REG_2__SCAN_IN | ~n32190;
  assign n43980 = ~n43979 | ~n43978;
  assign P3_U2749 = n43981 | n43980;
  assign n43988 = ~n43983 & ~n43982;
  assign n43986 = ~P3_DATAO_REG_17__SCAN_IN | ~n43984;
  assign n43985 = ~P3_UWORD_REG_1__SCAN_IN | ~n32190;
  assign n43987 = ~n43986 | ~n43985;
  assign P3_U2750 = n43988 | n43987;
  assign n43999 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n43989;
  assign n43991 = ~n43990 | ~n43994;
  assign n43997 = ~n43991 | ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n43995 = ~n43993 & ~n43992;
  assign n43996 = ~n43995 | ~n43994;
  assign n43998 = ~n43997 | ~n43996;
  assign P3_U2864 = n43999 | n43998;
  assign n44001 = ~n44003;
  assign n44006 = ~n44001 & ~n44000;
  assign n44004 = ~n44002 & ~P2_READREQUEST_REG_SCAN_IN;
  assign n44005 = ~n44004 & ~n44003;
  assign P2_U3612 = n44006 | n44005;
  assign n44010 = ~n44008 | ~n44021;
  assign n44009 = ~P1_EBX_REG_10__SCAN_IN | ~n44023;
  assign n44011 = ~n44010 | ~n44009;
  assign P1_U2862 = n44012 | n44011;
  assign n44018 = ~n44013 & ~n44019;
  assign n44016 = ~n44014 | ~n44021;
  assign n44015 = ~P1_EBX_REG_6__SCAN_IN | ~n44023;
  assign n44017 = ~n44016 | ~n44015;
  assign P1_U2866 = n44018 | n44017;
  assign n44027 = ~n44020 & ~n44019;
  assign n44025 = ~n44022 | ~n44021;
  assign n44024 = ~P1_EBX_REG_2__SCAN_IN | ~n44023;
  assign n44026 = ~n44025 | ~n44024;
  assign P1_U2870 = n44027 | n44026;
  assign n44033 = ~n44029 & ~n44091;
  assign n44031 = ~P1_DATAO_REG_15__SCAN_IN | ~n44092;
  assign n44030 = ~n44093 | ~P1_LWORD_REG_15__SCAN_IN;
  assign n44032 = ~n44031 | ~n44030;
  assign P1_U2921 = n44033 | n44032;
  assign n44038 = ~n44034 & ~n44091;
  assign n44036 = ~P1_DATAO_REG_14__SCAN_IN | ~n44092;
  assign n44035 = ~n44093 | ~P1_LWORD_REG_14__SCAN_IN;
  assign n44037 = ~n44036 | ~n44035;
  assign P1_U2922 = n44038 | n44037;
  assign n44043 = ~n44039 & ~n44091;
  assign n44041 = ~P1_DATAO_REG_12__SCAN_IN | ~n44092;
  assign n44040 = ~n44093 | ~P1_LWORD_REG_12__SCAN_IN;
  assign n44042 = ~n44041 | ~n44040;
  assign P1_U2924 = n44043 | n44042;
  assign n44048 = ~n44044 & ~n44091;
  assign n44046 = ~P1_DATAO_REG_10__SCAN_IN | ~n44092;
  assign n44045 = ~n44093 | ~P1_LWORD_REG_10__SCAN_IN;
  assign n44047 = ~n44046 | ~n44045;
  assign P1_U2926 = n44048 | n44047;
  assign n44053 = ~n44049 & ~n44091;
  assign n44051 = ~P1_DATAO_REG_9__SCAN_IN | ~n44092;
  assign n44050 = ~n44093 | ~P1_LWORD_REG_9__SCAN_IN;
  assign n44052 = ~n44051 | ~n44050;
  assign P1_U2927 = n44053 | n44052;
  assign n44058 = ~n44054 & ~n44091;
  assign n44056 = ~P1_DATAO_REG_8__SCAN_IN | ~n44092;
  assign n44055 = ~n44093 | ~P1_LWORD_REG_8__SCAN_IN;
  assign n44057 = ~n44056 | ~n44055;
  assign P1_U2928 = n44058 | n44057;
  assign n44062 = ~n24862 & ~n44091;
  assign n44060 = ~P1_DATAO_REG_7__SCAN_IN | ~n44092;
  assign n44059 = ~n44093 | ~P1_LWORD_REG_7__SCAN_IN;
  assign n44061 = ~n44060 | ~n44059;
  assign P1_U2929 = n44062 | n44061;
  assign n44067 = ~n44063 & ~n44091;
  assign n44065 = ~P1_DATAO_REG_6__SCAN_IN | ~n44092;
  assign n44064 = ~n44093 | ~P1_LWORD_REG_6__SCAN_IN;
  assign n44066 = ~n44065 | ~n44064;
  assign P1_U2930 = n44067 | n44066;
  assign n44072 = ~n44068 & ~n44091;
  assign n44070 = ~P1_DATAO_REG_5__SCAN_IN | ~n44092;
  assign n44069 = ~n44093 | ~P1_LWORD_REG_5__SCAN_IN;
  assign n44071 = ~n44070 | ~n44069;
  assign P1_U2931 = n44072 | n44071;
  assign n44077 = ~n44073 & ~n44091;
  assign n44075 = ~P1_DATAO_REG_4__SCAN_IN | ~n44092;
  assign n44074 = ~n44093 | ~P1_LWORD_REG_4__SCAN_IN;
  assign n44076 = ~n44075 | ~n44074;
  assign P1_U2932 = n44077 | n44076;
  assign n44081 = ~n24818 & ~n44091;
  assign n44079 = ~P1_DATAO_REG_3__SCAN_IN | ~n44092;
  assign n44078 = ~n44093 | ~P1_LWORD_REG_3__SCAN_IN;
  assign n44080 = ~n44079 | ~n44078;
  assign P1_U2933 = n44081 | n44080;
  assign n44085 = ~n24788 & ~n44091;
  assign n44083 = ~P1_DATAO_REG_2__SCAN_IN | ~n44092;
  assign n44082 = ~n44093 | ~P1_LWORD_REG_2__SCAN_IN;
  assign n44084 = ~n44083 | ~n44082;
  assign P1_U2934 = n44085 | n44084;
  assign n44090 = ~n44086 & ~n44091;
  assign n44088 = ~P1_DATAO_REG_1__SCAN_IN | ~n44092;
  assign n44087 = ~n44093 | ~P1_LWORD_REG_1__SCAN_IN;
  assign n44089 = ~n44088 | ~n44087;
  assign P1_U2935 = n44090 | n44089;
  assign n44097 = ~n24804 & ~n44091;
  assign n44095 = ~P1_DATAO_REG_0__SCAN_IN | ~n44092;
  assign n44094 = ~n44093 | ~P1_LWORD_REG_0__SCAN_IN;
  assign n44096 = ~n44095 | ~n44094;
  assign P1_U2936 = n44097 | n44096;
  assign n44101 = ~n44099;
  assign n44103 = ~n44101 & ~n44100;
  assign n44104 = ~n44103 & ~n44102;
  assign n44110 = ~n44105 & ~n44104;
  assign n44108 = ~n44106 | ~P1_STATE2_REG_1__SCAN_IN;
  assign n44109 = ~n44108 | ~n44107;
  assign P1_U3162 = n44110 | n44109;
endmodule


