// Benchmark "c3540_lock" written by ABC on Thu May 13 23:37:40 2021

module c3540_lock ( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G405  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G405;
  wire n1542, n1692, n1686, n1705, n1696, n1697, n1704, n1643, n1655, n1220,
    n920, n1257, n1657, n1452, n951, n1458, n875, n1530, n932, n1224,
    n1163, n876, n1713, n883, n892, n886, n880, n879, n884, n877, n878,
    n900, n881, n891, n890, n1687, n1306, n882, n898, n889, n888, n885,
    n1693, n887, n896, n894, n893, n895, n897, n899, n915, n1736, n1380,
    n1559, n1473, n901, n909, n903, n902, n907, n905, n904, n906, n908,
    n913, n911, n910, n912, n914, n916, n918, n1691, n1466, n1446, n917,
    n919, n960, n925, n1168, n1074, n921, n999, n1126, n1175, n1004, n924,
    n922, n1120, n923, n929, n1123, n927, n938, n1171, n926, n928, n953,
    n930, n936, n1133, n1153, n1296, n931, n1015, n1151, n1073, n933, n935,
    n1154, n934, n942, n1157, n940, n937, n1158, n939, n941, n946, n944,
    n945, n1164, n943, n955, n1118, n1273, n948, n947, n949, n950, n1191,
    n952, n1276, n1749, n954, n958, n956, n957, n1349, n959, n1203, n962,
    n961, n966, n964, n1176, n963, n965, n982, n975, n984, n967, n971,
    n969, n1131, n968, n970, n973, n972, n978, n977, n979, n974, n976,
    n983, n981, n980, n985, n1117, n1192, n987, n986, n1411, n1265, n1343,
    n1533, n989, n988, n996, n1016, n992, n1063, n991, n990, n994, n1068,
    n993, n995, n1010, n998, n1099, n997, n1009, n1003, n1001, n1000,
    n1077, n1002, n1006, n1005, n1008, n1007, n1236, n1237, n1012, n1011,
    n1013, n1014, n1515, n1019, n1017, n1018, n1023, n1021, n1020, n1022,
    n1025, n1024, n1096, n1027, n1093, n1026, n1538, n1028, n1029, n1463,
    n1653, n1246, n1031, n1030, n1033, n1032, n1035, n1034, n1535, n1113,
    n1037, n1036, n1038, n1039, n1589, n1040, n1044, n1042, n1041, n1043,
    n1046, n1045, n1098, n1054, n1049, n1047, n1048, n1051, n1050, n1053,
    n1052, n1240, n1056, n1055, n1509, n1059, n1057, n1058, n1060, n1061,
    n1241, n1062, n1067, n1065, n1064, n1066, n1070, n1069, n1097, n1072,
    n1085, n1071, n1084, n1076, n1075, n1081, n1254, n1079, n1078, n1080,
    n1083, n1082, n1524, n1110, n1541, n1087, n1086, n1088, n1089, n1544,
    n1090, n1091, n1235, n1107, n1092, n1094, n1095, n1104, n1101, n1100,
    n1102, n1103, n1105, n1106, n1269, n1251, n1350, n1111, n1108, n1245,
    n1109, n1532, n1112, n1739, n1195, n1250, n1115, n1114, n1272, n1116,
    n1361, n1119, n1148, n1167, n1453, n1122, n1121, n1130, n1125, n1124,
    n1128, n1231, n1127, n1129, n1258, n1132, n1137, n1135, n1134, n1136,
    n1139, n1138, n1142, n1141, n1143, n1140, n1261, n1149, n1277, n1145,
    n1144, n1146, n1147, n1259, n1150, n1188, n1152, n1156, n1155, n1162,
    n1160, n1159, n1161, n1183, n1166, n1182, n1165, n1337, n1174, n1170,
    n1169, n1173, n1172, n1180, n1738, n1178, n1177, n1179, n1181, n1189,
    n1334, n1185, n1184, n1186, n1187, n1335, n1190, n1742, n1197, n1194,
    n1193, n1268, n1196, n1282, n1740, n1198, n1404, n1199, n1201, n1200,
    n1202, G381, n1664, n1228, n1227, n1459, n1229, n1230, n1552, n1232,
    n1661, n1233, n1234, n1634, n1510, n1239, n1238, n1505, n1242, n1244,
    n1243, n1716, n1512, n1547, n1527, n1525, n1519, n1467, n1640, n1656,
    n1333, n1260, n1264, n1262, n1263, n1396, n1266, n1267, n1342, n1275,
    n1274, n1348, n1279, n1278, n1345, n1443, n1330, n1658, n1297, n1298,
    n1332, n1300, n1299, n1304, n1302, n1301, n1303, n1310, n1562, n1305,
    n1308, n1472, n1307, n1309, n1311, n1328, n1313, n1312, n1317, n1315,
    n1314, n1316, n1325, n1319, n1318, n1323, n1321, n1320, n1322, n1324,
    n1326, n1327, n1329, n1331, n1341, n1336, n1339, n1338, n1346, n1340,
    n1360, n1344, n1347, n1357, n1521, n1352, n1351, n1353, n1406, n1354,
    n1355, n1356, n1358, n1721, n1359, G375, n1363, n1362, n1364, n1403,
    n1366, n1365, n1379, n1368, n1367, n1369, n1377, n1371, n1370, n1375,
    n1373, n1372, n1374, n1376, n1378, n1394, n1414, n1673, n1382, n1381,
    n1390, n1384, n1383, n1388, n1604, n1385, n1386, n1387, n1389, n1391,
    n1392, n1393, n1395, n1398, n1397, n1399, n1401, n1400, n1402, n1409,
    n1405, n1407, n1408, G378, n1410, n1451, n1445, n1413, n1412, n1418,
    n1416, n1415, n1417, n1426, n1420, n1419, n1424, n1422, n1421, n1423,
    n1425, n1441, n1428, n1427, n1432, n1601, n1430, n1429, n1431, n1439,
    n1677, n1433, n1437, n1435, n1434, n1436, n1438, n1440, n1442, n1444,
    n1448, n1447, n1449, n1450, G384, n1717, n1669, n1735, n1455, n1454,
    n1456, n1457, n1461, n1460, n1462, n1663, n1465, n1464, n1469, n1468,
    n1470, n1504, n1581, n1471, n1484, n1474, n1482, n1476, n1475, n1480,
    n1478, n1477, n1479, n1481, n1483, n1501, n1486, n1485, n1487, n1495,
    n1489, n1488, n1493, n1491, n1490, n1492, n1494, n1499, n1497, n1496,
    n1498, n1500, n1502, n1503, n1507, n1590, n1506, n1508, n1518, n1511,
    n1513, n1514, n1641, n1516, n1517, n1523, n1520, n1649, n1522, G393,
    n1543, n1526, n1528, n1650, n1644, n1529, n1531, n1551, n1534, n1536,
    n1537, n1540, n1539, n1549, n1546, n1545, n1630, n1548, n1550, n1597,
    n1554, n1553, n1555, n1594, n1557, n1556, n1569, n1558, n1567, n1561,
    n1560, n1565, n1563, n1564, n1566, n1568, n1570, n1571, n1588, n1573,
    n1572, n1577, n1575, n1574, n1576, n1585, n1579, n1578, n1583, n1580,
    n1582, n1584, n1586, n1587, n1592, n1591, n1593, n1595, n1596, G387,
    n1599, n1598, n1612, n1600, n1610, n1603, n1602, n1608, n1606, n1605,
    n1607, n1609, n1611, n1628, n1674, n1613, n1614, n1622, n1616, n1615,
    n1620, n1618, n1617, n1619, n1621, n1626, n1624, n1623, n1625, n1627,
    n1629, n1632, n1631, n1633, n1639, n1636, n1635, n1637, n1638, n1648,
    n1642, n1646, n1645, n1647, n1652, n1651, G390, G355, n1654, n1723,
    n1660, n1659, n1668, n1662, n1666, n1665, n1667, n1670, n1715, n1672,
    n1671, n1685, n1675, n1683, n1676, n1681, n1679, n1678, n1680, n1682,
    n1684, n1711, n1689, n1688, n1690, n1703, n1695, n1694, n1701, n1699,
    n1698, n1700, n1702, n1709, n1707, n1706, n1708, n1710, n1712, n1714,
    n1719, n1718, n1720, n1722, G396, n1724, n1733, n1727, n1725, n1726,
    n1732, n1728, n1729, n1731, n1730, n1734, G405_Lock, keyinput_0,
    keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5, keyinput_6,
    keyinput_7, keyinput_8, keyinput_9, keyinput_10, keyinput_11,
    keyinput_12, keyinput_13, keyinput_14, keyinput_15, keyinput_16,
    keyinput_17, keyinput_18, keyinput_19, keyinput_20, keyinput_21,
    keyinput_22, keyinput_23, keyinput_24, keyinput_25, keyinput_26,
    keyinput_27, keyinput_28, keyinput_29, keyinput_30, keyinput_31,
    keyinput_32, keyinput_33, keyinput_34, keyinput_35, keyinput_36,
    keyinput_37, keyinput_38, keyinput_39, keyinput_40, keyinput_41,
    keyinput_42, keyinput_43, keyinput_44, keyinput_45, keyinput_46,
    keyinput_47, keyinput_48, keyinput_49, keyinput_50, keyinput_51,
    keyinput_52, keyinput_53, keyinput_54, keyinput_55, keyinput_56,
    keyinput_57, keyinput_58, keyinput_59, keyinput_60, keyinput_61,
    keyinput_62, keyinput_63, input_0, input_1, AND_1, input_2, OR_2,
    input_3, AND_3, input_4, OR_4, input_5, OR_5, input_6, OR_6, input_7,
    AND_7, input_8, OR_8, input_9, OR_9, input_10, AND_10, input_11,
    AND_11, input_12, AND_12, input_13, OR_13, input_14, OR_14, input_15,
    AND_15, input_16, AND_16, input_17, OR_17, input_18, OR_18, input_19,
    OR_19, input_20, OR_20, input_21, AND_21, input_22, AND_22, input_23,
    OR_23, input_24, OR_24, input_25, AND_25, input_26, OR_26, input_27,
    AND_27, input_28, AND_28, input_29, OR_29, input_30, AND_30, input_31,
    OR_31, input_32, input_33, AND_33, input_34, OR_34, input_35, AND_35,
    input_36, OR_36, input_37, OR_37, input_38, OR_38, input_39, AND_39,
    input_40, OR_40, input_41, OR_41, input_42, AND_42, input_43, AND_43,
    input_44, AND_44, input_45, OR_45, input_46, OR_46, input_47, AND_47,
    input_48, AND_48, input_49, OR_49, input_50, OR_50, input_51, OR_51,
    input_52, OR_52, input_53, AND_53, input_54, AND_54, input_55, OR_55,
    input_56, OR_56, input_57, AND_57, input_58, OR_58, input_59, AND_59,
    input_60, AND_60, input_61, OR_61, input_62, AND_62, input_63, OR_63,
    OR_63_INV, CASOP;
  assign n1542 = ~n1276 & ~n1749;
  assign n1692 = ~n892 & ~n889;
  assign n1686 = ~G200 & ~n880;
  assign n1705 = ~n884 & ~n877;
  assign n1696 = ~n892 & ~n891;
  assign n1697 = ~n890 & ~n889;
  assign n1704 = ~n883 & ~n880;
  assign n1643 = ~G41 & ~n1657;
  assign n1655 = ~n1643 & ~n1530;
  assign n1220 = ~G20 | ~G1;
  assign n920 = ~n1220;
  assign n1257 = ~G13;
  assign n1657 = ~n920 | ~n1257;
  assign n1452 = ~G20;
  assign n951 = ~n1452 | ~G13;
  assign n1458 = ~G45;
  assign n875 = n951 | n1458;
  assign n1530 = ~G1 | ~n875;
  assign n932 = ~G13 | ~G1;
  assign n1224 = ~n932;
  assign n1163 = ~G169;
  assign n876 = ~G20 | ~n1163;
  assign n1713 = ~n1224 | ~n876;
  assign n883 = ~G200;
  assign n892 = ~G20 | ~G179;
  assign n886 = ~n1452 & ~G190;
  assign n880 = n892 | n886;
  assign n879 = ~G132 | ~n1704;
  assign n884 = ~G20 | ~G200;
  assign n877 = ~G190 | ~n892;
  assign n878 = ~n1705 | ~G159;
  assign n900 = ~n879 | ~n878;
  assign n881 = ~n1686 | ~G137;
  assign n891 = ~G200 | ~n886;
  assign n890 = ~n892;
  assign n1687 = ~n891 & ~n890;
  assign n1306 = ~G58 | ~n1687;
  assign n882 = ~n881 | ~n1306;
  assign n898 = ~G33 & ~n882;
  assign n889 = ~n886 | ~n883;
  assign n888 = ~n1692 | ~G150;
  assign n885 = ~n892 | ~n884;
  assign n1693 = ~n886 & ~n885;
  assign n887 = ~n1693 | ~G50;
  assign n896 = ~n888 | ~n887;
  assign n894 = ~n1697 | ~G128;
  assign n893 = ~n1696 | ~G143;
  assign n895 = ~n894 | ~n893;
  assign n897 = ~n896 & ~n895;
  assign n899 = ~n898 | ~n897;
  assign n915 = ~n900 & ~n899;
  assign n1736 = ~G77;
  assign n1380 = ~n1687;
  assign n1559 = ~n1736 & ~n1380;
  assign n1473 = ~G87 | ~n1693;
  assign n901 = ~G33 | ~n1473;
  assign n909 = ~n1559 & ~n901;
  assign n903 = ~G283 | ~n1686;
  assign n902 = ~G294 | ~n1704;
  assign n907 = ~n903 | ~n902;
  assign n905 = ~G303 | ~n1697;
  assign n904 = ~G116 | ~n1696;
  assign n906 = ~n905 | ~n904;
  assign n908 = ~n907 & ~n906;
  assign n913 = ~n909 | ~n908;
  assign n911 = ~n1705 | ~G97;
  assign n910 = ~n1692 | ~G107;
  assign n912 = ~n911 | ~n910;
  assign n914 = ~n913 & ~n912;
  assign n916 = ~n915 & ~n914;
  assign n918 = ~n1713 & ~n916;
  assign n1691 = ~G33;
  assign n1466 = ~n1257 | ~n1691;
  assign n1446 = ~n1466 | ~n1713;
  assign n917 = ~G68 & ~n1446;
  assign n919 = ~n918 & ~n917;
  assign n960 = ~n1655 | ~n919;
  assign n925 = ~G1 & ~n1452;
  assign n1168 = ~G13 | ~n925;
  assign n1074 = ~n1168;
  assign n921 = ~n920 | ~G33;
  assign n999 = ~n932 | ~n921;
  assign n1126 = ~G20 | ~n999;
  assign n1175 = ~n1126;
  assign n1004 = ~n1074 & ~n1175;
  assign n924 = n1004 | G68;
  assign n922 = ~G33 | ~n1224;
  assign n1120 = ~G20 & ~n922;
  assign n923 = ~n1120 | ~G77;
  assign n929 = ~n924 | ~n923;
  assign n1123 = ~n925 & ~n999;
  assign n927 = ~n1123 | ~G68;
  assign n938 = ~n1224 | ~n1691;
  assign n1171 = ~G20 & ~n938;
  assign n926 = ~G50 | ~n1171;
  assign n928 = ~n927 | ~n926;
  assign n953 = n929 | n928;
  assign n930 = ~G41 & ~G45;
  assign n936 = ~G1 & ~n930;
  assign n1133 = ~G274 | ~n936;
  assign n1153 = ~n1133;
  assign n1296 = ~G41;
  assign n931 = ~n1296 & ~n1691;
  assign n1015 = ~n932 & ~n931;
  assign n1151 = ~G33 | ~n1015;
  assign n1073 = ~G97;
  assign n933 = ~n1151 & ~n1073;
  assign n935 = ~n1153 & ~n933;
  assign n1154 = ~G1698 & ~n938;
  assign n934 = ~n1154 | ~G226;
  assign n942 = ~n935 | ~n934;
  assign n1157 = ~n1015 & ~n936;
  assign n940 = ~n1157 | ~G238;
  assign n937 = ~G1698;
  assign n1158 = ~n938 & ~n937;
  assign n939 = ~G232 | ~n1158;
  assign n941 = ~n940 | ~n939;
  assign n946 = ~n942 & ~n941;
  assign n944 = ~n946 & ~n1163;
  assign n945 = ~n946;
  assign n1164 = ~G179;
  assign n943 = ~n945 & ~n1164;
  assign n955 = n944 | n943;
  assign n1118 = ~n953 | ~n955;
  assign n1273 = ~n1118;
  assign n948 = ~G200 | ~n945;
  assign n947 = ~G190 | ~n946;
  assign n949 = ~n948 | ~n947;
  assign n950 = ~n949 & ~n953;
  assign n1191 = ~n1273 & ~n950;
  assign n952 = ~G1 & ~n951;
  assign n1276 = ~G213 | ~n952;
  assign n1749 = ~G343;
  assign n954 = ~n1542 | ~n953;
  assign n958 = ~n1191 | ~n954;
  assign n956 = ~n954;
  assign n957 = ~n956 | ~n955;
  assign n1349 = ~n958 | ~n957;
  assign n959 = ~n1349 & ~n1466;
  assign n1203 = ~n960 & ~n959;
  assign n962 = ~n1074 | ~n1736;
  assign n961 = ~G87 | ~n1120;
  assign n966 = ~n962 | ~n961;
  assign n964 = ~n1171 | ~G58;
  assign n1176 = n1175 | n1123;
  assign n963 = ~G77 | ~n1176;
  assign n965 = ~n964 | ~n963;
  assign n982 = ~n966 & ~n965;
  assign n975 = ~n982;
  assign n984 = ~n975 | ~n1542;
  assign n967 = ~n1158 | ~G238;
  assign n971 = ~n967 | ~n1133;
  assign n969 = ~n1154 | ~G232;
  assign n1131 = ~n1151;
  assign n968 = ~n1131 | ~G107;
  assign n970 = ~n969 | ~n968;
  assign n973 = ~n971 & ~n970;
  assign n972 = ~G244 | ~n1157;
  assign n978 = ~n973 | ~n972;
  assign n977 = ~n978 | ~G200;
  assign n979 = ~n978;
  assign n974 = G190 & n979;
  assign n976 = ~n975 & ~n974;
  assign n983 = n977 & n976;
  assign n981 = ~n1164 & ~n978;
  assign n980 = ~n979 & ~n1163;
  assign n985 = ~n981 & ~n980;
  assign n1117 = ~n985 & ~n982;
  assign n1192 = ~n983 & ~n1117;
  assign n987 = n984 & n1192;
  assign n986 = ~n985 & ~n984;
  assign n1411 = ~n987 & ~n986;
  assign n1265 = ~n1411;
  assign n1343 = ~G330;
  assign n1533 = ~n1542;
  assign n989 = ~G250 | ~n1154;
  assign n988 = ~G257 | ~n1158;
  assign n996 = ~n989 | ~n988;
  assign n1016 = ~G1 & ~n1458;
  assign n992 = n1296 & n1016;
  assign n1063 = ~n992 | ~G274;
  assign n991 = ~n1063;
  assign n990 = G294 & n1131;
  assign n994 = ~n991 & ~n990;
  assign n1068 = ~n1015 & ~n992;
  assign n993 = ~n1068 | ~G264;
  assign n995 = ~n994 | ~n993;
  assign n1010 = ~n996 & ~n995;
  assign n998 = ~G169 & ~n1010;
  assign n1099 = ~n1010;
  assign n997 = ~G179 & ~n1099;
  assign n1009 = ~n998 & ~n997;
  assign n1003 = ~G116 | ~n1120;
  assign n1001 = n999 | n1074;
  assign n1000 = ~G1 & ~n1691;
  assign n1077 = ~n1001 & ~n1000;
  assign n1002 = ~n1077 | ~G107;
  assign n1006 = ~n1003 | ~n1002;
  assign n1005 = ~G107 & ~n1004;
  assign n1008 = ~n1006 & ~n1005;
  assign n1007 = ~G87 | ~n1171;
  assign n1236 = ~n1008 | ~n1007;
  assign n1237 = ~n1009 | ~n1236;
  assign n1012 = ~G200 | ~n1099;
  assign n1011 = ~n1010 | ~G190;
  assign n1013 = ~n1012 | ~n1011;
  assign n1014 = n1236 | n1013;
  assign n1515 = n1237 & n1014;
  assign n1019 = ~n1016 | ~G274;
  assign n1017 = ~n1016 & ~n1015;
  assign n1018 = ~G250 | ~n1017;
  assign n1023 = ~n1019 | ~n1018;
  assign n1021 = ~G238 | ~n1154;
  assign n1020 = ~G244 | ~n1158;
  assign n1022 = ~n1021 | ~n1020;
  assign n1025 = ~n1023 & ~n1022;
  assign n1024 = ~n1131 | ~G116;
  assign n1096 = ~n1025 | ~n1024;
  assign n1027 = ~G169 | ~n1096;
  assign n1093 = ~n1096;
  assign n1026 = ~G179 | ~n1093;
  assign n1538 = ~n1027 | ~n1026;
  assign n1028 = ~n1077 | ~G87;
  assign n1029 = ~n1028 | ~n1126;
  assign n1463 = ~G107;
  assign n1653 = ~n1463 | ~n1073;
  assign n1246 = n1653 | G87;
  assign n1031 = ~n1029 | ~n1246;
  assign n1030 = ~n1120 | ~G97;
  assign n1033 = ~n1031 | ~n1030;
  assign n1032 = ~G87 & ~n1168;
  assign n1035 = ~n1033 & ~n1032;
  assign n1034 = ~n1171 | ~G68;
  assign n1535 = ~n1035 | ~n1034;
  assign n1113 = ~n1538 | ~n1535;
  assign n1037 = ~G200 | ~n1096;
  assign n1036 = ~G190 | ~n1093;
  assign n1038 = ~n1037 | ~n1036;
  assign n1039 = n1535 | n1038;
  assign n1589 = ~n1113 | ~n1039;
  assign n1040 = ~n1131 | ~G303;
  assign n1044 = ~n1063 | ~n1040;
  assign n1042 = ~n1154 | ~G257;
  assign n1041 = ~n1158 | ~G264;
  assign n1043 = ~n1042 | ~n1041;
  assign n1046 = ~n1044 & ~n1043;
  assign n1045 = ~n1068 | ~G270;
  assign n1098 = ~n1046 | ~n1045;
  assign n1054 = ~n1163 | ~n1098;
  assign n1049 = ~n1120 | ~G283;
  assign n1047 = n1077 | n1175;
  assign n1048 = ~G116 | ~n1047;
  assign n1051 = ~n1049 | ~n1048;
  assign n1050 = ~G116 & ~n1168;
  assign n1053 = ~n1051 & ~n1050;
  assign n1052 = ~n1171 | ~G97;
  assign n1240 = ~n1053 | ~n1052;
  assign n1056 = ~n1054 | ~n1240;
  assign n1055 = ~G179 & ~n1098;
  assign n1509 = ~n1056 & ~n1055;
  assign n1059 = ~G200 | ~n1098;
  assign n1057 = ~n1098;
  assign n1058 = ~G190 | ~n1057;
  assign n1060 = ~n1059 | ~n1058;
  assign n1061 = ~n1240 & ~n1060;
  assign n1241 = ~n1509 & ~n1061;
  assign n1062 = ~n1131 | ~G283;
  assign n1067 = ~n1063 | ~n1062;
  assign n1065 = ~G244 | ~n1154;
  assign n1064 = ~G250 | ~n1158;
  assign n1066 = ~n1065 | ~n1064;
  assign n1070 = ~n1067 & ~n1066;
  assign n1069 = ~n1068 | ~G257;
  assign n1097 = ~n1070 | ~n1069;
  assign n1072 = ~G179 & ~n1097;
  assign n1085 = ~n1097;
  assign n1071 = ~G169 & ~n1085;
  assign n1084 = ~n1072 & ~n1071;
  assign n1076 = ~G107 | ~n1120;
  assign n1075 = ~n1074 | ~n1073;
  assign n1081 = ~n1076 | ~n1075;
  assign n1254 = G97 ^ ~G107;
  assign n1079 = ~n1254 | ~n1175;
  assign n1078 = ~G97 | ~n1077;
  assign n1080 = ~n1079 | ~n1078;
  assign n1083 = ~n1081 & ~n1080;
  assign n1082 = ~n1171 | ~G77;
  assign n1524 = ~n1083 | ~n1082;
  assign n1110 = ~n1084 | ~n1524;
  assign n1541 = ~n1110;
  assign n1087 = ~G200 | ~n1097;
  assign n1086 = ~G190 | ~n1085;
  assign n1088 = ~n1087 | ~n1086;
  assign n1089 = ~n1524 & ~n1088;
  assign n1544 = ~n1541 & ~n1089;
  assign n1090 = ~n1241 | ~n1544;
  assign n1091 = ~n1589 & ~n1090;
  assign n1235 = ~n1515 | ~n1091;
  assign n1107 = ~n1533 | ~n1235;
  assign n1092 = ~n1098 | ~n1097;
  assign n1094 = ~n1093 & ~n1092;
  assign n1095 = ~n1094 | ~n1099;
  assign n1104 = ~n1095 | ~n1164;
  assign n1101 = ~n1097 & ~n1096;
  assign n1100 = ~n1099 & ~n1098;
  assign n1102 = ~n1101 | ~n1100;
  assign n1103 = ~G179 | ~n1102;
  assign n1105 = ~n1104 | ~n1103;
  assign n1106 = ~n1542 | ~n1105;
  assign n1269 = ~n1107 | ~n1106;
  assign n1251 = ~n1343 & ~n1269;
  assign n1350 = n1265 & n1251;
  assign n1111 = ~n1589;
  assign n1108 = ~n1515 | ~n1509;
  assign n1245 = ~n1237 | ~n1108;
  assign n1109 = ~n1544 | ~n1245;
  assign n1532 = ~n1110 | ~n1109;
  assign n1112 = ~n1111 | ~n1532;
  assign n1739 = ~n1113 | ~n1112;
  assign n1195 = ~n1533 | ~n1739;
  assign n1250 = ~n1195;
  assign n1115 = ~n1250 | ~n1192;
  assign n1114 = ~n1117 | ~n1533;
  assign n1272 = ~n1115 | ~n1114;
  assign n1116 = ~n1350 & ~n1272;
  assign n1361 = n1116 ^ ~n1349;
  assign n1119 = ~n1191 | ~n1117;
  assign n1148 = ~n1119 | ~n1118;
  assign n1167 = ~n1120;
  assign n1453 = ~G68;
  assign n1122 = ~n1167 & ~n1453;
  assign n1121 = ~G58 & ~n1168;
  assign n1130 = ~n1122 & ~n1121;
  assign n1125 = ~G58 | ~n1123;
  assign n1124 = ~G159 | ~n1171;
  assign n1128 = ~n1125 | ~n1124;
  assign n1231 = G68 ^ G58;
  assign n1127 = ~n1231 & ~n1126;
  assign n1129 = ~n1128 & ~n1127;
  assign n1258 = ~n1130 | ~n1129;
  assign n1132 = ~n1131 | ~G87;
  assign n1137 = ~n1133 | ~n1132;
  assign n1135 = ~G223 | ~n1154;
  assign n1134 = ~G226 | ~n1158;
  assign n1136 = ~n1135 | ~n1134;
  assign n1139 = ~n1137 & ~n1136;
  assign n1138 = ~n1157 | ~G232;
  assign n1142 = ~n1139 | ~n1138;
  assign n1141 = ~G169 | ~n1142;
  assign n1143 = ~n1142;
  assign n1140 = ~G179 | ~n1143;
  assign n1261 = ~n1141 | ~n1140;
  assign n1149 = ~n1258 | ~n1261;
  assign n1277 = ~n1149;
  assign n1145 = ~G200 | ~n1142;
  assign n1144 = ~G190 | ~n1143;
  assign n1146 = ~n1145 | ~n1144;
  assign n1147 = ~n1146 & ~n1258;
  assign n1259 = ~n1277 & ~n1147;
  assign n1150 = ~n1148 | ~n1259;
  assign n1188 = ~n1150 | ~n1149;
  assign n1152 = ~n1151 & ~n1736;
  assign n1156 = ~n1153 & ~n1152;
  assign n1155 = ~n1154 | ~G222;
  assign n1162 = ~n1156 | ~n1155;
  assign n1160 = ~G226 | ~n1157;
  assign n1159 = ~G223 | ~n1158;
  assign n1161 = ~n1160 | ~n1159;
  assign n1183 = ~n1162 & ~n1161;
  assign n1166 = ~n1183 & ~n1163;
  assign n1182 = ~n1183;
  assign n1165 = ~n1182 & ~n1164;
  assign n1337 = ~n1166 & ~n1165;
  assign n1174 = ~G58;
  assign n1170 = ~n1167 & ~n1174;
  assign n1169 = ~G50 & ~n1168;
  assign n1173 = ~n1170 & ~n1169;
  assign n1172 = ~n1171 | ~G150;
  assign n1180 = ~n1173 | ~n1172;
  assign n1738 = ~n1453 | ~n1174;
  assign n1178 = ~n1175 | ~n1738;
  assign n1177 = ~G50 | ~n1176;
  assign n1179 = ~n1178 | ~n1177;
  assign n1181 = ~n1180 & ~n1179;
  assign n1189 = ~n1337 & ~n1181;
  assign n1334 = ~n1181;
  assign n1185 = ~G200 | ~n1182;
  assign n1184 = ~G190 | ~n1183;
  assign n1186 = ~n1185 | ~n1184;
  assign n1187 = ~n1334 & ~n1186;
  assign n1335 = ~n1189 & ~n1187;
  assign n1190 = n1188 & n1335;
  assign n1742 = ~n1190 & ~n1189;
  assign n1197 = ~n1742;
  assign n1194 = n1259 & n1335;
  assign n1193 = n1192 & n1191;
  assign n1268 = ~n1194 | ~n1193;
  assign n1196 = ~n1268 & ~n1195;
  assign n1282 = ~n1197 & ~n1196;
  assign n1740 = ~n1268;
  assign n1198 = ~n1251 | ~n1740;
  assign n1404 = ~n1282 | ~n1198;
  assign n1199 = n1361 ^ ~n1404;
  assign n1201 = ~n1199 | ~n1643;
  assign n1200 = ~n1361 | ~n1530;
  assign n1202 = ~n1201 | ~n1200;
  assign G381 = n1203 | n1202;
  assign n1664 = ~G50 | ~n1738;
  assign n1228 = G226 ^ G232;
  assign n1227 = G244 ^ ~G238;
  assign n1459 = n1228 ^ ~n1227;
  assign n1229 = G257 ^ ~G250;
  assign n1230 = n1229 ^ ~G270;
  assign n1552 = G264 ^ ~n1230;
  assign n1232 = G50 ^ ~n1231;
  assign n1661 = n1232 ^ ~n1736;
  assign n1233 = G87 ^ ~G116;
  assign n1234 = n1233 ^ ~G97;
  assign n1634 = G107 ^ ~n1234;
  assign n1510 = ~n1236 | ~n1542;
  assign n1239 = n1510 & n1515;
  assign n1238 = ~n1237 & ~n1533;
  assign n1505 = ~n1239 & ~n1238;
  assign n1242 = ~n1240 | ~n1542;
  assign n1244 = ~n1242 | ~n1241;
  assign n1243 = ~n1509 | ~n1542;
  assign n1716 = ~n1244 | ~n1243;
  assign n1512 = ~G330 | ~n1716;
  assign n1547 = ~n1505 & ~n1512;
  assign n1527 = ~n1547;
  assign n1525 = ~n1533 | ~n1245;
  assign n1519 = ~n1643;
  assign n1467 = ~G116 & ~n1246;
  assign n1640 = ~n1251 & ~n1250;
  assign n1656 = ~G116;
  assign n1333 = ~n1276;
  assign n1260 = ~n1333 | ~n1258;
  assign n1264 = ~n1259 | ~n1260;
  assign n1262 = ~n1260;
  assign n1263 = ~n1262 | ~n1261;
  assign n1396 = ~n1264 | ~n1263;
  assign n1266 = ~n1265 | ~n1396;
  assign n1267 = ~n1269 & ~n1266;
  assign n1342 = ~n1267 | ~n1349;
  assign n1275 = ~n1272 | ~n1349;
  assign n1274 = ~n1273 | ~n1533;
  assign n1348 = ~n1275 | ~n1274;
  assign n1279 = ~n1348 | ~n1396;
  assign n1278 = ~n1277 | ~n1276;
  assign n1345 = ~n1279 | ~n1278;
  assign n1443 = ~n1713;
  assign n1330 = ~n1443 | ~n1296;
  assign n1658 = ~n1466;
  assign n1297 = ~n1658 & ~G50;
  assign n1298 = ~n1330 | ~n1297;
  assign n1332 = ~n1655 | ~n1298;
  assign n1300 = ~n1704 | ~G116;
  assign n1299 = ~n1692 | ~G87;
  assign n1304 = ~n1300 | ~n1299;
  assign n1302 = ~n1697 | ~G283;
  assign n1301 = ~n1696 | ~G97;
  assign n1303 = ~n1302 | ~n1301;
  assign n1310 = ~n1304 & ~n1303;
  assign n1562 = ~G68 | ~n1693;
  assign n1305 = ~G107 | ~n1686;
  assign n1308 = ~n1562 | ~n1305;
  assign n1472 = ~G77 | ~n1705;
  assign n1307 = ~n1306 | ~n1472;
  assign n1309 = ~n1308 & ~n1307;
  assign n1311 = ~n1310 | ~n1309;
  assign n1328 = ~G33 | ~n1311;
  assign n1313 = ~G124 | ~n1697;
  assign n1312 = ~G137 | ~n1692;
  assign n1317 = ~n1313 | ~n1312;
  assign n1315 = ~G132 | ~n1696;
  assign n1314 = ~n1687 | ~G159;
  assign n1316 = ~n1315 | ~n1314;
  assign n1325 = ~n1317 & ~n1316;
  assign n1319 = ~G143 | ~n1705;
  assign n1318 = ~n1693 | ~G150;
  assign n1323 = ~n1319 | ~n1318;
  assign n1321 = ~G125 | ~n1704;
  assign n1320 = ~G128 | ~n1686;
  assign n1322 = ~n1321 | ~n1320;
  assign n1324 = ~n1323 & ~n1322;
  assign n1326 = ~n1325 | ~n1324;
  assign n1327 = ~n1691 | ~n1326;
  assign n1329 = ~n1328 | ~n1327;
  assign n1331 = ~n1330 & ~n1329;
  assign n1341 = ~n1332 & ~n1331;
  assign n1336 = ~n1334 | ~n1333;
  assign n1339 = n1336 & n1335;
  assign n1338 = ~n1337 & ~n1336;
  assign n1346 = ~n1339 & ~n1338;
  assign n1340 = ~n1658 | ~n1346;
  assign n1360 = ~n1341 | ~n1340;
  assign n1344 = ~n1343 & ~n1342;
  assign n1347 = ~n1345 & ~n1344;
  assign n1357 = n1347 ^ ~n1346;
  assign n1521 = ~n1530;
  assign n1352 = ~n1348;
  assign n1351 = ~n1350 | ~n1349;
  assign n1353 = ~n1352 | ~n1351;
  assign n1406 = n1396 ^ n1353;
  assign n1354 = ~n1361 | ~n1406;
  assign n1355 = ~n1521 | ~n1354;
  assign n1356 = ~n1404 & ~n1355;
  assign n1358 = ~n1357 & ~n1356;
  assign n1721 = ~n1655;
  assign n1359 = ~n1358 | ~n1721;
  assign G375 = ~n1360 | ~n1359;
  assign n1363 = n1361 ^ n1406;
  assign n1362 = ~n1404;
  assign n1364 = ~n1363 | ~n1362;
  assign n1403 = ~n1519 & ~n1364;
  assign n1366 = ~G128 | ~n1704;
  assign n1365 = ~n1705 | ~G150;
  assign n1379 = ~n1366 | ~n1365;
  assign n1368 = ~G132 | ~n1686;
  assign n1367 = ~n1687 | ~G50;
  assign n1369 = ~n1368 | ~n1367;
  assign n1377 = ~G33 & ~n1369;
  assign n1371 = ~G143 | ~n1692;
  assign n1370 = ~n1693 | ~G159;
  assign n1375 = ~n1371 | ~n1370;
  assign n1373 = ~G137 | ~n1696;
  assign n1372 = ~G125 | ~n1697;
  assign n1374 = ~n1373 | ~n1372;
  assign n1376 = ~n1375 & ~n1374;
  assign n1378 = ~n1377 | ~n1376;
  assign n1394 = ~n1379 & ~n1378;
  assign n1414 = ~n1453 & ~n1380;
  assign n1673 = ~G87 | ~n1705;
  assign n1382 = ~n1704 | ~G283;
  assign n1381 = ~n1686 | ~G116;
  assign n1390 = ~n1382 | ~n1381;
  assign n1384 = G97 & n1692;
  assign n1383 = G294 & n1697;
  assign n1388 = ~n1384 & ~n1383;
  assign n1604 = G77 & n1693;
  assign n1385 = ~G107 | ~n1696;
  assign n1386 = ~G33 | ~n1385;
  assign n1387 = ~n1604 & ~n1386;
  assign n1389 = ~n1388 | ~n1387;
  assign n1391 = ~n1390 & ~n1389;
  assign n1392 = ~n1673 | ~n1391;
  assign n1393 = ~n1414 & ~n1392;
  assign n1395 = ~n1394 & ~n1393;
  assign n1398 = ~n1395 & ~n1713;
  assign n1397 = ~n1396 & ~n1466;
  assign n1399 = ~n1398 & ~n1397;
  assign n1401 = ~n1655 | ~n1399;
  assign n1400 = ~n1446 & ~G58;
  assign n1402 = ~n1401 & ~n1400;
  assign n1409 = ~n1403 & ~n1402;
  assign n1405 = ~n1404 | ~n1643;
  assign n1407 = ~n1405 | ~n1521;
  assign n1408 = ~n1407 | ~n1406;
  assign G378 = ~n1409 | ~n1408;
  assign n1410 = n1411 ^ n1640;
  assign n1451 = ~n1655 & ~n1410;
  assign n1445 = ~n1411 | ~n1658;
  assign n1413 = ~G132 | ~n1697;
  assign n1412 = ~n1696 | ~G150;
  assign n1418 = ~n1413 | ~n1412;
  assign n1416 = ~G33 & ~n1414;
  assign n1415 = ~n1686 | ~G143;
  assign n1417 = ~n1416 | ~n1415;
  assign n1426 = ~n1418 & ~n1417;
  assign n1420 = ~G137 | ~n1704;
  assign n1419 = ~n1705 | ~G50;
  assign n1424 = ~n1420 | ~n1419;
  assign n1422 = ~n1692 | ~G159;
  assign n1421 = ~n1693 | ~G58;
  assign n1423 = ~n1422 | ~n1421;
  assign n1425 = ~n1424 & ~n1423;
  assign n1441 = ~n1426 | ~n1425;
  assign n1428 = ~G311 | ~n1697;
  assign n1427 = ~n1692 | ~G116;
  assign n1432 = ~n1428 | ~n1427;
  assign n1601 = G87 & n1687;
  assign n1430 = ~n1601 & ~n1691;
  assign n1429 = ~G283 | ~n1696;
  assign n1431 = ~n1430 | ~n1429;
  assign n1439 = ~n1432 & ~n1431;
  assign n1677 = ~G97 | ~n1693;
  assign n1433 = ~G294 | ~n1686;
  assign n1437 = ~n1677 | ~n1433;
  assign n1435 = ~n1704 | ~G303;
  assign n1434 = ~n1705 | ~G107;
  assign n1436 = ~n1435 | ~n1434;
  assign n1438 = ~n1437 & ~n1436;
  assign n1440 = ~n1439 | ~n1438;
  assign n1442 = ~n1441 | ~n1440;
  assign n1444 = ~n1443 | ~n1442;
  assign n1448 = ~n1445 | ~n1444;
  assign n1447 = ~G77 & ~n1446;
  assign n1449 = ~n1448 & ~n1447;
  assign n1450 = ~n1721 & ~n1449;
  assign G384 = ~n1451 & ~n1450;
  assign n1717 = ~n1658 | ~n1452;
  assign n1669 = ~n1713 | ~n1717;
  assign n1735 = ~G50;
  assign n1455 = ~n1467 | ~n1735;
  assign n1454 = ~n1736 & ~n1453;
  assign n1456 = ~n1455 & ~n1454;
  assign n1457 = ~n1456 | ~G58;
  assign n1461 = ~n1458 | ~n1457;
  assign n1460 = ~G45 | ~n1459;
  assign n1462 = ~n1461 | ~n1460;
  assign n1663 = ~n1657 & ~n1691;
  assign n1465 = ~n1462 | ~n1663;
  assign n1464 = ~n1463 | ~n1657;
  assign n1469 = ~n1465 | ~n1464;
  assign n1468 = ~n1467 & ~n1466;
  assign n1470 = ~n1469 & ~n1468;
  assign n1504 = ~n1669 & ~n1470;
  assign n1581 = ~G97 | ~n1687;
  assign n1471 = ~G50 | ~n1686;
  assign n1484 = ~n1581 | ~n1471;
  assign n1474 = ~n1473 | ~n1472;
  assign n1482 = ~G33 & ~n1474;
  assign n1476 = ~n1704 | ~G159;
  assign n1475 = ~n1692 | ~G68;
  assign n1480 = ~n1476 | ~n1475;
  assign n1478 = ~n1697 | ~G150;
  assign n1477 = ~n1696 | ~G58;
  assign n1479 = ~n1478 | ~n1477;
  assign n1481 = ~n1480 & ~n1479;
  assign n1483 = ~n1482 | ~n1481;
  assign n1501 = ~n1484 & ~n1483;
  assign n1486 = ~G317 | ~n1686;
  assign n1485 = ~n1687 | ~G116;
  assign n1487 = ~n1486 | ~n1485;
  assign n1495 = ~n1691 & ~n1487;
  assign n1489 = ~n1693 | ~G283;
  assign n1488 = ~n1692 | ~G303;
  assign n1493 = ~n1489 | ~n1488;
  assign n1491 = ~G311 | ~n1696;
  assign n1490 = ~G326 | ~n1697;
  assign n1492 = ~n1491 | ~n1490;
  assign n1494 = ~n1493 & ~n1492;
  assign n1499 = ~n1495 | ~n1494;
  assign n1497 = ~G322 | ~n1704;
  assign n1496 = ~n1705 | ~G294;
  assign n1498 = ~n1497 | ~n1496;
  assign n1500 = ~n1499 & ~n1498;
  assign n1502 = ~n1501 & ~n1500;
  assign n1503 = ~n1713 & ~n1502;
  assign n1507 = ~n1504 & ~n1503;
  assign n1590 = ~n1717;
  assign n1506 = ~n1505 | ~n1590;
  assign n1508 = ~n1507 | ~n1506;
  assign n1518 = ~n1721 & ~n1508;
  assign n1511 = ~n1509 | ~n1533;
  assign n1513 = ~n1511 | ~n1510;
  assign n1514 = n1513 ^ ~n1512;
  assign n1641 = n1515 ^ n1514;
  assign n1516 = ~n1640 | ~n1643;
  assign n1517 = ~n1641 & ~n1516;
  assign n1523 = ~n1518 & ~n1517;
  assign n1520 = n1519 | n1640;
  assign n1649 = ~n1521 | ~n1520;
  assign n1522 = ~n1641 | ~n1649;
  assign G393 = ~n1523 | ~n1522;
  assign n1543 = ~n1542 | ~n1524;
  assign n1526 = ~n1525 | ~n1543;
  assign n1528 = n1527 ^ n1526;
  assign n1650 = n1544 ^ ~n1528;
  assign n1644 = ~n1650 | ~n1641;
  assign n1529 = ~n1640 | ~n1644;
  assign n1531 = ~n1530 & ~n1529;
  assign n1551 = ~n1655 & ~n1531;
  assign n1534 = ~n1533 | ~n1532;
  assign n1536 = n1534 ^ ~n1589;
  assign n1537 = ~n1542 | ~n1535;
  assign n1540 = ~n1536 | ~n1537;
  assign n1539 = n1538 | n1537;
  assign n1549 = ~n1540 | ~n1539;
  assign n1546 = ~n1542 | ~n1541;
  assign n1545 = ~n1544 | ~n1543;
  assign n1630 = ~n1546 | ~n1545;
  assign n1548 = ~n1547 | ~n1630;
  assign n1550 = n1549 ^ n1548;
  assign n1597 = ~n1551 | ~n1550;
  assign n1554 = ~n1663 | ~n1552;
  assign n1553 = ~G87 | ~n1657;
  assign n1555 = ~n1554 | ~n1553;
  assign n1594 = ~n1555 & ~n1669;
  assign n1557 = ~G143 | ~n1704;
  assign n1556 = ~n1705 | ~G58;
  assign n1569 = ~n1557 | ~n1556;
  assign n1558 = n1686 & G150;
  assign n1567 = ~n1559 & ~n1558;
  assign n1561 = ~G137 | ~n1697;
  assign n1560 = ~n1692 | ~G50;
  assign n1565 = ~n1561 | ~n1560;
  assign n1563 = ~G159 | ~n1696;
  assign n1564 = ~n1563 | ~n1562;
  assign n1566 = ~n1565 & ~n1564;
  assign n1568 = ~n1567 | ~n1566;
  assign n1570 = ~n1569 & ~n1568;
  assign n1571 = ~G33 & ~n1570;
  assign n1588 = ~n1713 & ~n1571;
  assign n1573 = ~n1692 | ~G283;
  assign n1572 = ~n1693 | ~G107;
  assign n1577 = ~n1573 | ~n1572;
  assign n1575 = ~G317 | ~n1697;
  assign n1574 = ~n1696 | ~G294;
  assign n1576 = ~n1575 | ~n1574;
  assign n1585 = ~n1577 & ~n1576;
  assign n1579 = ~G311 | ~n1704;
  assign n1578 = ~n1705 | ~G116;
  assign n1583 = ~n1579 | ~n1578;
  assign n1580 = ~G303 | ~n1686;
  assign n1582 = ~n1581 | ~n1580;
  assign n1584 = ~n1583 & ~n1582;
  assign n1586 = ~n1585 | ~n1584;
  assign n1587 = ~G33 | ~n1586;
  assign n1592 = ~n1588 | ~n1587;
  assign n1591 = ~n1590 | ~n1589;
  assign n1593 = ~n1592 | ~n1591;
  assign n1595 = ~n1594 & ~n1593;
  assign n1596 = ~n1595 | ~n1655;
  assign G387 = ~n1597 | ~n1596;
  assign n1599 = ~n1704 | ~G150;
  assign n1598 = ~n1705 | ~G68;
  assign n1612 = ~n1599 | ~n1598;
  assign n1600 = n1696 & G50;
  assign n1610 = ~n1601 & ~n1600;
  assign n1603 = ~G143 | ~n1697;
  assign n1602 = ~n1692 | ~G58;
  assign n1608 = ~n1603 | ~n1602;
  assign n1606 = ~G33 & ~n1604;
  assign n1605 = ~G159 | ~n1686;
  assign n1607 = ~n1606 | ~n1605;
  assign n1609 = ~n1608 & ~n1607;
  assign n1611 = ~n1610 | ~n1609;
  assign n1628 = ~n1612 & ~n1611;
  assign n1674 = ~G107 | ~n1687;
  assign n1613 = ~n1686 | ~G311;
  assign n1614 = ~n1674 | ~n1613;
  assign n1622 = ~n1691 & ~n1614;
  assign n1616 = ~n1693 | ~G116;
  assign n1615 = ~n1692 | ~G294;
  assign n1620 = ~n1616 | ~n1615;
  assign n1618 = ~G322 | ~n1697;
  assign n1617 = ~n1696 | ~G303;
  assign n1619 = ~n1618 | ~n1617;
  assign n1621 = ~n1620 & ~n1619;
  assign n1626 = ~n1622 | ~n1621;
  assign n1624 = ~G317 | ~n1704;
  assign n1623 = ~n1705 | ~G283;
  assign n1625 = ~n1624 | ~n1623;
  assign n1627 = ~n1626 & ~n1625;
  assign n1629 = ~n1628 & ~n1627;
  assign n1632 = ~n1713 & ~n1629;
  assign n1631 = ~n1717 & ~n1630;
  assign n1633 = ~n1632 & ~n1631;
  assign n1639 = ~n1655 | ~n1633;
  assign n1636 = ~n1663 | ~n1634;
  assign n1635 = ~G97 | ~n1657;
  assign n1637 = ~n1636 | ~n1635;
  assign n1638 = ~n1669 & ~n1637;
  assign n1648 = ~n1639 & ~n1638;
  assign n1642 = n1641 & n1640;
  assign n1646 = ~n1650 & ~n1642;
  assign n1645 = ~n1644 | ~n1643;
  assign n1647 = ~n1646 & ~n1645;
  assign n1652 = ~n1648 & ~n1647;
  assign n1651 = ~n1650 | ~n1649;
  assign G390 = ~n1652 | ~n1651;
  assign G355 = ~G87 | ~n1653;
  assign n1654 = G330 ^ n1716;
  assign n1723 = ~n1655 & ~n1654;
  assign n1660 = ~n1657 | ~n1656;
  assign n1659 = ~n1658 | ~G355;
  assign n1668 = ~n1660 | ~n1659;
  assign n1662 = ~G45 | ~n1661;
  assign n1666 = ~n1663 | ~n1662;
  assign n1665 = ~G45 & ~n1664;
  assign n1667 = ~n1666 & ~n1665;
  assign n1670 = ~n1668 & ~n1667;
  assign n1715 = ~n1670 & ~n1669;
  assign n1672 = ~n1704 | ~G50;
  assign n1671 = ~n1686 | ~G58;
  assign n1685 = ~n1672 | ~n1671;
  assign n1675 = ~n1674 | ~n1673;
  assign n1683 = ~G33 & ~n1675;
  assign n1676 = ~G77 | ~n1692;
  assign n1681 = ~n1677 | ~n1676;
  assign n1679 = ~n1697 | ~G159;
  assign n1678 = ~n1696 | ~G68;
  assign n1680 = ~n1679 | ~n1678;
  assign n1682 = ~n1681 & ~n1680;
  assign n1684 = ~n1683 | ~n1682;
  assign n1711 = ~n1685 & ~n1684;
  assign n1689 = ~G322 | ~n1686;
  assign n1688 = ~n1687 | ~G283;
  assign n1690 = ~n1689 | ~n1688;
  assign n1703 = ~n1691 & ~n1690;
  assign n1695 = ~G311 | ~n1692;
  assign n1694 = ~n1693 | ~G294;
  assign n1701 = ~n1695 | ~n1694;
  assign n1699 = ~G317 | ~n1696;
  assign n1698 = ~G329 | ~n1697;
  assign n1700 = ~n1699 | ~n1698;
  assign n1702 = ~n1701 & ~n1700;
  assign n1709 = ~n1703 | ~n1702;
  assign n1707 = ~G326 | ~n1704;
  assign n1706 = ~n1705 | ~G303;
  assign n1708 = ~n1707 | ~n1706;
  assign n1710 = ~n1709 & ~n1708;
  assign n1712 = ~n1711 & ~n1710;
  assign n1714 = ~n1713 & ~n1712;
  assign n1719 = n1715 | n1714;
  assign n1718 = ~n1717 & ~n1716;
  assign n1720 = ~n1719 & ~n1718;
  assign n1722 = ~n1721 & ~n1720;
  assign G396 = ~n1723 & ~n1722;
  assign n1724 = ~G213 | ~n1749;
  assign n1733 = G375 ^ G378;
  assign n1727 = ~n1724 | ~n1733;
  assign n1725 = ~n1724;
  assign n1726 = ~n1725 | ~G2897;
  assign n1732 = ~n1727 | ~n1726;
  assign n1728 = G387 ^ G390;
  assign n1729 = G393 ^ ~n1728;
  assign n1731 = G384 ^ ~n1729;
  assign n1730 = G381 ^ ~G396;
  assign n1734 = n1731 ^ ~n1730;
  assign G405_Lock = n1732 ^ ~n1734;
  assign keyinput_0 = 1'b0;
  assign keyinput_1 = 1'b1;
  assign keyinput_2 = 1'b1;
  assign keyinput_3 = 1'b1;
  assign keyinput_4 = 1'b0;
  assign keyinput_5 = 1'b0;
  assign keyinput_6 = 1'b0;
  assign keyinput_7 = 1'b0;
  assign keyinput_8 = 1'b1;
  assign keyinput_9 = 1'b1;
  assign keyinput_10 = 1'b1;
  assign keyinput_11 = 1'b0;
  assign keyinput_12 = 1'b1;
  assign keyinput_13 = 1'b1;
  assign keyinput_14 = 1'b0;
  assign keyinput_15 = 1'b1;
  assign keyinput_16 = 1'b1;
  assign keyinput_17 = 1'b1;
  assign keyinput_18 = 1'b0;
  assign keyinput_19 = 1'b1;
  assign keyinput_20 = 1'b0;
  assign keyinput_21 = 1'b0;
  assign keyinput_22 = 1'b0;
  assign keyinput_23 = 1'b1;
  assign keyinput_24 = 1'b0;
  assign keyinput_25 = 1'b0;
  assign keyinput_26 = 1'b1;
  assign keyinput_27 = 1'b0;
  assign keyinput_28 = 1'b1;
  assign keyinput_29 = 1'b0;
  assign keyinput_30 = 1'b0;
  assign keyinput_31 = 1'b0;
  assign keyinput_32 = 1'b0;
  assign keyinput_33 = 1'b1;
  assign keyinput_34 = 1'b0;
  assign keyinput_35 = 1'b1;
  assign keyinput_36 = 1'b0;
  assign keyinput_37 = 1'b1;
  assign keyinput_38 = 1'b0;
  assign keyinput_39 = 1'b0;
  assign keyinput_40 = 1'b1;
  assign keyinput_41 = 1'b0;
  assign keyinput_42 = 1'b0;
  assign keyinput_43 = 1'b0;
  assign keyinput_44 = 1'b1;
  assign keyinput_45 = 1'b1;
  assign keyinput_46 = 1'b1;
  assign keyinput_47 = 1'b1;
  assign keyinput_48 = 1'b0;
  assign keyinput_49 = 1'b0;
  assign keyinput_50 = 1'b0;
  assign keyinput_51 = 1'b1;
  assign keyinput_52 = 1'b1;
  assign keyinput_53 = 1'b1;
  assign keyinput_54 = 1'b1;
  assign keyinput_55 = 1'b0;
  assign keyinput_56 = 1'b1;
  assign keyinput_57 = 1'b0;
  assign keyinput_58 = 1'b0;
  assign keyinput_59 = 1'b1;
  assign keyinput_60 = 1'b1;
  assign keyinput_61 = 1'b1;
  assign keyinput_62 = 1'b0;
  assign keyinput_63 = 1'b0;
  assign input_0 = keyinput_0 ^ G1;
  assign input_1 = keyinput_1 ^ G13;
  assign AND_1 = input_0 & input_1;
  assign input_2 = keyinput_2 ^ G20;
  assign OR_2 = input_2 | AND_1;
  assign input_3 = keyinput_3 ^ G33;
  assign AND_3 = input_3 & OR_2;
  assign input_4 = keyinput_4 ^ G41;
  assign OR_4 = input_4 | AND_3;
  assign input_5 = keyinput_5 ^ G45;
  assign OR_5 = input_5 | OR_4;
  assign input_6 = keyinput_6 ^ G50;
  assign OR_6 = input_6 | OR_5;
  assign input_7 = keyinput_7 ^ G58;
  assign AND_7 = input_7 & OR_6;
  assign input_8 = keyinput_8 ^ G68;
  assign OR_8 = input_8 | AND_7;
  assign input_9 = keyinput_9 ^ G77;
  assign OR_9 = input_9 | OR_8;
  assign input_10 = keyinput_10 ^ G87;
  assign AND_10 = input_10 & OR_9;
  assign input_11 = keyinput_11 ^ G97;
  assign AND_11 = input_11 & AND_10;
  assign input_12 = keyinput_12 ^ G107;
  assign AND_12 = input_12 & AND_11;
  assign input_13 = keyinput_13 ^ G116;
  assign OR_13 = input_13 | AND_12;
  assign input_14 = keyinput_14 ^ G124;
  assign OR_14 = input_14 | OR_13;
  assign input_15 = keyinput_15 ^ G125;
  assign AND_15 = input_15 & OR_14;
  assign input_16 = keyinput_16 ^ G128;
  assign AND_16 = input_16 & AND_15;
  assign input_17 = keyinput_17 ^ G132;
  assign OR_17 = input_17 | AND_16;
  assign input_18 = keyinput_18 ^ G137;
  assign OR_18 = input_18 | OR_17;
  assign input_19 = keyinput_19 ^ G143;
  assign OR_19 = input_19 | OR_18;
  assign input_20 = keyinput_20 ^ G150;
  assign OR_20 = input_20 | OR_19;
  assign input_21 = keyinput_21 ^ G159;
  assign AND_21 = input_21 & OR_20;
  assign input_22 = keyinput_22 ^ G169;
  assign AND_22 = input_22 & AND_21;
  assign input_23 = keyinput_23 ^ G179;
  assign OR_23 = input_23 | AND_22;
  assign input_24 = keyinput_24 ^ G190;
  assign OR_24 = input_24 | OR_23;
  assign input_25 = keyinput_25 ^ G200;
  assign AND_25 = input_25 & OR_24;
  assign input_26 = keyinput_26 ^ G213;
  assign OR_26 = input_26 | AND_25;
  assign input_27 = keyinput_27 ^ G222;
  assign AND_27 = input_27 & OR_26;
  assign input_28 = keyinput_28 ^ G223;
  assign AND_28 = input_28 & AND_27;
  assign input_29 = keyinput_29 ^ G226;
  assign OR_29 = input_29 | AND_28;
  assign input_30 = keyinput_30 ^ G232;
  assign AND_30 = input_30 & OR_29;
  assign input_31 = keyinput_31 ^ G238;
  assign OR_31 = input_31 | AND_30;
  assign input_32 = keyinput_32 ^ G1;
  assign input_33 = keyinput_33 ^ G13;
  assign AND_33 = input_32 & input_33;
  assign input_34 = keyinput_34 ^ G20;
  assign OR_34 = input_34 | AND_33;
  assign input_35 = keyinput_35 ^ G33;
  assign AND_35 = input_35 & OR_34;
  assign input_36 = keyinput_36 ^ G41;
  assign OR_36 = input_36 | AND_35;
  assign input_37 = keyinput_37 ^ G45;
  assign OR_37 = input_37 | OR_36;
  assign input_38 = keyinput_38 ^ G50;
  assign OR_38 = input_38 | OR_37;
  assign input_39 = keyinput_39 ^ G58;
  assign AND_39 = input_39 & OR_38;
  assign input_40 = keyinput_40 ^ G68;
  assign OR_40 = input_40 | AND_39;
  assign input_41 = keyinput_41 ^ G77;
  assign OR_41 = input_41 | OR_40;
  assign input_42 = keyinput_42 ^ G87;
  assign AND_42 = input_42 & OR_41;
  assign input_43 = keyinput_43 ^ G97;
  assign AND_43 = input_43 & AND_42;
  assign input_44 = keyinput_44 ^ G107;
  assign AND_44 = input_44 & AND_43;
  assign input_45 = keyinput_45 ^ G116;
  assign OR_45 = input_45 | AND_44;
  assign input_46 = keyinput_46 ^ G124;
  assign OR_46 = input_46 | OR_45;
  assign input_47 = keyinput_47 ^ G125;
  assign AND_47 = input_47 & OR_46;
  assign input_48 = keyinput_48 ^ G128;
  assign AND_48 = input_48 & AND_47;
  assign input_49 = keyinput_49 ^ G132;
  assign OR_49 = input_49 | AND_48;
  assign input_50 = keyinput_50 ^ G137;
  assign OR_50 = input_50 | OR_49;
  assign input_51 = keyinput_51 ^ G143;
  assign OR_51 = input_51 | OR_50;
  assign input_52 = keyinput_52 ^ G150;
  assign OR_52 = input_52 | OR_51;
  assign input_53 = keyinput_53 ^ G159;
  assign AND_53 = input_53 & OR_52;
  assign input_54 = keyinput_54 ^ G169;
  assign AND_54 = input_54 & AND_53;
  assign input_55 = keyinput_55 ^ G179;
  assign OR_55 = input_55 | AND_54;
  assign input_56 = keyinput_56 ^ G190;
  assign OR_56 = input_56 | OR_55;
  assign input_57 = keyinput_57 ^ G200;
  assign AND_57 = input_57 & OR_56;
  assign input_58 = keyinput_58 ^ G213;
  assign OR_58 = input_58 | AND_57;
  assign input_59 = keyinput_59 ^ G222;
  assign AND_59 = input_59 & OR_58;
  assign input_60 = keyinput_60 ^ G223;
  assign AND_60 = input_60 & AND_59;
  assign input_61 = keyinput_61 ^ G226;
  assign OR_61 = input_61 | AND_60;
  assign input_62 = keyinput_62 ^ G232;
  assign AND_62 = input_62 & OR_61;
  assign input_63 = keyinput_63 ^ G238;
  assign OR_63 = input_63 | AND_62;
  assign OR_63_INV = ~OR_63;
  assign CASOP = OR_31 & OR_63_INV;
  assign G405 = G405_Lock ^ CASOP;
endmodule


