// Benchmark "c7552" written by ABC on Thu Mar  5 01:07:52 2020

module c7552 ( 
    G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
    G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
    G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
    G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
    G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134,
    G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156,
    G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496,
    G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253,
    G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743,
    G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432,
    G4437, G4526, G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41,
    G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63,
    G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81,
    G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106,
    G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130,
    G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166,
    G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190,
    G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202,
    G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214,
    G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226,
    G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238,
    G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486,
    G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239,
    G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729,
    G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420,
    G4427, G4432, G4437, G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire G400, G1184, G1501, G2857, G4442, G4514, G401, G573, G574, G575,
    G1178, G1186, G1192, G1198, G1205, G1206, G1207, G1210, G1458, G1461,
    G1464, G1471, G1475, G1482, G1488, G1495, G1499, G1500, G1503, G1512,
    G1518, G1524, G1535, G1541, G2207, G2210, G2213, G2220, G2226, G2232,
    G2238, G2241, G2249, G2255, G2258, G2828, G3700, G3703, G3707, G3713,
    G3719, G3725, G3731, G3739, G3745, G3751, G4121, G4396, G4402, G4407,
    G4412, G4417, G4422, G4429, G4434, G4439, G4833, G2876, G2878, G1519,
    G2871, G2883, G280, G4839, G572, G581, G587, G601, G606, G650, G657,
    G671, G678, G777, G1115, G1336, G1350, G1477, G1507, G1514, G1530,
    G2259, G2833, G2872, G2886, G2892, G2905, G2909, G3622, G3635, G3755,
    G4640, G4653, G4873, G4876, G4881, G4889, G4905, G4916, G4921, G5175,
    G5178, G5186, G5191, G5199, G5215, G5223, G5393, G5401, G5409, G5417,
    G5425, G5433, G5441, G5449, G5457, G5745, G5753, G5761, G5769, G5777,
    G5785, G5793, G5801, G5809, G5865, G5873, G5881, G5889, G5897, G5905,
    G5913, G5921, G5985, G5993, G6001, G6009, G6017, G6025, G6033, G6041,
    G6514, G6554, G6567, G6575, G6583, G6591, G6599, G6607, G6615, G6623,
    G6631, G6853, G6861, G6869, G6877, G6885, G6893, G6901, G6909, G6917,
    G784, G1014, G3221, G4913, G4929, G5183, G5231, G6511, G615, G594,
    G611, G617, G619, G621, G623, G625, G627, G664, G685, G691, G693, G695,
    G697, G699, G701, G703, G705, G707, G709, G4879, G4880, G4887, G4895,
    G4911, G4920, G4927, G5181, G5182, G5190, G5197, G5205, G5221, G5229,
    G1343, G1357, G1364, G1366, G1368, G1370, G1372, G1374, G1376, G1378,
    G1380, G1382, G5399, G5407, G5415, G5423, G5431, G5439, G5447, G5455,
    G5463, G5751, G5759, G5767, G5775, G5783, G5791, G5799, G5807, G5815,
    G2019, G2032, G2117, G2130, G2266, G2272, G2286, G2288, G2290, G2292,
    G2294, G5871, G5879, G5887, G5895, G5903, G5911, G5919, G5927, G5991,
    G5999, G6007, G6015, G6023, G6031, G6039, G6047, G2899, G2914, G2919,
    G2921, G2923, G2925, G2927, G2929, G2931, G6518, G3173, G6558, G6573,
    G6581, G6589, G6597, G6605, G6613, G6621, G6629, G6637, G3629, G3642,
    G3649, G3651, G3653, G3655, G3657, G3659, G3661, G3663, G3762, G3768,
    G3782, G3784, G3786, G3788, G3790, G6859, G6867, G6875, G6883, G6891,
    G6899, G6907, G6915, G6923, G4094, G4107, G4444, G4457, G4647, G4660,
    G4667, G4669, G4671, G4673, G4675, G4677, G4679, G4681, G4683, G4685,
    G4897, G5207, G6551, G763, G764, G4919, G886, G1005, G1006, G5189,
    G1018, G5237, G6517, G3169, G4935, G4970, G5239, G577, G616, G618,
    G620, G622, G624, G626, G628, G692, G694, G696, G698, G700, G702, G704,
    G706, G708, G710, G765, G4903, G885, G1007, G1017, G5213, G1363, G1365,
    G1367, G1369, G1371, G1373, G1375, G1377, G1379, G1381, G2026, G2039,
    G2046, G2048, G2050, G2052, G2054, G2056, G2058, G2060, G2062, G2064,
    G2124, G2137, G2144, G2146, G2148, G2150, G2152, G2154, G2156, G2158,
    G2160, G2162, G2279, G2285, G2287, G2289, G2291, G2293, G2296, G2298,
    G2300, G2302, G2304, G2918, G2920, G2922, G2924, G2926, G2928, G2930,
    G2932, G3168, G6557, G3211, G3648, G3650, G3652, G3654, G3656, G3658,
    G3660, G3662, G3665, G3666, G3775, G3781, G3783, G3785, G3787, G3789,
    G3792, G3794, G3796, G3798, G3800, G4101, G4114, G4123, G4126, G4129,
    G4132, G4135, G4138, G4141, G4144, G4147, G4150, G4451, G4464, G4471,
    G4473, G4475, G4477, G4479, G4481, G4483, G4485, G4487, G4489, G4666,
    G4668, G4670, G4672, G4674, G4676, G4678, G4680, G4682, G4684, G579,
    G629, G633, G637, G641, G645, G711, G715, G719, G723, G727, G731, G737,
    G745, G751, G757, G887, G1019, G5245, G1383, G1387, G1391, G1395,
    G1399, G1406, G1412, G1418, G2305, G2308, G2312, G2316, G2933, G2938,
    G2942, G2946, G2950, G3170, G3210, G3667, G3670, G3673, G3676, G3679,
    G3682, G3686, G3801, G3804, G3807, G3810, G3813, G4525, G4686, G4689,
    G4692, G4695, G4698, G4701, G4704, G4707, G4710, G4976, G5271, G5274,
    G5305, G5308, G5318, G6690, G6711, G6714, G7252, G7296, G7466, G907,
    G913, G915, G916, G1116, G2045, G2047, G2049, G2051, G2053, G2055,
    G2057, G2059, G2061, G2063, G2143, G2145, G2147, G2149, G2151, G2153,
    G2155, G2157, G2159, G2161, G2295, G2297, G2299, G2301, G2303, G3212,
    G3791, G3793, G3795, G3797, G3799, G4122, G4125, G4128, G4131, G4134,
    G4137, G4140, G4143, G4146, G4149, G4470, G4472, G4474, G4476, G4478,
    G4480, G4482, G4484, G4486, G4488, G4962, G5003, G5234, G5242, G5250,
    G5284, G802, G821, G845, G868, G877, G902, G908, G914, G917, G953,
    G1023, G1035, G1050, G1068, G1086, G1102, G1108, G1117, G5322, G1553,
    G1567, G1584, G1590, G1606, G1624, G1647, G1669, G1677, G1802, G1816,
    G1834, G1841, G1866, G1880, G1897, G1914, G1929, G2065, G2069, G2073,
    G2077, G2081, G2085, G2091, G2099, G2105, G2111, G2163, G2167, G2171,
    G2175, G2179, G2186, G2192, G2198, G2320, G2323, G2329, G2335, G2962,
    G2970, G2977, G2979, G2989, G2998, G3006, G3013, G3015, G3183, G3192,
    G3200, G3207, G3209, G3216, G3222, G6694, G3695, G3816, G3821, G3828,
    G3833, G3838, G4151, G4154, G4157, G4160, G4163, G4166, G4169, G4172,
    G4175, G7256, G7300, G4490, G4493, G4496, G4499, G4502, G4505, G4508,
    G4511, G7470, G4884, G4892, G4900, G4908, G4924, G4952, G4983, G4993,
    G5011, G5194, G5202, G5210, G5218, G5226, G5247, G5255, G5258, G5263,
    G5266, G5277, G5278, G5281, G5289, G5292, G5297, G5300, G5311, G5312,
    G5315, G5323, G5326, G5331, G5334, G5339, G5342, G5349, G5352, G5396,
    G5404, G5412, G5420, G5428, G5436, G5444, G5452, G5460, G5465, G5581,
    G5748, G5756, G5764, G5772, G5780, G5788, G5796, G5804, G5812, G5849,
    G5929, G6049, G6367, G6370, G6375, G6378, G6383, G6386, G6391, G6394,
    G6399, G6402, G6407, G6410, G6415, G6418, G6423, G6426, G6431, G6434,
    G6442, G6450, G6458, G6466, G6498, G6519, G6522, G6527, G6530, G6535,
    G6538, G6543, G6546, G6559, G6562, G6687, G6695, G6698, G6703, G6706,
    G6717, G6718, G6724, G6768, G7208, G7221, G7229, G7232, G7239, G7242,
    G7249, G7257, G7260, G7268, G7293, G7301, G7304, G7309, G7312, G7317,
    G7320, G7327, G7330, G7396, G7404, G7412, G7425, G7463, G7471, G7474,
    G7479, G7482, G7487, G7490, G7497, G7500, G7507, G7510, G7554, G1152,
    G5238, G1156, G5246, G5254, G5288, G3223, G4942, G4966, G5007, G5279,
    G5280, G5313, G5314, G6719, G6720, G790, G4888, G803, G4896, G825,
    G4904, G851, G4912, G893, G4928, G906, G912, G1024, G5198, G1036,
    G5206, G1053, G5214, G1072, G5222, G1091, G5230, G1112, G1121, G1153,
    G1157, G5253, G1216, G5261, G5262, G5269, G5270, G5287, G1239, G5295,
    G5296, G5303, G5304, G5321, G1262, G5329, G5330, G5337, G5338, G1544,
    G5400, G1554, G5408, G1571, G5416, G1596, G5424, G1607, G5432, G1628,
    G5440, G1653, G5448, G1685, G5456, G1693, G5464, G1793, G5752, G1803,
    G5760, G1820, G5768, G1848, G5776, G1857, G5784, G1867, G5792, G1883,
    G5800, G1901, G5808, G1919, G5816, G5855, G2351, G2366, G2384, G2391,
    G2417, G2431, G2448, G2465, G5935, G2597, G2612, G2629, G2635, G2652,
    G2670, G2693, G2715, G6055, G6373, G6374, G6381, G6382, G6389, G6390,
    G6397, G6398, G6405, G6406, G6413, G6414, G6421, G6422, G6429, G6430,
    G6437, G6438, G6446, G3059, G6454, G3068, G6462, G3076, G3079, G6470,
    G3090, G3099, G3107, G3114, G3116, G6502, G6525, G6526, G6533, G6534,
    G6541, G6542, G6549, G6550, G6565, G6566, G3220, G3292, G3308, G3327,
    G3335, G3362, G3376, G3393, G3410, G3425, G6693, G3503, G6701, G6702,
    G6709, G6710, G6728, G6772, G3853, G3868, G3885, G3891, G3908, G3926,
    G3949, G3971, G3979, G7212, G7227, G7255, G4202, G7263, G7264, G7272,
    G7299, G4225, G7307, G7308, G7315, G7316, G4297, G4305, G4312, G4314,
    G4324, G7400, G4333, G7408, G4341, G7416, G4348, G4349, G7431, G4389,
    G7469, G4530, G7477, G7478, G7485, G7486, G7513, G7514, G7558, G4932,
    G4956, G4973, G4987, G4997, G5017, G5099, G5345, G5346, G5355, G5356,
    G5372, G5380, G5471, G5523, G5587, G5669, G5857, G5868, G5876, G5884,
    G5892, G5900, G5908, G5916, G5924, G5969, G5988, G5996, G6004, G6012,
    G6020, G6028, G6036, G6044, G6057, G6439, G6447, G6455, G6463, G6471,
    G6474, G6479, G6482, G6487, G6490, G6495, G6503, G6506, G6570, G6578,
    G6586, G6594, G6602, G6610, G6618, G6626, G6634, G6671, G6721, G6729,
    G6732, G6737, G6740, G6745, G6748, G6755, G6758, G6765, G6773, G6776,
    G6781, G6784, G6789, G6792, G6799, G6802, G6832, G6856, G6864, G6872,
    G6880, G6888, G6896, G6904, G6912, G6920, G6925, G7041, G7205, G7213,
    G7216, G7224, G7235, G7236, G7245, G7246, G7265, G7273, G7276, G7283,
    G7286, G7323, G7324, G7333, G7334, G7361, G7364, G7369, G7372, G7377,
    G7380, G7385, G7388, G7393, G7401, G7409, G7417, G7420, G7428, G7493,
    G7494, G7503, G7504, G7515, G7518, G7523, G7526, G7531, G7534, G7541,
    G7544, G7551, G7559, G7562, G7567, G7570, G7575, G7578, G7585, G7588,
    G1176, G957, G791, G804, G826, G852, G894, G1025, G1037, G1054, G1073,
    G1092, G1154, G1158, G1215, G1224, G1225, G1233, G1234, G1238, G1247,
    G1248, G1256, G1257, G1261, G1270, G1271, G1279, G1280, G1545, G1555,
    G1572, G1597, G1608, G1629, G1654, G1686, G1694, G1794, G1804, G1821,
    G1849, G1858, G1868, G1884, G1902, G1920, G2954, G2955, G2963, G2964,
    G2971, G2972, G2980, G2981, G2990, G2991, G2999, G3000, G3007, G3008,
    G3016, G3017, G3019, G3020, G3174, G3175, G3184, G3185, G3193, G3194,
    G3201, G3202, G3213, G3214, G3227, G3502, G3511, G3512, G3520, G3521,
    G4201, G4210, G4211, G4224, G4233, G4234, G4242, G4243, G4529, G4538,
    G4539, G4547, G4548, G4552, G4553, G4946, G5347, G5348, G5357, G5358,
    G7237, G7238, G7247, G7248, G7325, G7326, G7335, G7336, G7495, G7496,
    G7505, G7506, G3244, G792, G805, G827, G853, G895, G1026, G1038, G1055,
    G1074, G1093, G1155, G1217, G1226, G1235, G1240, G1249, G1258, G1263,
    G1272, G1281, G5376, G5384, G1546, G1556, G1573, G1598, G1609, G1630,
    G1655, G1687, G1695, G1795, G1805, G1822, G1850, G1859, G1869, G1885,
    G1903, G1921, G5863, G2341, G5872, G2352, G5880, G2370, G5888, G2398,
    G5896, G2407, G5904, G2418, G5912, G2434, G5920, G2452, G5928, G2481,
    G5975, G2587, G5992, G2598, G6000, G2616, G6008, G2641, G6016, G2653,
    G6024, G2674, G6032, G2699, G6040, G2724, G2732, G6048, G2956, G2965,
    G2973, G2982, G2992, G3001, G3009, G3018, G3021, G6445, G3051, G6453,
    G3061, G6461, G3070, G6469, G3081, G6477, G6478, G6485, G6486, G6493,
    G6494, G6501, G3118, G6509, G6510, G3176, G3186, G3195, G3203, G3215,
    G3281, G6574, G3293, G6582, G3312, G6590, G3342, G6598, G3351, G6606,
    G3363, G6614, G3379, G6622, G3397, G6630, G3415, G6638, G6677, G3504,
    G3513, G3522, G6727, G3526, G6735, G6736, G6743, G6744, G6771, G3549,
    G6779, G6780, G6787, G6788, G6836, G3843, G6860, G3854, G6868, G3872,
    G6876, G3897, G6884, G3909, G6892, G3930, G6900, G3955, G6908, G3987,
    G6916, G3995, G6924, G7211, G4179, G7219, G7220, G4196, G7228, G4203,
    G4212, G7271, G4220, G4226, G4235, G4244, G7367, G7368, G7375, G7376,
    G7383, G7384, G7391, G7392, G7399, G4326, G7407, G4335, G7415, G4343,
    G7423, G7424, G4353, G7432, G4531, G4540, G4549, G4554, G7521, G7522,
    G7529, G7530, G7557, G4576, G7565, G7566, G7573, G7574, G4936, G4937,
    G4977, G4978, G5105, G5359, G5362, G5529, G5675, G5932, G5977, G6052,
    G6063, G6115, G6173, G6679, G6751, G6752, G6761, G6762, G6795, G6796,
    G6805, G6806, G6931, G6983, G7047, G7129, G7279, G7280, G7289, G7290,
    G7337, G7340, G7353, G7356, G7537, G7538, G7547, G7548, G7581, G7582,
    G7591, G7592, G7595, G7598, G2342, G2353, G2371, G2399, G2408, G2419,
    G2435, G2453, G2588, G2599, G2617, G2642, G2654, G2675, G2700, G2733,
    G3050, G3060, G3069, G3080, G3091, G3092, G3100, G3101, G3108, G3109,
    G3117, G3120, G3121, G3282, G3294, G3313, G3343, G3352, G3364, G3380,
    G3398, G3416, G3525, G3534, G3535, G3543, G3544, G3548, G3557, G3558,
    G3566, G3567, G3844, G3855, G3873, G3898, G3910, G3931, G3956, G3988,
    G3996, G4178, G4187, G4188, G4197, G4219, G4289, G4290, G4298, G4299,
    G4306, G4307, G4315, G4316, G4325, G4334, G4342, G4350, G4351, G4354,
    G4561, G4562, G4570, G4571, G4575, G4584, G4585, G4593, G4594, G4938,
    G4979, G6753, G6754, G6763, G6764, G6797, G6798, G6807, G6808, G7281,
    G7282, G7291, G7292, G7539, G7540, G7549, G7550, G7583, G7584, G7593,
    G7594, G1856, G920, G925, G926, G927, G928, G937, G938, G939, G940,
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G956, G1122,
    G1125, G1126, G1127, G1128, G1132, G1133, G1134, G1137, G1138, G1141,
    G1221, G1230, G1244, G1253, G1267, G1276, G1284, G1288, G1292, G1296,
    G1300, G1304, G1702, G1705, G1706, G1707, G1709, G1710, G1711, G1712,
    G1713, G1714, G1718, G1722, G1723, G1724, G1725, G1733, G1734, G1735,
    G1736, G1737, G1738, G1739, G1740, G1741, G1742, G1743, G1744, G1745,
    G1749, G1750, G1935, G1938, G1939, G1940, G1942, G1943, G1944, G1945,
    G1946, G1947, G1948, G1949, G1950, G1953, G1954, G1955, G1956, G1960,
    G1961, G1962, G1965, G1966, G1969, G2343, G2354, G2372, G2400, G2409,
    G2420, G2436, G2454, G2470, G5936, G5983, G2589, G2600, G2618, G2643,
    G2655, G2676, G2701, G2734, G2740, G6056, G3022, G3025, G3026, G3027,
    G3029, G3030, G3031, G3032, G3033, G3052, G3062, G3071, G3082, G3093,
    G3102, G3110, G3119, G3122, G3228, G3231, G3232, G3233, G3234, G3283,
    G3295, G3314, G3344, G3353, G3365, G3381, G3399, G3417, G6685, G3508,
    G3517, G3527, G3536, G3545, G3550, G3559, G3568, G3571, G3575, G3845,
    G3856, G3874, G3899, G3911, G3932, G3957, G3989, G3997, G4180, G4189,
    G4198, G4207, G4216, G4221, G4230, G4239, G4263, G4267, G4291, G4300,
    G4308, G4317, G4327, G4336, G4344, G4352, G4355, G4535, G4544, G4558,
    G4563, G4572, G4577, G4586, G4595, G4598, G4602, G4716, G4724, G4732,
    G4740, G4748, G4756, G4764, G4772, G4780, G4788, G4939, G4980, G5044,
    G5054, G5064, G5074, G5084, G5094, G5132, G5142, G5152, G5162, G5365,
    G5366, G5488, G5498, G5508, G5518, G5546, G5556, G5566, G5576, G5614,
    G5624, G5634, G5644, G5654, G5664, G5702, G5712, G5722, G5732, G5820,
    G5828, G5836, G5844, G5852, G5860, G6121, G6179, G6261, G7359, G7360,
    G7343, G7344, G6809, G6812, G6819, G6822, G6989, G7135, G7345, G7348,
    G7601, G7602, G7603, G7606, G7611, G7614, G929, G950, G1129, G1708,
    G1715, G1726, G1746, G1941, G1957, G2471, G2741, G3028, G3034, G3235,
    G5014, G5034, G5102, G5122, G5367, G5368, G5478, G5536, G5584, G5604,
    G5672, G5692, G5817, G5825, G5833, G5841, G6340, G6341, G6350, G6351,
    G7436, G7437, G4720, G4728, G4736, G4744, G4752, G4760, G4768, G4776,
    G4784, G4792, G3350, G2406, G924, G5088, G5098, G997, G1146, G1287,
    G1291, G1295, G1299, G1303, G1307, G1309, G1312, G1315, G1318, G1321,
    G1324, G1721, G5522, G5580, G5658, G5668, G1788, G1974, G5824, G5832,
    G5840, G5848, G1999, G5856, G2003, G5864, G2472, G2487, G2492, G2493,
    G2494, G2500, G2501, G2502, G2503, G2504, G2505, G2506, G2507, G2511,
    G2512, G2513, G2514, G2518, G2519, G2520, G2523, G2524, G2527, G2742,
    G2749, G2754, G2755, G2756, G2762, G2763, G2764, G2765, G2766, G2767,
    G2776, G2777, G2778, G2779, G2788, G2789, G2790, G2792, G2793, G2794,
    G2795, G2796, G2798, G2799, G2800, G2804, G3035, G3045, G3123, G3128,
    G3129, G3130, G3136, G3139, G3140, G3141, G3142, G3249, G3431, G3434,
    G3435, G3436, G3438, G3439, G3440, G3441, G3442, G3443, G3444, G3445,
    G3446, G3449, G3450, G3451, G3452, G3456, G3457, G3458, G3460, G3461,
    G3463, G3531, G3540, G3554, G3563, G3574, G3578, G3579, G3583, G3587,
    G3591, G3596, G3599, G4004, G4007, G4008, G4009, G4011, G4012, G4013,
    G4014, G4015, G4016, G4020, G4024, G4025, G4026, G4027, G4035, G4036,
    G4037, G4038, G4039, G4040, G4041, G4042, G4043, G4044, G4045, G4046,
    G4047, G4051, G4052, G4184, G4193, G4247, G4251, G4255, G4259, G4266,
    G4270, G4284, G4287, G4356, G4361, G4362, G4363, G4369, G4372, G4373,
    G4374, G4375, G4567, G4581, G4590, G4601, G4605, G4606, G4610, G4614,
    G4618, G4623, G4626, G4796, G4804, G4812, G4820, G4828, G4844, G4852,
    G4860, G4868, G4945, G4948, G4986, G4989, G5048, G5058, G5068, G5078,
    G5166, G5136, G5146, G5156, G5388, G5492, G5502, G5512, G5550, G5560,
    G5570, G5618, G5628, G5638, G5648, G5736, G5706, G5716, G5726, G5940,
    G5948, G5956, G5964, G5972, G5980, G6080, G6090, G6100, G6110, G6138,
    G6148, G6158, G6168, G6216, G6226, G6236, G6246, G6256, G6267, G6304,
    G6314, G6324, G6342, G6352, G7351, G7352, G6642, G6650, G6658, G6666,
    G6674, G6682, G6815, G6816, G6825, G6826, G6948, G6958, G6968, G6978,
    G7006, G7016, G7026, G7036, G7074, G7084, G7094, G7104, G7114, G7124,
    G7162, G7172, G7182, G7192, G7438, G7617, G7618, G7609, G7610, G1151,
    G1002, G933, G1308, G1311, G1314, G1317, G1320, G1323, G1730, G1789,
    G1981, G5823, G1986, G5831, G1989, G5839, G1993, G5847, G1996, G2000,
    G2004, G2495, G2515, G2757, G2768, G2780, G2801, G3046, G3131, G3143,
    G3238, G3258, G3437, G3453, G3595, G3598, G4010, G4017, G4028, G4048,
    G4283, G4286, G4364, G4376, G4622, G4625, G4947, G4988, G5018, G5019,
    G5024, G5038, G5106, G5107, G5112, G5126, G5468, G5482, G5526, G5540,
    G5588, G5589, G5594, G5608, G5676, G5677, G5682, G5696, G5937, G5945,
    G5953, G5961, G6070, G6128, G6264, G6284, G6360, G6361, G6639, G6647,
    G6655, G6663, G6817, G6818, G6827, G6828, G6938, G6996, G7044, G7064,
    G7132, G7152, G7446, G7447, G7456, G7457, G241, G265, G2005, G4800,
    G4808, G4816, G4824, G4832, G4848, G4856, G4864, G4872, G1310, G1313,
    G1316, G1319, G1322, G1325, G5392, G1790, G1982, G1985, G1988, G1992,
    G1995, G2001, G2491, G2508, G2522, G2526, G2529, G2531, G5944, G5952,
    G5960, G5968, G2555, G5976, G2559, G5984, G2753, G2771, G2791, G2797,
    G2807, G6114, G6172, G6250, G6260, G6346, G6356, G3127, G3156, G3259,
    G3466, G6646, G6654, G6662, G6670, G3483, G6678, G3487, G6686, G3582,
    G3586, G3590, G3594, G3597, G3600, G3602, G3605, G3608, G3611, G4023,
    G6982, G7040, G7118, G7128, G4089, G4250, G4254, G4258, G4262, G4272,
    G4275, G4278, G4281, G4285, G4288, G4360, G4380, G4386, G7442, G4609,
    G4613, G4617, G4621, G4624, G4627, G4629, G4632, G4635, G4638, G4836,
    G4949, G4990, G5020, G5108, G5590, G5678, G6084, G6094, G6104, G6142,
    G6152, G6162, G6206, G6220, G6230, G6240, G6328, G6294, G6308, G6318,
    G6362, G6840, G6848, G6952, G6962, G6972, G7010, G7020, G7030, G7078,
    G7088, G7098, G7108, G7196, G7166, G7176, G7186, G7448, G7458, G254,
    G260, G1987, G1994, G2002, G962, G1751, G1990, G1997, G2499, G2536,
    G5943, G2542, G5951, G2545, G5959, G2549, G5967, G2552, G2556, G2560,
    G2761, G2784, G2853, G3135, G3146, G3163, G3467, G6645, G3470, G6653,
    G3473, G6661, G3477, G6669, G3480, G3484, G3488, G3601, G3604, G3607,
    G3610, G4032, G4090, G4271, G4274, G4277, G4280, G4368, G4379, G4387,
    G4628, G4631, G4634, G4637, G4841, G4849, G4857, G4865, G5021, G5028,
    G5109, G5116, G5369, G5377, G5385, G5472, G5473, G5530, G5531, G5591,
    G5598, G5679, G5686, G6060, G6074, G6118, G6132, G6176, G6186, G6196,
    G6268, G6269, G6274, G6288, G6337, G6829, G6928, G6942, G6986, G7000,
    G7048, G7049, G7054, G7068, G7136, G7137, G7142, G7156, G7433, G242,
    G3151, G257, G263, G266, G1991, G1998, G3489, G371, G4840, G2561,
    G2532, G2537, G2541, G2544, G2548, G2551, G2557, G2563, G2577, G2775,
    G2806, G2808, G2852, G2854, G6366, G4381, G3164, G3241, G3468, G3469,
    G3472, G3476, G3479, G3485, G3603, G3606, G3609, G3612, G6844, G6852,
    G4091, G4273, G4276, G4279, G4282, G4382, G4388, G7452, G7462, G4630,
    G4633, G4636, G4639, G4955, G4958, G4996, G4999, G5474, G5532, G6210,
    G6270, G6298, G7050, G7138, G3471, G3478, G3486, G372, G2543, G2550,
    G2558, G4847, G387, G4855, G390, G4863, G393, G4871, G396, G965, G5375,
    G1327, G5383, G1330, G5391, G1333, G1754, G2546, G2553, G2564, G2809,
    G2813, G6345, G2860, G3474, G3481, G6835, G3614, G4053, G7441, G4516,
    G4957, G4998, G5027, G5030, G5115, G5118, G5475, G5533, G5597, G5600,
    G5685, G5688, G6064, G6065, G6122, G6123, G6180, G6181, G6190, G6200,
    G6271, G6278, G6347, G6357, G6837, G6845, G6932, G6933, G6990, G6991,
    G7051, G7058, G7139, G7146, G7443, G7453, G243, G244, G245, G255, G256,
    G261, G262, G267, G268, G269, G3475, G3482, G2547, G2554, G386, G389,
    G392, G395, G1326, G1329, G1332, G1436, G1440, G1445, G1450, G1454,
    G2859, G4385, G3148, G3239, G3240, G3265, G3267, G3270, G3274, G3277,
    G3613, G4515, G4959, G5000, G5029, G5117, G5599, G5687, G6066, G6124,
    G6182, G6934, G6992, G375, G378, G381, G384, G1328, G1331, G1334,
    G1447, G1766, G2571, G2579, G2812, G2816, G2851, G2861, G6355, G2863,
    G6365, G2866, G3147, G3242, G3271, G3279, G3615, G6843, G3617, G6851,
    G3620, G4056, G4517, G7451, G4519, G7461, G4522, G5031, G5119, G5481,
    G5484, G5539, G5542, G5601, G5689, G6067, G6125, G6183, G6277, G6280,
    G6935, G6993, G7057, G7060, G7145, G7148, G4968, G5009, G2850, G2862,
    G2865, G3149, G3243, G3616, G3619, G4518, G4521, G4965, G5006, G5483,
    G5541, G6279, G7059, G7147, G374, G377, G380, G383, G955, G4967, G5008,
    G975, G1136, G1140, G1143, G1145, G1160, G1771, G1964, G1968, G1971,
    G1973, G2007, G2578, G2864, G2867, G3150, G3245, G3618, G3621, G4067,
    G4520, G4523, G4713, G4753, G5037, G5040, G5125, G5128, G5485, G5543,
    G5607, G5610, G5695, G5698, G6073, G6076, G6131, G6134, G6189, G6192,
    G6281, G6941, G6944, G6999, G7002, G7061, G7149, G958, G967, G971,
    G1161, G2008, G2580, G2868, G3152, G4443, G4524, G4721, G4729, G4737,
    G4745, G4761, G4769, G4777, G4785, G5039, G5127, G5609, G5697, G6075,
    G6133, G6191, G6943, G7001, G3248, G248, G4719, G294, G4759, G323,
    G980, G4072, G5041, G5129, G5491, G5494, G5549, G5552, G5611, G5699,
    G6077, G6135, G6193, G6287, G6290, G6945, G7003, G7067, G7070, G7155,
    G7158, G247, G3155, G251, G272, G961, G275, G293, G297, G300, G303,
    G306, G4727, G309, G4735, G312, G4743, G315, G4751, G318, G322, G4767,
    G326, G4775, G329, G4783, G332, G4791, G335, G2881, G993, G994, G1166,
    G1171, G1174, G2014, G3459, G3462, G3464, G3465, G3490, G4793, G5493,
    G5551, G6289, G7069, G7157, G250, G274, G308, G311, G314, G317, G325,
    G328, G331, G334, G417, G991, G992, G3491, G4801, G4809, G4817, G4825,
    G5047, G5050, G5135, G5138, G5495, G5553, G5617, G5620, G5705, G5708,
    G6083, G6086, G6141, G6144, G6199, G6202, G6291, G6951, G6954, G7009,
    G7012, G7071, G7159, G271, G296, G299, G302, G305, G4799, G343, G1170,
    G1173, G5049, G5137, G5167, G5619, G5707, G6085, G6143, G6201, G6953,
    G7011, G342, G346, G349, G352, G355, G4807, G358, G4815, G361, G4823,
    G364, G4831, G367, G1172, G1175, G3497, G5051, G5139, G5501, G5504,
    G5559, G5562, G5621, G5709, G6087, G6145, G6203, G6297, G6300, G6955,
    G7013, G7077, G7080, G7165, G7168, G357, G360, G363, G366, G5173,
    G5503, G5561, G6299, G7079, G7167, G345, G348, G351, G354, G5057,
    G5060, G5145, G5148, G5505, G5563, G5627, G5630, G5715, G5718, G6093,
    G6096, G6151, G6154, G6209, G6212, G6301, G6961, G6964, G7019, G7022,
    G7081, G7169, G5059, G5147, G5629, G5717, G6095, G6153, G6211, G6963,
    G7021, G5061, G5149, G5511, G5514, G5569, G5572, G5631, G5719, G6097,
    G6155, G6213, G6307, G6310, G6965, G7023, G7087, G7090, G7175, G7178,
    G5513, G5571, G6309, G7089, G7177, G5067, G5070, G5155, G5158, G5515,
    G5573, G5637, G5640, G5725, G5728, G6103, G6106, G6161, G6164, G6219,
    G6222, G6311, G6971, G6974, G7029, G7032, G7091, G7179, G5069, G5157,
    G5639, G5727, G6105, G6163, G6221, G6973, G7031, G5521, G1756, G5579,
    G1761, G5071, G5159, G5641, G5729, G6107, G6165, G6223, G6317, G6320,
    G6975, G7033, G7097, G7100, G7185, G7188, G1755, G1760, G6319, G7099,
    G7187, G1757, G1762, G6113, G2818, G6171, G2823, G6981, G4058, G7039,
    G4063, G5077, G5080, G5165, G5090, G5647, G5650, G5735, G5660, G6229,
    G6232, G6321, G7101, G7189, G2817, G2822, G4057, G4062, G5079, G5089,
    G5649, G5659, G6231, G1782, G1783, G1784, G1785, G2819, G2824, G4059,
    G4064, G5081, G5091, G5651, G5661, G6233, G6327, G6252, G7107, G7110,
    G7195, G7120, G5737, G6251, G7109, G7119, G5087, G985, G5097, G988,
    G5657, G1776, G5667, G1779, G2844, G2845, G2846, G2847, G4083, G4084,
    G4085, G4086, G6239, G6242, G6253, G7111, G7121, G984, G987, G1775,
    G1778, G5743, G6241, G6329, G7197, G986, G989, G1777, G1780, G6259,
    G2841, G7117, G4077, G7127, G4080, G6243, G990, G996, G1781, G1787,
    G2840, G6335, G4076, G4079, G7203, G995, G1786, G6249, G2838, G2842,
    G4078, G4081, G2837, G2843, G4082, G4088, G5170, G5740, G2839, G2848,
    G4087, G1791, G1003, G5174, G5744, G2849, G7200, G1792, G1004, G6332,
    G320, G337, G4092, G7204, G4093, G2855, G6336, G369, G2856, G398;
  assign G2 = G1;
  assign G3 = G1;
  assign G400 = ~G57;
  assign G1184 = G134 & G133;
  assign G450 = G1459;
  assign G448 = G1469;
  assign G444 = G1480;
  assign G442 = G1486;
  assign G440 = G1492;
  assign G438 = G1496;
  assign G1501 = G199 & G188 & G162 & G172;
  assign G496 = G2208;
  assign G494 = G2218;
  assign G492 = G2224;
  assign G490 = G2230;
  assign G488 = G2236;
  assign G486 = G2239;
  assign G484 = G2247;
  assign G482 = G2253;
  assign G480 = G2256;
  assign G2857 = G240 & G228 & G150 & G184;
  assign G560 = G3698;
  assign G542 = G3701;
  assign G558 = G3705;
  assign G556 = G3711;
  assign G554 = G3717;
  assign G552 = G3723;
  assign G550 = G3729;
  assign G548 = G3737;
  assign G546 = G3743;
  assign G544 = G3749;
  assign G540 = G4393;
  assign G538 = G4400;
  assign G536 = G4405;
  assign G534 = G4410;
  assign G532 = G4415;
  assign G530 = G4420;
  assign G528 = G4427;
  assign G526 = G4432;
  assign G524 = G4437;
  assign G4442 = G186 & G185 & G183 & G182;
  assign G4514 = G230 & G218 & G210 & G152;
  assign G279 = ~G15;
  assign G401 = ~G5;
  assign G573 = G1;
  assign G574 = ~G5;
  assign G575 = ~G5;
  assign G1178 = ~G2236;
  assign G1186 = ~G2253;
  assign G1192 = ~G2256;
  assign G1198 = G38;
  assign G1205 = G15;
  assign G1206 = ~G12 | ~G9;
  assign G1207 = ~G12 | ~G9;
  assign G1210 = G38;
  assign G1458 = ~G1455;
  assign G1461 = ~G1459;
  assign G436 = G1462;
  assign G1464 = ~G1462;
  assign G1471 = ~G1469;
  assign G1475 = G106;
  assign G1482 = ~G1480;
  assign G1488 = ~G1486;
  assign G1495 = ~G1492;
  assign G1499 = ~G1496;
  assign G1500 = ~G106;
  assign G1503 = G18;
  assign G1512 = G18;
  assign G1518 = G4528 & G1492;
  assign G1524 = G18;
  assign G1535 = ~G18;
  assign G1541 = ~G4528 | ~G1496;
  assign G2207 = ~G2204;
  assign G2210 = ~G2208;
  assign G478 = G2211;
  assign G2213 = ~G2211;
  assign G2220 = ~G2218;
  assign G2226 = ~G2224;
  assign G2232 = ~G2230;
  assign G2238 = ~G2236;
  assign G2241 = ~G2239;
  assign G2249 = ~G2247;
  assign G2255 = ~G2253;
  assign G2258 = ~G2256;
  assign G2828 = G4526;
  assign G3700 = ~G3698;
  assign G3703 = ~G3701;
  assign G3707 = ~G3705;
  assign G3713 = ~G3711;
  assign G3719 = ~G3717;
  assign G3725 = ~G3723;
  assign G3731 = ~G3729;
  assign G3739 = ~G3737;
  assign G3745 = ~G3743;
  assign G3751 = ~G3749;
  assign G4121 = ~G4393;
  assign G522 = G4394;
  assign G4396 = ~G4394;
  assign G4402 = ~G4400;
  assign G4407 = ~G4405;
  assign G4412 = ~G4410;
  assign G4417 = ~G4415;
  assign G4422 = ~G4420;
  assign G4429 = ~G4427;
  assign G4434 = ~G4432;
  assign G4439 = ~G4437;
  assign G4833 = G4526;
  assign G402 = ~G400 | ~G401;
  assign G404 = ~G2857;
  assign G406 = ~G4514;
  assign G408 = ~G4442;
  assign G410 = ~G1501;
  assign G2876 = G2857 & G4514;
  assign G2878 = G4442 & G1501;
  assign G432 = G573;
  assign G446 = G1475;
  assign G1519 = ~G1518;
  assign G2871 = G4528 & G1458;
  assign G2883 = ~G4528 | ~G2207;
  assign G280 = G1184 & G575;
  assign G284 = ~G1197 | ~G574;
  assign G286 = ~G1205;
  assign G289 = ~G1197 | ~G574;
  assign G292 = ~G1184 | ~G575;
  assign G341 = ~G1205;
  assign G4839 = ~G4833;
  assign G572 = G573;
  assign G581 = G1206;
  assign G587 = G1512;
  assign G601 = G1206;
  assign G606 = G1512;
  assign G650 = G1206;
  assign G657 = G1512;
  assign G671 = G1207;
  assign G678 = G1503;
  assign G777 = G1541 & G1198;
  assign G1115 = G1541 & G1198;
  assign G1336 = G1512;
  assign G1350 = G1503;
  assign G1477 = ~G1475;
  assign G1507 = ~G1503;
  assign G1514 = ~G1512;
  assign G1530 = ~G1524;
  assign G2259 = G1535;
  assign G2833 = ~G2828;
  assign G2872 = ~G2871;
  assign G2886 = G1207;
  assign G2892 = G1503;
  assign G2905 = G1207;
  assign G2909 = G1503;
  assign G3622 = G1524;
  assign G3635 = G1524;
  assign G3755 = G1535;
  assign G4640 = G1524;
  assign G4653 = G1524;
  assign G4873 = G1541;
  assign G4876 = G1198;
  assign G4881 = G1488;
  assign G4889 = G1482;
  assign G4905 = G1471;
  assign G4916 = G1198;
  assign G4921 = G1464;
  assign G5175 = G1541;
  assign G5178 = G1198;
  assign G5186 = G1198;
  assign G5191 = G1488;
  assign G5199 = G1482;
  assign G5215 = G1471;
  assign G5223 = G1464;
  assign G5393 = G1192;
  assign G5401 = G1186;
  assign G5409 = G2249;
  assign G5417 = G1178;
  assign G5425 = G2232;
  assign G5433 = G2226;
  assign G5441 = G2220;
  assign G5449 = G2241;
  assign G5457 = G2213;
  assign G5745 = G1192;
  assign G5753 = G1186;
  assign G5761 = G2249;
  assign G5769 = G2241;
  assign G5777 = G1178;
  assign G5785 = G2232;
  assign G5793 = G2226;
  assign G5801 = G2220;
  assign G5809 = G2213;
  assign G5865 = G3751;
  assign G5873 = G3745;
  assign G5881 = G3739;
  assign G5889 = G3731;
  assign G5897 = G3725;
  assign G5905 = G3719;
  assign G5913 = G3713;
  assign G5921 = G3707;
  assign G5985 = G3751;
  assign G5993 = G3745;
  assign G6001 = G3739;
  assign G6009 = G3725;
  assign G6017 = G3719;
  assign G6025 = G3713;
  assign G6033 = G3707;
  assign G6041 = G3731;
  assign G6514 = G1210;
  assign G6554 = G1210;
  assign G6567 = G4439;
  assign G6575 = G4434;
  assign G6583 = G4429;
  assign G6591 = G4422;
  assign G6599 = G4417;
  assign G6607 = G4412;
  assign G6615 = G4407;
  assign G6623 = G4402;
  assign G6631 = G4396;
  assign G6853 = G4439;
  assign G6861 = G4434;
  assign G6869 = G4429;
  assign G6877 = G4417;
  assign G6885 = G4412;
  assign G6893 = G4407;
  assign G6901 = G4402;
  assign G6909 = G4422;
  assign G6917 = G4396;
  assign G281 = ~G280;
  assign G453 = G572;
  assign G784 = G1519 & G1198;
  assign G1014 = G1198 & G1519;
  assign G3221 = G2883 & G1210;
  assign G4913 = G1519;
  assign G4929 = ~G1519 & ~G1198;
  assign G5183 = G1519;
  assign G5231 = ~G1198 & ~G1519;
  assign G6511 = G2883;
  assign G278 = G163 & G572;
  assign G615 = G170 & G587;
  assign G594 = ~G587;
  assign G611 = ~G606;
  assign G617 = G169 & G587;
  assign G619 = G168 & G587;
  assign G621 = G167 & G587;
  assign G623 = G166 & G606;
  assign G625 = G165 & G606;
  assign G627 = G164 & G606;
  assign G664 = ~G657;
  assign G685 = ~G678;
  assign G691 = G177 & G657;
  assign G693 = G176 & G657;
  assign G695 = G175 & G657;
  assign G697 = G174 & G657;
  assign G699 = G173 & G657;
  assign G701 = G157 & G678;
  assign G703 = G156 & G678;
  assign G705 = G155 & G678;
  assign G707 = G154 & G678;
  assign G709 = G153 & G678;
  assign G4879 = ~G4873;
  assign G4880 = ~G4876;
  assign G4887 = ~G4881;
  assign G4895 = ~G4889;
  assign G4911 = ~G4905;
  assign G4920 = ~G4916;
  assign G4927 = ~G4921;
  assign G5181 = ~G5175;
  assign G5182 = ~G5178;
  assign G5190 = ~G5186;
  assign G5197 = ~G5191;
  assign G5205 = ~G5199;
  assign G5221 = ~G5215;
  assign G5229 = ~G5223;
  assign G1343 = ~G1336;
  assign G1357 = ~G1350;
  assign G1364 = G181 & G1336;
  assign G1366 = G171 & G1336;
  assign G1368 = G180 & G1336;
  assign G1370 = G179 & G1336;
  assign G1372 = G178 & G1336;
  assign G1374 = G161 & G1350;
  assign G1376 = G151 & G1350;
  assign G1378 = G160 & G1350;
  assign G1380 = G159 & G1350;
  assign G1382 = G158 & G1350;
  assign G5399 = ~G5393;
  assign G5407 = ~G5401;
  assign G5415 = ~G5409;
  assign G5423 = ~G5417;
  assign G5431 = ~G5425;
  assign G5439 = ~G5433;
  assign G5447 = ~G5441;
  assign G5455 = ~G5449;
  assign G5463 = ~G5457;
  assign G5751 = ~G5745;
  assign G5759 = ~G5753;
  assign G5767 = ~G5761;
  assign G5775 = ~G5769;
  assign G5783 = ~G5777;
  assign G5791 = ~G5785;
  assign G5799 = ~G5793;
  assign G5807 = ~G5801;
  assign G5815 = ~G5809;
  assign G2019 = G1514;
  assign G2032 = G1507;
  assign G2117 = G1514;
  assign G2130 = G1507;
  assign G2266 = ~G2259;
  assign G2272 = G1507;
  assign G2286 = G44 & G2259;
  assign G2288 = G41 & G2259;
  assign G2290 = G29 & G2259;
  assign G2292 = G26 & G2259;
  assign G2294 = G23 & G2259;
  assign G5871 = ~G5865;
  assign G5879 = ~G5873;
  assign G5887 = ~G5881;
  assign G5895 = ~G5889;
  assign G5903 = ~G5897;
  assign G5911 = ~G5905;
  assign G5919 = ~G5913;
  assign G5927 = ~G5921;
  assign G5991 = ~G5985;
  assign G5999 = ~G5993;
  assign G6007 = ~G6001;
  assign G6015 = ~G6009;
  assign G6023 = ~G6017;
  assign G6031 = ~G6025;
  assign G6039 = ~G6033;
  assign G6047 = ~G6041;
  assign G2899 = ~G2892;
  assign G2914 = ~G2909;
  assign G2919 = G209 & G2892;
  assign G2921 = G216 & G2892;
  assign G2923 = G215 & G2892;
  assign G2925 = G214 & G2892;
  assign G2927 = G213 & G2909;
  assign G2929 = G212 & G2909;
  assign G2931 = G211 & G2909;
  assign G6518 = ~G6514;
  assign G3173 = G2872 & G1210;
  assign G6558 = ~G6554;
  assign G6573 = ~G6567;
  assign G6581 = ~G6575;
  assign G6589 = ~G6583;
  assign G6597 = ~G6591;
  assign G6605 = ~G6599;
  assign G6613 = ~G6607;
  assign G6621 = ~G6615;
  assign G6629 = ~G6623;
  assign G6637 = ~G6631;
  assign G3629 = ~G3622;
  assign G3642 = ~G3635;
  assign G3649 = G1461 & G3622;
  assign G3651 = G1464 & G3622;
  assign G3653 = G1471 & G3622;
  assign G3655 = G1500 & G3622;
  assign G3657 = G1482 & G3622;
  assign G3659 = G1488 & G3635;
  assign G3661 = G1495 & G3635;
  assign G3663 = G1499 & G3635;
  assign G3762 = ~G3755;
  assign G3768 = G1507;
  assign G3782 = G47 & G3755;
  assign G3784 = G35 & G3755;
  assign G3786 = G32 & G3755;
  assign G3788 = G50 & G3755;
  assign G3790 = G66 & G3755;
  assign G6859 = ~G6853;
  assign G6867 = ~G6861;
  assign G6875 = ~G6869;
  assign G6883 = ~G6877;
  assign G6891 = ~G6885;
  assign G6899 = ~G6893;
  assign G6907 = ~G6901;
  assign G6915 = ~G6909;
  assign G6923 = ~G6917;
  assign G4094 = G1530;
  assign G4107 = G1530;
  assign G4444 = G1530;
  assign G4457 = G1530;
  assign G4647 = ~G4640;
  assign G4660 = ~G4653;
  assign G4667 = G2210 & G4640;
  assign G4669 = G2213 & G4640;
  assign G4671 = G2220 & G4640;
  assign G4673 = G2226 & G4640;
  assign G4675 = G2232 & G4640;
  assign G4677 = G2238 & G4653;
  assign G4679 = G2241 & G4653;
  assign G4681 = G2249 & G4653;
  assign G4683 = G2255 & G4653;
  assign G4685 = G2258 & G4653;
  assign G4897 = G1477;
  assign G5207 = G1477;
  assign G6551 = G2872;
  assign G763 = ~G4876 | ~G4879;
  assign G764 = ~G4873 | ~G4880;
  assign G4919 = ~G4913;
  assign G886 = ~G4913 | ~G4920;
  assign G1005 = ~G5178 | ~G5181;
  assign G1006 = ~G5175 | ~G5182;
  assign G5189 = ~G5183;
  assign G1018 = ~G5183 | ~G5190;
  assign G5237 = ~G5231;
  assign G6517 = ~G6511;
  assign G3169 = ~G6511 | ~G6518;
  assign G4935 = ~G4929;
  assign G4970 = G784;
  assign G5239 = G1014;
  assign G577 = G594 | G615;
  assign G616 = G594 | G587;
  assign G618 = G594 | G617;
  assign G620 = G594 | G619;
  assign G622 = G594 | G621;
  assign G624 = G611 | G623;
  assign G626 = G611 | G625;
  assign G628 = G611 | G627;
  assign G692 = G664 | G691;
  assign G694 = G664 | G693;
  assign G696 = G664 | G695;
  assign G698 = G664 | G697;
  assign G700 = G664 | G699;
  assign G702 = G685 | G701;
  assign G704 = G685 | G703;
  assign G706 = G685 | G705;
  assign G708 = G685 | G707;
  assign G710 = G685 | G709;
  assign G765 = ~G763 | ~G764;
  assign G4903 = ~G4897;
  assign G885 = ~G4916 | ~G4919;
  assign G1007 = ~G1005 | ~G1006;
  assign G1017 = ~G5186 | ~G5189;
  assign G5213 = ~G5207;
  assign G1363 = G141 & G1343;
  assign G1365 = G147 & G1343;
  assign G1367 = G138 & G1343;
  assign G1369 = G144 & G1343;
  assign G1371 = G135 & G1343;
  assign G1373 = G141 & G1357;
  assign G1375 = G147 & G1357;
  assign G1377 = G138 & G1357;
  assign G1379 = G144 & G1357;
  assign G1381 = G135 & G1357;
  assign G2026 = ~G2019;
  assign G2039 = ~G2032;
  assign G2046 = G103 & G2019;
  assign G2048 = G130 & G2019;
  assign G2050 = G127 & G2019;
  assign G2052 = G124 & G2019;
  assign G2054 = G100 & G2019;
  assign G2056 = G103 & G2032;
  assign G2058 = G130 & G2032;
  assign G2060 = G127 & G2032;
  assign G2062 = G124 & G2032;
  assign G2064 = G100 & G2032;
  assign G2124 = ~G2117;
  assign G2137 = ~G2130;
  assign G2144 = G115 & G2117;
  assign G2146 = G118 & G2117;
  assign G2148 = G97 & G2117;
  assign G2150 = G94 & G2117;
  assign G2152 = G121 & G2117;
  assign G2154 = G115 & G2130;
  assign G2156 = G118 & G2130;
  assign G2158 = G97 & G2130;
  assign G2160 = G94 & G2130;
  assign G2162 = G121 & G2130;
  assign G2279 = ~G2272;
  assign G2285 = G208 & G2266;
  assign G2287 = G198 & G2266;
  assign G2289 = G207 & G2266;
  assign G2291 = G206 & G2266;
  assign G2293 = G205 & G2266;
  assign G2296 = G44 & G2272;
  assign G2298 = G41 & G2272;
  assign G2300 = G29 & G2272;
  assign G2302 = G26 & G2272;
  assign G2304 = G23 & G2272;
  assign G2918 = G2899 | G2892;
  assign G2920 = G2899 | G2919;
  assign G2922 = G2899 | G2921;
  assign G2924 = G2899 | G2923;
  assign G2926 = G2899 | G2925;
  assign G2928 = G2914 | G2927;
  assign G2930 = G2914 | G2929;
  assign G2932 = G2914 | G2931;
  assign G3168 = ~G6514 | ~G6517;
  assign G6557 = ~G6551;
  assign G3211 = ~G6551 | ~G6558;
  assign G3648 = G114 & G3629;
  assign G3650 = G113 & G3629;
  assign G3652 = G111 & G3629;
  assign G3654 = G87 & G3629;
  assign G3656 = G112 & G3629;
  assign G3658 = G88 & G3642;
  assign G3660 = G1455 & G3642;
  assign G3662 = G2204 & G3642;
  assign G3665 = G3703 & G3642;
  assign G3666 = G70 & G3642;
  assign G3775 = ~G3768;
  assign G3781 = G193 & G3762;
  assign G3783 = G192 & G3762;
  assign G3785 = G191 & G3762;
  assign G3787 = G190 & G3762;
  assign G3789 = G189 & G3762;
  assign G3792 = G47 & G3768;
  assign G3794 = G35 & G3768;
  assign G3796 = G32 & G3768;
  assign G3798 = G50 & G3768;
  assign G3800 = G66 & G3768;
  assign G4101 = ~G4094;
  assign G4114 = ~G4107;
  assign G4123 = G58 & G4094;
  assign G4126 = G77 & G4094;
  assign G4129 = G78 & G4094;
  assign G4132 = G59 & G4094;
  assign G4135 = G81 & G4094;
  assign G4138 = G80 & G4107;
  assign G4141 = G79 & G4107;
  assign G4144 = G60 & G4107;
  assign G4147 = G61 & G4107;
  assign G4150 = G62 & G4107;
  assign G4451 = ~G4444;
  assign G4464 = ~G4457;
  assign G4471 = G69 & G4444;
  assign G4473 = G70 & G4444;
  assign G4475 = G74 & G4444;
  assign G4477 = G76 & G4444;
  assign G4479 = G75 & G4444;
  assign G4481 = G73 & G4457;
  assign G4483 = G53 & G4457;
  assign G4485 = G54 & G4457;
  assign G4487 = G55 & G4457;
  assign G4489 = G56 & G4457;
  assign G4666 = G82 & G4647;
  assign G4668 = G65 & G4647;
  assign G4670 = G83 & G4647;
  assign G4672 = G84 & G4647;
  assign G4674 = G85 & G4647;
  assign G4676 = G64 & G4660;
  assign G4678 = G63 & G4660;
  assign G4680 = G86 & G4660;
  assign G4682 = G109 & G4660;
  assign G4684 = G110 & G4660;
  assign G579 = G577 & G581;
  assign G629 = G616 & G581;
  assign G633 = G618 & G581;
  assign G637 = G620 & G581;
  assign G641 = G622 & G581;
  assign G645 = G624 & G601;
  assign G711 = G692 & G650;
  assign G715 = G694 & G650;
  assign G719 = G696 & G650;
  assign G723 = G698 & G650;
  assign G727 = G700 & G650;
  assign G731 = G702 & G671;
  assign G737 = G704 & G671;
  assign G745 = G706 & G671;
  assign G751 = G708 & G671;
  assign G757 = G710 & G671;
  assign G887 = ~G885 | ~G886;
  assign G1019 = ~G1017 | ~G1018;
  assign G5245 = ~G5239;
  assign G1383 = G1365 | G1366;
  assign G1387 = G1367 | G1368;
  assign G1391 = G1369 | G1370;
  assign G1395 = G1371 | G1372;
  assign G1399 = G1375 | G1376;
  assign G1406 = G1377 | G1378;
  assign G1412 = G1379 | G1380;
  assign G1418 = G1381 | G1382;
  assign G2305 = G2287 | G2288;
  assign G2308 = G2289 | G2290;
  assign G2312 = G2291 | G2292;
  assign G2316 = G2293 | G2294;
  assign G2933 = G2920 & G2886;
  assign G2938 = G2922 & G2886;
  assign G2942 = G2924 & G2886;
  assign G2946 = G2926 & G2886;
  assign G2950 = G2928 & G2905;
  assign G3170 = ~G3168 | ~G3169;
  assign G3210 = ~G6554 | ~G6557;
  assign G3667 = G3650 | G3651;
  assign G3670 = G3652 | G3653;
  assign G3673 = G3654 | G3655;
  assign G3676 = G3656 | G3657;
  assign G3679 = G3658 | G3659;
  assign G3682 = G3665 | G3635;
  assign G3686 = G3666 | G3635;
  assign G3801 = G3781 | G3782;
  assign G3804 = G3783 | G3784;
  assign G3807 = G3785 | G3786;
  assign G3810 = G3787 | G3788;
  assign G3813 = G3789 | G3790;
  assign G4525 = G2918 & G2886;
  assign G4686 = G4668 | G4669;
  assign G4689 = G4670 | G4671;
  assign G4692 = G4672 | G4673;
  assign G4695 = G4674 | G4675;
  assign G4698 = G4676 | G4677;
  assign G4701 = G4678 | G4679;
  assign G4704 = G4680 | G4681;
  assign G4707 = G4682 | G4683;
  assign G4710 = G4684 | G4685;
  assign G4976 = ~G4970;
  assign G5271 = G2932 & G2905;
  assign G5274 = G2930 & G2905;
  assign G5305 = G628 & G601;
  assign G5308 = G626 & G601;
  assign G5318 = G1373 | G1374;
  assign G6690 = G3648 | G3649;
  assign G6711 = G3662 | G3663;
  assign G6714 = G3660 | G3661;
  assign G7252 = G2285 | G2286;
  assign G7296 = G1363 | G1364;
  assign G7466 = G4666 | G4667;
  assign G907 = G765 & G784;
  assign G913 = G765 & G784;
  assign G915 = G765 & G784;
  assign G916 = G765 & G784;
  assign G1116 = G1007 & G1014;
  assign G2045 = G204 & G2026;
  assign G2047 = G203 & G2026;
  assign G2049 = G202 & G2026;
  assign G2051 = G201 & G2026;
  assign G2053 = G200 & G2026;
  assign G2055 = G235 & G2039;
  assign G2057 = G234 & G2039;
  assign G2059 = G233 & G2039;
  assign G2061 = G232 & G2039;
  assign G2063 = G231 & G2039;
  assign G2143 = G197 & G2124;
  assign G2145 = G187 & G2124;
  assign G2147 = G196 & G2124;
  assign G2149 = G195 & G2124;
  assign G2151 = G194 & G2124;
  assign G2153 = G227 & G2137;
  assign G2155 = G217 & G2137;
  assign G2157 = G226 & G2137;
  assign G2159 = G225 & G2137;
  assign G2161 = G224 & G2137;
  assign G2295 = G239 & G2279;
  assign G2297 = G229 & G2279;
  assign G2299 = G238 & G2279;
  assign G2301 = G237 & G2279;
  assign G2303 = G236 & G2279;
  assign G3212 = ~G3210 | ~G3211;
  assign G3791 = G223 & G3775;
  assign G3793 = G222 & G3775;
  assign G3795 = G221 & G3775;
  assign G3797 = G220 & G3775;
  assign G3799 = G219 & G3775;
  assign G4122 = G4121 & G4101;
  assign G4125 = G4396 & G4101;
  assign G4128 = G4402 & G4101;
  assign G4131 = G4407 & G4101;
  assign G4134 = G4412 & G4101;
  assign G4137 = G4417 & G4114;
  assign G4140 = G4422 & G4114;
  assign G4143 = G4429 & G4114;
  assign G4146 = G4434 & G4114;
  assign G4149 = G4439 & G4114;
  assign G4470 = G3700 & G4451;
  assign G4472 = G3703 & G4451;
  assign G4474 = G3707 & G4451;
  assign G4476 = G3713 & G4451;
  assign G4478 = G3719 & G4451;
  assign G4480 = G3725 & G4464;
  assign G4482 = G3731 & G4464;
  assign G4484 = G3739 & G4464;
  assign G4486 = G3745 & G4464;
  assign G4488 = G3751 & G4464;
  assign G4962 = G765;
  assign G5003 = G765;
  assign G5234 = G1007;
  assign G5242 = G1007;
  assign G5250 = ~G4525;
  assign G5284 = ~G579;
  assign G802 = G1488 & G2950;
  assign G821 = G1482 & G2946;
  assign G845 = G1477 & G2942;
  assign G868 = G1471 & G2938;
  assign G877 = G1464 & G2933;
  assign G902 = G887 & G765;
  assign G908 = G777 | G907;
  assign G914 = G887 & G765;
  assign G917 = G777 | G916;
  assign G953 = G887 & G765;
  assign G1023 = ~G1019;
  assign G1035 = G1488 & G2950;
  assign G1050 = G1482 & G2946;
  assign G1068 = G1477 & G2942;
  assign G1086 = G1471 & G2938;
  assign G1102 = G1464 & G2933;
  assign G1108 = G1019 & G1007;
  assign G1117 = G1115 | G1116;
  assign G5322 = ~G5318;
  assign G1553 = G1192 & G757;
  assign G1567 = G1186 & G751;
  assign G1584 = G2249 & G745;
  assign G1590 = G2241 & G737;
  assign G1606 = G1178 & G731;
  assign G1624 = G2232 & G1418;
  assign G1647 = G2226 & G1412;
  assign G1669 = G2220 & G1406;
  assign G1677 = G2213 & G1399;
  assign G1802 = G1192 & G757;
  assign G1816 = G1186 & G751;
  assign G1834 = G2249 & G745;
  assign G1841 = G737 & G2241;
  assign G1866 = G1178 & G731;
  assign G1880 = G2232 & G1418;
  assign G1897 = G2226 & G1412;
  assign G1914 = G2220 & G1406;
  assign G1929 = G2213 & G1399;
  assign G2065 = G2045 | G2046;
  assign G2069 = G2047 | G2048;
  assign G2073 = G2049 | G2050;
  assign G2077 = G2051 | G2052;
  assign G2081 = G2053 | G2054;
  assign G2085 = G2055 | G2056;
  assign G2091 = G2057 | G2058;
  assign G2099 = G2059 | G2060;
  assign G2105 = G2061 | G2062;
  assign G2111 = G2063 | G2064;
  assign G2163 = G2145 | G2146;
  assign G2167 = G2147 | G2148;
  assign G2171 = G2149 | G2150;
  assign G2175 = G2151 | G2152;
  assign G2179 = G2155 | G2156;
  assign G2186 = G2157 | G2158;
  assign G2192 = G2159 | G2160;
  assign G2198 = G2161 | G2162;
  assign G2320 = G2297 | G2298;
  assign G2323 = G2299 | G2300;
  assign G2329 = G2301 | G2302;
  assign G2335 = G2303 | G2304;
  assign G2962 = G4710 & G727;
  assign G2970 = G4707 & G723;
  assign G2977 = G4704 & G719;
  assign G2979 = G4701 & G715;
  assign G2989 = G4698 & G711;
  assign G2998 = G4695 & G1395;
  assign G3006 = G4692 & G1391;
  assign G3013 = G4689 & G1387;
  assign G3015 = G4686 & G1383;
  assign G3183 = G3679 & G645;
  assign G3192 = G3676 & G641;
  assign G3200 = G3673 & G637;
  assign G3207 = G3670 & G633;
  assign G3209 = G3667 & G629;
  assign G3216 = G3212 & G3170;
  assign G3222 = G3170 & G3173;
  assign G6694 = ~G6690;
  assign G3695 = G1535 & G2305;
  assign G3816 = G3791 | G3792;
  assign G3821 = G3793 | G3794;
  assign G3828 = G3795 | G3796;
  assign G3833 = G3797 | G3798;
  assign G3838 = G3799 | G3800;
  assign G4151 = G4125 | G4126;
  assign G4154 = G4128 | G4129;
  assign G4157 = G4131 | G4132;
  assign G4160 = G4134 | G4135;
  assign G4163 = G4137 | G4138;
  assign G4166 = G4140 | G4141;
  assign G4169 = G4143 | G4144;
  assign G4172 = G4146 | G4147;
  assign G4175 = G4149 | G4150;
  assign G7256 = ~G7252;
  assign G7300 = ~G7296;
  assign G4490 = G4474 | G4475;
  assign G4493 = G4476 | G4477;
  assign G4496 = G4478 | G4479;
  assign G4499 = G4480 | G4481;
  assign G4502 = G4482 | G4483;
  assign G4505 = G4484 | G4485;
  assign G4508 = G4486 | G4487;
  assign G4511 = G4488 | G4489;
  assign G7470 = ~G7466;
  assign G4884 = G2950;
  assign G4892 = G2946;
  assign G4900 = G2942;
  assign G4908 = G2938;
  assign G4924 = G2933;
  assign G4952 = G887;
  assign G4983 = ~G777 & ~G915;
  assign G4993 = G887;
  assign G5011 = ~G1464 & ~G2933;
  assign G5194 = G2950;
  assign G5202 = G2946;
  assign G5210 = G2942;
  assign G5218 = G2938;
  assign G5226 = G2933;
  assign G5247 = G2933;
  assign G5255 = G2942;
  assign G5258 = G2938;
  assign G5263 = G2950;
  assign G5266 = G2946;
  assign G5277 = ~G5271;
  assign G5278 = ~G5274;
  assign G5281 = G629;
  assign G5289 = G637;
  assign G5292 = G633;
  assign G5297 = G645;
  assign G5300 = G641;
  assign G5311 = ~G5305;
  assign G5312 = ~G5308;
  assign G5315 = G1399;
  assign G5323 = G1412;
  assign G5326 = G1406;
  assign G5331 = G731;
  assign G5334 = G1418;
  assign G5339 = G745;
  assign G5342 = G737;
  assign G5349 = G757;
  assign G5352 = G751;
  assign G5396 = G757;
  assign G5404 = G751;
  assign G5412 = G745;
  assign G5420 = G731;
  assign G5428 = G1418;
  assign G5436 = G1412;
  assign G5444 = G1406;
  assign G5452 = G737;
  assign G5460 = G1399;
  assign G5465 = ~G2241 & ~G737;
  assign G5581 = ~G2213 & ~G1399;
  assign G5748 = G757;
  assign G5756 = G751;
  assign G5764 = G745;
  assign G5772 = G737;
  assign G5780 = G731;
  assign G5788 = G1418;
  assign G5796 = G1412;
  assign G5804 = G1406;
  assign G5812 = G1399;
  assign G5849 = ~G737 & ~G2241;
  assign G5929 = G3682;
  assign G6049 = G3682;
  assign G6367 = G4710;
  assign G6370 = G727;
  assign G6375 = G4707;
  assign G6378 = G723;
  assign G6383 = G4704;
  assign G6386 = G719;
  assign G6391 = G4698;
  assign G6394 = G711;
  assign G6399 = G4695;
  assign G6402 = G1395;
  assign G6407 = G4692;
  assign G6410 = G1391;
  assign G6415 = G4689;
  assign G6418 = G1387;
  assign G6423 = G4701;
  assign G6426 = G715;
  assign G6431 = G4686;
  assign G6434 = G1383;
  assign G6442 = G3813;
  assign G6450 = G3810;
  assign G6458 = G3807;
  assign G6466 = G3801;
  assign G6498 = G3804;
  assign G6519 = G3679;
  assign G6522 = G645;
  assign G6527 = G3676;
  assign G6530 = G641;
  assign G6535 = G3673;
  assign G6538 = G637;
  assign G6543 = G3670;
  assign G6546 = G633;
  assign G6559 = G3667;
  assign G6562 = G629;
  assign G6687 = G3667;
  assign G6695 = G3673;
  assign G6698 = G3670;
  assign G6703 = G3679;
  assign G6706 = G3676;
  assign G6717 = ~G6711;
  assign G6718 = ~G6714;
  assign G6724 = G2153 | G2154;
  assign G6768 = G2295 | G2296;
  assign G7208 = G2143 | G2144;
  assign G7221 = G3801;
  assign G7229 = G3807;
  assign G7232 = G3804;
  assign G7239 = G3813;
  assign G7242 = G3810;
  assign G7249 = G2305;
  assign G7257 = G2312;
  assign G7260 = G2308;
  assign G7268 = G2316;
  assign G7293 = G1383;
  assign G7301 = G1391;
  assign G7304 = G1387;
  assign G7309 = G711;
  assign G7312 = G1395;
  assign G7317 = G719;
  assign G7320 = G715;
  assign G7327 = G727;
  assign G7330 = G723;
  assign G7396 = G2316;
  assign G7404 = G2312;
  assign G7412 = G2308;
  assign G7425 = G3686;
  assign G7463 = G4686;
  assign G7471 = G4692;
  assign G7474 = G4689;
  assign G7479 = G4698;
  assign G7482 = G4695;
  assign G7487 = G4704;
  assign G7490 = G4701;
  assign G7497 = G4710;
  assign G7500 = G4707;
  assign G7507 = G4472 | G4473;
  assign G7510 = G4470 | G4471;
  assign G7554 = G4122 | G4123;
  assign G1152 = ~G5234 | ~G5237;
  assign G5238 = ~G5234;
  assign G1156 = ~G5242 | ~G5245;
  assign G5246 = ~G5242;
  assign G5254 = ~G5250;
  assign G5288 = ~G5284;
  assign G3223 = G3221 | G3222;
  assign G4942 = G914 | G777 | G913;
  assign G4966 = ~G4962;
  assign G5007 = ~G5003;
  assign G5279 = ~G5274 | ~G5277;
  assign G5280 = ~G5271 | ~G5278;
  assign G5313 = ~G5308 | ~G5311;
  assign G5314 = ~G5305 | ~G5312;
  assign G6719 = ~G6714 | ~G6717;
  assign G6720 = ~G6711 | ~G6718;
  assign G790 = ~G4884 | ~G4887;
  assign G4888 = ~G4884;
  assign G803 = ~G4892 | ~G4895;
  assign G4896 = ~G4892;
  assign G825 = ~G4900 | ~G4903;
  assign G4904 = ~G4900;
  assign G851 = ~G4908 | ~G4911;
  assign G4912 = ~G4908;
  assign G893 = ~G4924 | ~G4927;
  assign G4928 = ~G4924;
  assign G906 = ~G902;
  assign G912 = ~G908;
  assign G1024 = ~G5194 | ~G5197;
  assign G5198 = ~G5194;
  assign G1036 = ~G5202 | ~G5205;
  assign G5206 = ~G5202;
  assign G1053 = ~G5210 | ~G5213;
  assign G5214 = ~G5210;
  assign G1072 = ~G5218 | ~G5221;
  assign G5222 = ~G5218;
  assign G1091 = ~G5226 | ~G5229;
  assign G5230 = ~G5226;
  assign G1112 = ~G1108;
  assign G1121 = ~G1117;
  assign G1153 = ~G5231 | ~G5238;
  assign G1157 = ~G5239 | ~G5246;
  assign G5253 = ~G5247;
  assign G1216 = ~G5247 | ~G5254;
  assign G5261 = ~G5255;
  assign G5262 = ~G5258;
  assign G5269 = ~G5263;
  assign G5270 = ~G5266;
  assign G5287 = ~G5281;
  assign G1239 = ~G5281 | ~G5288;
  assign G5295 = ~G5289;
  assign G5296 = ~G5292;
  assign G5303 = ~G5297;
  assign G5304 = ~G5300;
  assign G5321 = ~G5315;
  assign G1262 = ~G5315 | ~G5322;
  assign G5329 = ~G5323;
  assign G5330 = ~G5326;
  assign G5337 = ~G5331;
  assign G5338 = ~G5334;
  assign G1544 = ~G5396 | ~G5399;
  assign G5400 = ~G5396;
  assign G1554 = ~G5404 | ~G5407;
  assign G5408 = ~G5404;
  assign G1571 = ~G5412 | ~G5415;
  assign G5416 = ~G5412;
  assign G1596 = ~G5420 | ~G5423;
  assign G5424 = ~G5420;
  assign G1607 = ~G5428 | ~G5431;
  assign G5432 = ~G5428;
  assign G1628 = ~G5436 | ~G5439;
  assign G5440 = ~G5436;
  assign G1653 = ~G5444 | ~G5447;
  assign G5448 = ~G5444;
  assign G1685 = ~G5452 | ~G5455;
  assign G5456 = ~G5452;
  assign G1693 = ~G5460 | ~G5463;
  assign G5464 = ~G5460;
  assign G1793 = ~G5748 | ~G5751;
  assign G5752 = ~G5748;
  assign G1803 = ~G5756 | ~G5759;
  assign G5760 = ~G5756;
  assign G1820 = ~G5764 | ~G5767;
  assign G5768 = ~G5764;
  assign G1848 = ~G5772 | ~G5775;
  assign G5776 = ~G5772;
  assign G1857 = ~G5780 | ~G5783;
  assign G5784 = ~G5780;
  assign G1867 = ~G5788 | ~G5791;
  assign G5792 = ~G5788;
  assign G1883 = ~G5796 | ~G5799;
  assign G5800 = ~G5796;
  assign G1901 = ~G5804 | ~G5807;
  assign G5808 = ~G5804;
  assign G1919 = ~G5812 | ~G5815;
  assign G5816 = ~G5812;
  assign G5855 = ~G5849;
  assign G2351 = G3751 & G2111;
  assign G2366 = G3745 & G2105;
  assign G2384 = G3739 & G2099;
  assign G2391 = G2091 & G3731;
  assign G2417 = G3725 & G2085;
  assign G2431 = G3719 & G2335;
  assign G2448 = G3713 & G2329;
  assign G2465 = G3707 & G2323;
  assign G5935 = ~G5929;
  assign G2597 = G3751 & G2111;
  assign G2612 = G3745 & G2105;
  assign G2629 = G3739 & G2099;
  assign G2635 = G3731 & G2091;
  assign G2652 = G3725 & G2085;
  assign G2670 = G3719 & G2335;
  assign G2693 = G3713 & G2329;
  assign G2715 = G3707 & G2323;
  assign G6055 = ~G6049;
  assign G6373 = ~G6367;
  assign G6374 = ~G6370;
  assign G6381 = ~G6375;
  assign G6382 = ~G6378;
  assign G6389 = ~G6383;
  assign G6390 = ~G6386;
  assign G6397 = ~G6391;
  assign G6398 = ~G6394;
  assign G6405 = ~G6399;
  assign G6406 = ~G6402;
  assign G6413 = ~G6407;
  assign G6414 = ~G6410;
  assign G6421 = ~G6415;
  assign G6422 = ~G6418;
  assign G6429 = ~G6423;
  assign G6430 = ~G6426;
  assign G6437 = ~G6431;
  assign G6438 = ~G6434;
  assign G6446 = ~G6442;
  assign G3059 = G4175 & G3813;
  assign G6454 = ~G6450;
  assign G3068 = G4172 & G3810;
  assign G6462 = ~G6458;
  assign G3076 = G4169 & G3807;
  assign G3079 = G4166 & G3804;
  assign G6470 = ~G6466;
  assign G3090 = G4163 & G3801;
  assign G3099 = G4160 & G2175;
  assign G3107 = G4157 & G2171;
  assign G3114 = G4154 & G2167;
  assign G3116 = G4151 & G2163;
  assign G6502 = ~G6498;
  assign G6525 = ~G6519;
  assign G6526 = ~G6522;
  assign G6533 = ~G6527;
  assign G6534 = ~G6530;
  assign G6541 = ~G6535;
  assign G6542 = ~G6538;
  assign G6549 = ~G6543;
  assign G6550 = ~G6546;
  assign G6565 = ~G6559;
  assign G6566 = ~G6562;
  assign G3220 = ~G3216;
  assign G3292 = G4439 & G3838;
  assign G3308 = G4434 & G3833;
  assign G3327 = G4429 & G3828;
  assign G3335 = G3821 & G4422;
  assign G3362 = G4417 & G3816;
  assign G3376 = G4412 & G2198;
  assign G3393 = G4407 & G2192;
  assign G3410 = G4402 & G2186;
  assign G3425 = G4396 & G2179;
  assign G6693 = ~G6687;
  assign G3503 = ~G6687 | ~G6694;
  assign G6701 = ~G6695;
  assign G6702 = ~G6698;
  assign G6709 = ~G6703;
  assign G6710 = ~G6706;
  assign G6728 = ~G6724;
  assign G6772 = ~G6768;
  assign G3853 = G4439 & G3838;
  assign G3868 = G4434 & G3833;
  assign G3885 = G4429 & G3828;
  assign G3891 = G4422 & G3821;
  assign G3908 = G4417 & G3816;
  assign G3926 = G4412 & G2198;
  assign G3949 = G4407 & G2192;
  assign G3971 = G4402 & G2186;
  assign G3979 = G4396 & G2179;
  assign G7212 = ~G7208;
  assign G7227 = ~G7221;
  assign G7255 = ~G7249;
  assign G4202 = ~G7249 | ~G7256;
  assign G7263 = ~G7257;
  assign G7264 = ~G7260;
  assign G7272 = ~G7268;
  assign G7299 = ~G7293;
  assign G4225 = ~G7293 | ~G7300;
  assign G7307 = ~G7301;
  assign G7308 = ~G7304;
  assign G7315 = ~G7309;
  assign G7316 = ~G7312;
  assign G4297 = G4511 & G2081;
  assign G4305 = G4508 & G2077;
  assign G4312 = G4505 & G2073;
  assign G4314 = G4502 & G2069;
  assign G4324 = G4499 & G2065;
  assign G7400 = ~G7396;
  assign G4333 = G4496 & G2316;
  assign G7408 = ~G7404;
  assign G4341 = G4493 & G2312;
  assign G7416 = ~G7412;
  assign G4348 = G4490 & G2308;
  assign G4349 = G3686 & G3695;
  assign G7431 = ~G7425;
  assign G4389 = G2320 & G1535;
  assign G7469 = ~G7463;
  assign G4530 = ~G7463 | ~G7470;
  assign G7477 = ~G7471;
  assign G7478 = ~G7474;
  assign G7485 = ~G7479;
  assign G7486 = ~G7482;
  assign G7513 = ~G7507;
  assign G7514 = ~G7510;
  assign G7558 = ~G7554;
  assign G4932 = G917 | G953;
  assign G4956 = ~G4952;
  assign G4973 = ~G917;
  assign G4987 = ~G4983;
  assign G4997 = ~G4993;
  assign G5017 = ~G5011;
  assign G5099 = G877;
  assign G5345 = ~G5339;
  assign G5346 = ~G5342;
  assign G5355 = ~G5349;
  assign G5356 = ~G5352;
  assign G5372 = ~G5279 | ~G5280;
  assign G5380 = ~G5313 | ~G5314;
  assign G5471 = ~G5465;
  assign G5523 = G1590;
  assign G5587 = ~G5581;
  assign G5669 = G1677;
  assign G5857 = G1841;
  assign G5868 = G2111;
  assign G5876 = G2105;
  assign G5884 = G2099;
  assign G5892 = G2091;
  assign G5900 = G2085;
  assign G5908 = G2335;
  assign G5916 = G2329;
  assign G5924 = G2323;
  assign G5969 = ~G2091 & ~G3731;
  assign G5988 = G2111;
  assign G5996 = G2105;
  assign G6004 = G2099;
  assign G6012 = G2085;
  assign G6020 = G2335;
  assign G6028 = G2329;
  assign G6036 = G2323;
  assign G6044 = G2091;
  assign G6057 = ~G3731 & ~G2091;
  assign G6439 = G4175;
  assign G6447 = G4172;
  assign G6455 = G4169;
  assign G6463 = G4163;
  assign G6471 = G4160;
  assign G6474 = G2175;
  assign G6479 = G4157;
  assign G6482 = G2171;
  assign G6487 = G4154;
  assign G6490 = G2167;
  assign G6495 = G4166;
  assign G6503 = G4151;
  assign G6506 = G2163;
  assign G6570 = G3838;
  assign G6578 = G3833;
  assign G6586 = G3828;
  assign G6594 = G3821;
  assign G6602 = G3816;
  assign G6610 = G2198;
  assign G6618 = G2192;
  assign G6626 = G2186;
  assign G6634 = G2179;
  assign G6671 = ~G3821 & ~G4422;
  assign G6721 = G2179;
  assign G6729 = G2192;
  assign G6732 = G2186;
  assign G6737 = G3816;
  assign G6740 = G2198;
  assign G6745 = G3828;
  assign G6748 = G3821;
  assign G6755 = G3838;
  assign G6758 = G3833;
  assign G6765 = G2320;
  assign G6773 = G2329;
  assign G6776 = G2323;
  assign G6781 = G2085;
  assign G6784 = G2335;
  assign G6789 = G2099;
  assign G6792 = G2091;
  assign G6799 = G2111;
  assign G6802 = G2105;
  assign G6832 = ~G6719 | ~G6720;
  assign G6856 = G3838;
  assign G6864 = G3833;
  assign G6872 = G3828;
  assign G6880 = G3816;
  assign G6888 = G2198;
  assign G6896 = G2192;
  assign G6904 = G2186;
  assign G6912 = G3821;
  assign G6920 = G2179;
  assign G6925 = ~G4422 & ~G3821;
  assign G7041 = ~G4396 & ~G2179;
  assign G7205 = G2163;
  assign G7213 = G2171;
  assign G7216 = G2167;
  assign G7224 = G2175;
  assign G7235 = ~G7229;
  assign G7236 = ~G7232;
  assign G7245 = ~G7239;
  assign G7246 = ~G7242;
  assign G7265 = G2065;
  assign G7273 = G2073;
  assign G7276 = G2069;
  assign G7283 = G2081;
  assign G7286 = G2077;
  assign G7323 = ~G7317;
  assign G7324 = ~G7320;
  assign G7333 = ~G7327;
  assign G7334 = ~G7330;
  assign G7361 = G4511;
  assign G7364 = G2081;
  assign G7369 = G4508;
  assign G7372 = G2077;
  assign G7377 = G4505;
  assign G7380 = G2073;
  assign G7385 = G4499;
  assign G7388 = G2065;
  assign G7393 = G4496;
  assign G7401 = G4493;
  assign G7409 = G4490;
  assign G7417 = G4502;
  assign G7420 = G2069;
  assign G7428 = G3695;
  assign G7493 = ~G7487;
  assign G7494 = ~G7490;
  assign G7503 = ~G7497;
  assign G7504 = ~G7500;
  assign G7515 = G4493;
  assign G7518 = G4490;
  assign G7523 = G4499;
  assign G7526 = G4496;
  assign G7531 = G4505;
  assign G7534 = G4502;
  assign G7541 = G4511;
  assign G7544 = G4508;
  assign G7551 = G4151;
  assign G7559 = G4157;
  assign G7562 = G4154;
  assign G7567 = G4163;
  assign G7570 = G4160;
  assign G7575 = G4169;
  assign G7578 = G4166;
  assign G7585 = G4175;
  assign G7588 = G4172;
  assign G1176 = ~G1121 | ~G1112;
  assign G957 = ~G912 | ~G906;
  assign G791 = ~G4881 | ~G4888;
  assign G804 = ~G4889 | ~G4896;
  assign G826 = ~G4897 | ~G4904;
  assign G852 = ~G4905 | ~G4912;
  assign G894 = ~G4921 | ~G4928;
  assign G1025 = ~G5191 | ~G5198;
  assign G1037 = ~G5199 | ~G5206;
  assign G1054 = ~G5207 | ~G5214;
  assign G1073 = ~G5215 | ~G5222;
  assign G1092 = ~G5223 | ~G5230;
  assign G1154 = ~G1152 | ~G1153;
  assign G1158 = ~G1156 | ~G1157;
  assign G1215 = ~G5250 | ~G5253;
  assign G1224 = ~G5258 | ~G5261;
  assign G1225 = ~G5255 | ~G5262;
  assign G1233 = ~G5266 | ~G5269;
  assign G1234 = ~G5263 | ~G5270;
  assign G1238 = ~G5284 | ~G5287;
  assign G1247 = ~G5292 | ~G5295;
  assign G1248 = ~G5289 | ~G5296;
  assign G1256 = ~G5300 | ~G5303;
  assign G1257 = ~G5297 | ~G5304;
  assign G1261 = ~G5318 | ~G5321;
  assign G1270 = ~G5326 | ~G5329;
  assign G1271 = ~G5323 | ~G5330;
  assign G1279 = ~G5334 | ~G5337;
  assign G1280 = ~G5331 | ~G5338;
  assign G1545 = ~G5393 | ~G5400;
  assign G1555 = ~G5401 | ~G5408;
  assign G1572 = ~G5409 | ~G5416;
  assign G1597 = ~G5417 | ~G5424;
  assign G1608 = ~G5425 | ~G5432;
  assign G1629 = ~G5433 | ~G5440;
  assign G1654 = ~G5441 | ~G5448;
  assign G1686 = ~G5449 | ~G5456;
  assign G1694 = ~G5457 | ~G5464;
  assign G1794 = ~G5745 | ~G5752;
  assign G1804 = ~G5753 | ~G5760;
  assign G1821 = ~G5761 | ~G5768;
  assign G1849 = ~G5769 | ~G5776;
  assign G1858 = ~G5777 | ~G5784;
  assign G1868 = ~G5785 | ~G5792;
  assign G1884 = ~G5793 | ~G5800;
  assign G1902 = ~G5801 | ~G5808;
  assign G1920 = ~G5809 | ~G5816;
  assign G2954 = ~G6370 | ~G6373;
  assign G2955 = ~G6367 | ~G6374;
  assign G2963 = ~G6378 | ~G6381;
  assign G2964 = ~G6375 | ~G6382;
  assign G2971 = ~G6386 | ~G6389;
  assign G2972 = ~G6383 | ~G6390;
  assign G2980 = ~G6394 | ~G6397;
  assign G2981 = ~G6391 | ~G6398;
  assign G2990 = ~G6402 | ~G6405;
  assign G2991 = ~G6399 | ~G6406;
  assign G2999 = ~G6410 | ~G6413;
  assign G3000 = ~G6407 | ~G6414;
  assign G3007 = ~G6418 | ~G6421;
  assign G3008 = ~G6415 | ~G6422;
  assign G3016 = ~G6426 | ~G6429;
  assign G3017 = ~G6423 | ~G6430;
  assign G3019 = ~G6434 | ~G6437;
  assign G3020 = ~G6431 | ~G6438;
  assign G3174 = ~G6522 | ~G6525;
  assign G3175 = ~G6519 | ~G6526;
  assign G3184 = ~G6530 | ~G6533;
  assign G3185 = ~G6527 | ~G6534;
  assign G3193 = ~G6538 | ~G6541;
  assign G3194 = ~G6535 | ~G6542;
  assign G3201 = ~G6546 | ~G6549;
  assign G3202 = ~G6543 | ~G6550;
  assign G3213 = ~G6562 | ~G6565;
  assign G3214 = ~G6559 | ~G6566;
  assign G3227 = ~G3223;
  assign G3502 = ~G6690 | ~G6693;
  assign G3511 = ~G6698 | ~G6701;
  assign G3512 = ~G6695 | ~G6702;
  assign G3520 = ~G6706 | ~G6709;
  assign G3521 = ~G6703 | ~G6710;
  assign G4201 = ~G7252 | ~G7255;
  assign G4210 = ~G7260 | ~G7263;
  assign G4211 = ~G7257 | ~G7264;
  assign G4224 = ~G7296 | ~G7299;
  assign G4233 = ~G7304 | ~G7307;
  assign G4234 = ~G7301 | ~G7308;
  assign G4242 = ~G7312 | ~G7315;
  assign G4243 = ~G7309 | ~G7316;
  assign G4529 = ~G7466 | ~G7469;
  assign G4538 = ~G7474 | ~G7477;
  assign G4539 = ~G7471 | ~G7478;
  assign G4547 = ~G7482 | ~G7485;
  assign G4548 = ~G7479 | ~G7486;
  assign G4552 = ~G7510 | ~G7513;
  assign G4553 = ~G7507 | ~G7514;
  assign G4946 = ~G4942;
  assign G5347 = ~G5342 | ~G5345;
  assign G5348 = ~G5339 | ~G5346;
  assign G5357 = ~G5352 | ~G5355;
  assign G5358 = ~G5349 | ~G5356;
  assign G7237 = ~G7232 | ~G7235;
  assign G7238 = ~G7229 | ~G7236;
  assign G7247 = ~G7242 | ~G7245;
  assign G7248 = ~G7239 | ~G7246;
  assign G7325 = ~G7320 | ~G7323;
  assign G7326 = ~G7317 | ~G7324;
  assign G7335 = ~G7330 | ~G7333;
  assign G7336 = ~G7327 | ~G7334;
  assign G7495 = ~G7490 | ~G7493;
  assign G7496 = ~G7487 | ~G7494;
  assign G7505 = ~G7500 | ~G7503;
  assign G7506 = ~G7497 | ~G7504;
  assign G3244 = ~G3227 | ~G3220;
  assign G792 = ~G790 | ~G791;
  assign G805 = ~G803 | ~G804;
  assign G827 = ~G825 | ~G826;
  assign G853 = ~G851 | ~G852;
  assign G895 = ~G893 | ~G894;
  assign G1026 = ~G1024 | ~G1025;
  assign G1038 = ~G1036 | ~G1037;
  assign G1055 = ~G1053 | ~G1054;
  assign G1074 = ~G1072 | ~G1073;
  assign G1093 = ~G1091 | ~G1092;
  assign G1155 = ~G1154;
  assign G1217 = ~G1215 | ~G1216;
  assign G1226 = ~G1224 | ~G1225;
  assign G1235 = ~G1233 | ~G1234;
  assign G1240 = ~G1238 | ~G1239;
  assign G1249 = ~G1247 | ~G1248;
  assign G1258 = ~G1256 | ~G1257;
  assign G1263 = ~G1261 | ~G1262;
  assign G1272 = ~G1270 | ~G1271;
  assign G1281 = ~G1279 | ~G1280;
  assign G5376 = ~G5372;
  assign G5384 = ~G5380;
  assign G1546 = ~G1544 | ~G1545;
  assign G1556 = ~G1554 | ~G1555;
  assign G1573 = ~G1571 | ~G1572;
  assign G1598 = ~G1596 | ~G1597;
  assign G1609 = ~G1607 | ~G1608;
  assign G1630 = ~G1628 | ~G1629;
  assign G1655 = ~G1653 | ~G1654;
  assign G1687 = ~G1685 | ~G1686;
  assign G1695 = ~G1693 | ~G1694;
  assign G1795 = ~G1793 | ~G1794;
  assign G1805 = ~G1803 | ~G1804;
  assign G1822 = ~G1820 | ~G1821;
  assign G1850 = ~G1848 | ~G1849;
  assign G1859 = ~G1857 | ~G1858;
  assign G1869 = ~G1867 | ~G1868;
  assign G1885 = ~G1883 | ~G1884;
  assign G1903 = ~G1901 | ~G1902;
  assign G1921 = ~G1919 | ~G1920;
  assign G5863 = ~G5857;
  assign G2341 = ~G5868 | ~G5871;
  assign G5872 = ~G5868;
  assign G2352 = ~G5876 | ~G5879;
  assign G5880 = ~G5876;
  assign G2370 = ~G5884 | ~G5887;
  assign G5888 = ~G5884;
  assign G2398 = ~G5892 | ~G5895;
  assign G5896 = ~G5892;
  assign G2407 = ~G5900 | ~G5903;
  assign G5904 = ~G5900;
  assign G2418 = ~G5908 | ~G5911;
  assign G5912 = ~G5908;
  assign G2434 = ~G5916 | ~G5919;
  assign G5920 = ~G5916;
  assign G2452 = ~G5924 | ~G5927;
  assign G5928 = ~G5924;
  assign G2481 = G3682 & G4389;
  assign G5975 = ~G5969;
  assign G2587 = ~G5988 | ~G5991;
  assign G5992 = ~G5988;
  assign G2598 = ~G5996 | ~G5999;
  assign G6000 = ~G5996;
  assign G2616 = ~G6004 | ~G6007;
  assign G6008 = ~G6004;
  assign G2641 = ~G6012 | ~G6015;
  assign G6016 = ~G6012;
  assign G2653 = ~G6020 | ~G6023;
  assign G6024 = ~G6020;
  assign G2674 = ~G6028 | ~G6031;
  assign G6032 = ~G6028;
  assign G2699 = ~G6036 | ~G6039;
  assign G6040 = ~G6036;
  assign G2724 = G3682 & G4389;
  assign G2732 = ~G6044 | ~G6047;
  assign G6048 = ~G6044;
  assign G2956 = ~G2954 | ~G2955;
  assign G2965 = ~G2963 | ~G2964;
  assign G2973 = ~G2971 | ~G2972;
  assign G2982 = ~G2980 | ~G2981;
  assign G2992 = ~G2990 | ~G2991;
  assign G3001 = ~G2999 | ~G3000;
  assign G3009 = ~G3007 | ~G3008;
  assign G3018 = ~G3016 | ~G3017;
  assign G3021 = ~G3019 | ~G3020;
  assign G6445 = ~G6439;
  assign G3051 = ~G6439 | ~G6446;
  assign G6453 = ~G6447;
  assign G3061 = ~G6447 | ~G6454;
  assign G6461 = ~G6455;
  assign G3070 = ~G6455 | ~G6462;
  assign G6469 = ~G6463;
  assign G3081 = ~G6463 | ~G6470;
  assign G6477 = ~G6471;
  assign G6478 = ~G6474;
  assign G6485 = ~G6479;
  assign G6486 = ~G6482;
  assign G6493 = ~G6487;
  assign G6494 = ~G6490;
  assign G6501 = ~G6495;
  assign G3118 = ~G6495 | ~G6502;
  assign G6509 = ~G6503;
  assign G6510 = ~G6506;
  assign G3176 = ~G3174 | ~G3175;
  assign G3186 = ~G3184 | ~G3185;
  assign G3195 = ~G3193 | ~G3194;
  assign G3203 = ~G3201 | ~G3202;
  assign G3215 = ~G3213 | ~G3214;
  assign G3281 = ~G6570 | ~G6573;
  assign G6574 = ~G6570;
  assign G3293 = ~G6578 | ~G6581;
  assign G6582 = ~G6578;
  assign G3312 = ~G6586 | ~G6589;
  assign G6590 = ~G6586;
  assign G3342 = ~G6594 | ~G6597;
  assign G6598 = ~G6594;
  assign G3351 = ~G6602 | ~G6605;
  assign G6606 = ~G6602;
  assign G3363 = ~G6610 | ~G6613;
  assign G6614 = ~G6610;
  assign G3379 = ~G6618 | ~G6621;
  assign G6622 = ~G6618;
  assign G3397 = ~G6626 | ~G6629;
  assign G6630 = ~G6626;
  assign G3415 = ~G6634 | ~G6637;
  assign G6638 = ~G6634;
  assign G6677 = ~G6671;
  assign G3504 = ~G3502 | ~G3503;
  assign G3513 = ~G3511 | ~G3512;
  assign G3522 = ~G3520 | ~G3521;
  assign G6727 = ~G6721;
  assign G3526 = ~G6721 | ~G6728;
  assign G6735 = ~G6729;
  assign G6736 = ~G6732;
  assign G6743 = ~G6737;
  assign G6744 = ~G6740;
  assign G6771 = ~G6765;
  assign G3549 = ~G6765 | ~G6772;
  assign G6779 = ~G6773;
  assign G6780 = ~G6776;
  assign G6787 = ~G6781;
  assign G6788 = ~G6784;
  assign G6836 = ~G6832;
  assign G3843 = ~G6856 | ~G6859;
  assign G6860 = ~G6856;
  assign G3854 = ~G6864 | ~G6867;
  assign G6868 = ~G6864;
  assign G3872 = ~G6872 | ~G6875;
  assign G6876 = ~G6872;
  assign G3897 = ~G6880 | ~G6883;
  assign G6884 = ~G6880;
  assign G3909 = ~G6888 | ~G6891;
  assign G6892 = ~G6888;
  assign G3930 = ~G6896 | ~G6899;
  assign G6900 = ~G6896;
  assign G3955 = ~G6904 | ~G6907;
  assign G6908 = ~G6904;
  assign G3987 = ~G6912 | ~G6915;
  assign G6916 = ~G6912;
  assign G3995 = ~G6920 | ~G6923;
  assign G6924 = ~G6920;
  assign G7211 = ~G7205;
  assign G4179 = ~G7205 | ~G7212;
  assign G7219 = ~G7213;
  assign G7220 = ~G7216;
  assign G4196 = ~G7224 | ~G7227;
  assign G7228 = ~G7224;
  assign G4203 = ~G4201 | ~G4202;
  assign G4212 = ~G4210 | ~G4211;
  assign G7271 = ~G7265;
  assign G4220 = ~G7265 | ~G7272;
  assign G4226 = ~G4224 | ~G4225;
  assign G4235 = ~G4233 | ~G4234;
  assign G4244 = ~G4242 | ~G4243;
  assign G7367 = ~G7361;
  assign G7368 = ~G7364;
  assign G7375 = ~G7369;
  assign G7376 = ~G7372;
  assign G7383 = ~G7377;
  assign G7384 = ~G7380;
  assign G7391 = ~G7385;
  assign G7392 = ~G7388;
  assign G7399 = ~G7393;
  assign G4326 = ~G7393 | ~G7400;
  assign G7407 = ~G7401;
  assign G4335 = ~G7401 | ~G7408;
  assign G7415 = ~G7409;
  assign G4343 = ~G7409 | ~G7416;
  assign G7423 = ~G7417;
  assign G7424 = ~G7420;
  assign G4353 = ~G7428 | ~G7431;
  assign G7432 = ~G7428;
  assign G4531 = ~G4529 | ~G4530;
  assign G4540 = ~G4538 | ~G4539;
  assign G4549 = ~G4547 | ~G4548;
  assign G4554 = ~G4552 | ~G4553;
  assign G7521 = ~G7515;
  assign G7522 = ~G7518;
  assign G7529 = ~G7523;
  assign G7530 = ~G7526;
  assign G7557 = ~G7551;
  assign G4576 = ~G7551 | ~G7558;
  assign G7565 = ~G7559;
  assign G7566 = ~G7562;
  assign G7573 = ~G7567;
  assign G7574 = ~G7570;
  assign G4936 = ~G4932;
  assign G4937 = ~G4932 | ~G4935;
  assign G4977 = ~G4973;
  assign G4978 = ~G4973 | ~G4976;
  assign G5105 = ~G5099;
  assign G5359 = ~G5357 | ~G5358;
  assign G5362 = ~G5347 | ~G5348;
  assign G5529 = ~G5523;
  assign G5675 = ~G5669;
  assign G5932 = G4389;
  assign G5977 = G2391;
  assign G6052 = G4389;
  assign G6063 = ~G6057;
  assign G6115 = G2635;
  assign G6173 = ~G3682 & ~G4389;
  assign G6679 = G3335;
  assign G6751 = ~G6745;
  assign G6752 = ~G6748;
  assign G6761 = ~G6755;
  assign G6762 = ~G6758;
  assign G6795 = ~G6789;
  assign G6796 = ~G6792;
  assign G6805 = ~G6799;
  assign G6806 = ~G6802;
  assign G6931 = ~G6925;
  assign G6983 = G3891;
  assign G7047 = ~G7041;
  assign G7129 = G3979;
  assign G7279 = ~G7273;
  assign G7280 = ~G7276;
  assign G7289 = ~G7283;
  assign G7290 = ~G7286;
  assign G7337 = ~G7247 | ~G7248;
  assign G7340 = ~G7237 | ~G7238;
  assign G7353 = ~G7335 | ~G7336;
  assign G7356 = ~G7325 | ~G7326;
  assign G7537 = ~G7531;
  assign G7538 = ~G7534;
  assign G7547 = ~G7541;
  assign G7548 = ~G7544;
  assign G7581 = ~G7575;
  assign G7582 = ~G7578;
  assign G7591 = ~G7585;
  assign G7592 = ~G7588;
  assign G7595 = ~G7505 | ~G7506;
  assign G7598 = ~G7495 | ~G7496;
  assign G2342 = ~G5865 | ~G5872;
  assign G2353 = ~G5873 | ~G5880;
  assign G2371 = ~G5881 | ~G5888;
  assign G2399 = ~G5889 | ~G5896;
  assign G2408 = ~G5897 | ~G5904;
  assign G2419 = ~G5905 | ~G5912;
  assign G2435 = ~G5913 | ~G5920;
  assign G2453 = ~G5921 | ~G5928;
  assign G2588 = ~G5985 | ~G5992;
  assign G2599 = ~G5993 | ~G6000;
  assign G2617 = ~G6001 | ~G6008;
  assign G2642 = ~G6009 | ~G6016;
  assign G2654 = ~G6017 | ~G6024;
  assign G2675 = ~G6025 | ~G6032;
  assign G2700 = ~G6033 | ~G6040;
  assign G2733 = ~G6041 | ~G6048;
  assign G3050 = ~G6442 | ~G6445;
  assign G3060 = ~G6450 | ~G6453;
  assign G3069 = ~G6458 | ~G6461;
  assign G3080 = ~G6466 | ~G6469;
  assign G3091 = ~G6474 | ~G6477;
  assign G3092 = ~G6471 | ~G6478;
  assign G3100 = ~G6482 | ~G6485;
  assign G3101 = ~G6479 | ~G6486;
  assign G3108 = ~G6490 | ~G6493;
  assign G3109 = ~G6487 | ~G6494;
  assign G3117 = ~G6498 | ~G6501;
  assign G3120 = ~G6506 | ~G6509;
  assign G3121 = ~G6503 | ~G6510;
  assign G3282 = ~G6567 | ~G6574;
  assign G3294 = ~G6575 | ~G6582;
  assign G3313 = ~G6583 | ~G6590;
  assign G3343 = ~G6591 | ~G6598;
  assign G3352 = ~G6599 | ~G6606;
  assign G3364 = ~G6607 | ~G6614;
  assign G3380 = ~G6615 | ~G6622;
  assign G3398 = ~G6623 | ~G6630;
  assign G3416 = ~G6631 | ~G6638;
  assign G3525 = ~G6724 | ~G6727;
  assign G3534 = ~G6732 | ~G6735;
  assign G3535 = ~G6729 | ~G6736;
  assign G3543 = ~G6740 | ~G6743;
  assign G3544 = ~G6737 | ~G6744;
  assign G3548 = ~G6768 | ~G6771;
  assign G3557 = ~G6776 | ~G6779;
  assign G3558 = ~G6773 | ~G6780;
  assign G3566 = ~G6784 | ~G6787;
  assign G3567 = ~G6781 | ~G6788;
  assign G3844 = ~G6853 | ~G6860;
  assign G3855 = ~G6861 | ~G6868;
  assign G3873 = ~G6869 | ~G6876;
  assign G3898 = ~G6877 | ~G6884;
  assign G3910 = ~G6885 | ~G6892;
  assign G3931 = ~G6893 | ~G6900;
  assign G3956 = ~G6901 | ~G6908;
  assign G3988 = ~G6909 | ~G6916;
  assign G3996 = ~G6917 | ~G6924;
  assign G4178 = ~G7208 | ~G7211;
  assign G4187 = ~G7216 | ~G7219;
  assign G4188 = ~G7213 | ~G7220;
  assign G4197 = ~G7221 | ~G7228;
  assign G4219 = ~G7268 | ~G7271;
  assign G4289 = ~G7364 | ~G7367;
  assign G4290 = ~G7361 | ~G7368;
  assign G4298 = ~G7372 | ~G7375;
  assign G4299 = ~G7369 | ~G7376;
  assign G4306 = ~G7380 | ~G7383;
  assign G4307 = ~G7377 | ~G7384;
  assign G4315 = ~G7388 | ~G7391;
  assign G4316 = ~G7385 | ~G7392;
  assign G4325 = ~G7396 | ~G7399;
  assign G4334 = ~G7404 | ~G7407;
  assign G4342 = ~G7412 | ~G7415;
  assign G4350 = ~G7420 | ~G7423;
  assign G4351 = ~G7417 | ~G7424;
  assign G4354 = ~G7425 | ~G7432;
  assign G4561 = ~G7518 | ~G7521;
  assign G4562 = ~G7515 | ~G7522;
  assign G4570 = ~G7526 | ~G7529;
  assign G4571 = ~G7523 | ~G7530;
  assign G4575 = ~G7554 | ~G7557;
  assign G4584 = ~G7562 | ~G7565;
  assign G4585 = ~G7559 | ~G7566;
  assign G4593 = ~G7570 | ~G7573;
  assign G4594 = ~G7567 | ~G7574;
  assign G4938 = ~G4929 | ~G4936;
  assign G4979 = ~G4970 | ~G4977;
  assign G6753 = ~G6748 | ~G6751;
  assign G6754 = ~G6745 | ~G6752;
  assign G6763 = ~G6758 | ~G6761;
  assign G6764 = ~G6755 | ~G6762;
  assign G6797 = ~G6792 | ~G6795;
  assign G6798 = ~G6789 | ~G6796;
  assign G6807 = ~G6802 | ~G6805;
  assign G6808 = ~G6799 | ~G6806;
  assign G7281 = ~G7276 | ~G7279;
  assign G7282 = ~G7273 | ~G7280;
  assign G7291 = ~G7286 | ~G7289;
  assign G7292 = ~G7283 | ~G7290;
  assign G7539 = ~G7534 | ~G7537;
  assign G7540 = ~G7531 | ~G7538;
  assign G7549 = ~G7544 | ~G7547;
  assign G7550 = ~G7541 | ~G7548;
  assign G7583 = ~G7578 | ~G7581;
  assign G7584 = ~G7575 | ~G7582;
  assign G7593 = ~G7588 | ~G7591;
  assign G7594 = ~G7585 | ~G7592;
  assign G1856 = ~G1850;
  assign G920 = G792 & G805 & G827 & G895 & G853;
  assign G925 = G792 & G821;
  assign G926 = G845 & G805 & G792;
  assign G927 = G805 & G868 & G827 & G792;
  assign G928 = G805 & G877 & G792 & G853 & G827;
  assign G937 = G805 & G845;
  assign G938 = G805 & G827 & G868;
  assign G939 = G805 & G877 & G853 & G827;
  assign G940 = G853 & G805 & G895 & G827;
  assign G941 = G805 & G845;
  assign G942 = G805 & G827 & G868;
  assign G943 = G805 & G877 & G853 & G827;
  assign G944 = G827 & G868;
  assign G945 = G877 & G853 & G827;
  assign G946 = G853 & G895 & G827;
  assign G947 = G827 & G868;
  assign G948 = G877 & G853 & G827;
  assign G949 = G853 & G877;
  assign G956 = G895 & G853;
  assign G1122 = G1074 & G1026 & G1055 & G1038 & G1093;
  assign G1125 = G1026 & G1050;
  assign G1126 = G1068 & G1038 & G1026;
  assign G1127 = G1038 & G1086 & G1055 & G1026;
  assign G1128 = G1038 & G1102 & G1026 & G1074 & G1055;
  assign G1132 = G1038 & G1068;
  assign G1133 = G1038 & G1055 & G1086;
  assign G1134 = G1038 & G1102 & G1074 & G1055;
  assign G1137 = G1086 & G1055;
  assign G1138 = G1102 & G1074 & G1055;
  assign G1141 = G1074 & G1102;
  assign G1221 = ~G1217;
  assign G1230 = ~G1226;
  assign G1244 = ~G1240;
  assign G1253 = ~G1249;
  assign G1267 = ~G1263;
  assign G1276 = ~G1272;
  assign G1284 = G1235;
  assign G1288 = G1235;
  assign G1292 = G1258;
  assign G1296 = G1258;
  assign G1300 = G1281;
  assign G1304 = G1281;
  assign G1702 = G1546 & G1556 & G1687 & G1573;
  assign G1705 = G1546 & G1567;
  assign G1706 = G1584 & G1556 & G1546;
  assign G1707 = G1556 & G1590 & G1573 & G1546;
  assign G1709 = G1556 & G1584;
  assign G1710 = G1556 & G1573 & G1590;
  assign G1711 = G1556 & G1687 & G1573;
  assign G1712 = G1556 & G1584;
  assign G1713 = G1556 & G1573 & G1590;
  assign G1714 = G1573 & G1590;
  assign G1718 = G1598 & G1609 & G1630 & G1695 & G1655;
  assign G1722 = G1598 & G1624;
  assign G1723 = G1647 & G1609 & G1598;
  assign G1724 = G1609 & G1669 & G1630 & G1598;
  assign G1725 = G1609 & G1677 & G1598 & G1655 & G1630;
  assign G1733 = G1609 & G1647;
  assign G1734 = G1609 & G1630 & G1669;
  assign G1735 = G1609 & G1677 & G1655 & G1630;
  assign G1736 = G1655 & G1609 & G1695 & G1630;
  assign G1737 = G1609 & G1647;
  assign G1738 = G1609 & G1630 & G1669;
  assign G1739 = G1609 & G1677 & G1655 & G1630;
  assign G1740 = G1630 & G1669;
  assign G1741 = G1677 & G1655 & G1630;
  assign G1742 = G1655 & G1695 & G1630;
  assign G1743 = G1630 & G1669;
  assign G1744 = G1677 & G1655 & G1630;
  assign G1745 = G1655 & G1677;
  assign G1749 = G1687 & G1573;
  assign G1750 = G1695 & G1655;
  assign G1935 = G1795 & G1822 & G1805 & G1850;
  assign G1938 = G1795 & G1816;
  assign G1939 = G1834 & G1805 & G1795;
  assign G1940 = G1805 & G1841 & G1822 & G1795;
  assign G1942 = G1805 & G1834;
  assign G1943 = G1805 & G1822 & G1841;
  assign G1944 = G1805 & G1850 & G1822;
  assign G1945 = G1805 & G1834;
  assign G1946 = G1805 & G1841 & G1822;
  assign G1947 = G1822 & G1841;
  assign G1948 = G1850 & G1822;
  assign G1949 = G1822 & G1841;
  assign G1950 = G1903 & G1859 & G1885 & G1869 & G1921;
  assign G1953 = G1859 & G1880;
  assign G1954 = G1897 & G1869 & G1859;
  assign G1955 = G1869 & G1914 & G1885 & G1859;
  assign G1956 = G1869 & G1929 & G1859 & G1903 & G1885;
  assign G1960 = G1869 & G1897;
  assign G1961 = G1869 & G1885 & G1914;
  assign G1962 = G1869 & G1929 & G1903 & G1885;
  assign G1965 = G1914 & G1885;
  assign G1966 = G1929 & G1903 & G1885;
  assign G1969 = G1903 & G1929;
  assign G2343 = ~G2341 | ~G2342;
  assign G2354 = ~G2352 | ~G2353;
  assign G2372 = ~G2370 | ~G2371;
  assign G2400 = ~G2398 | ~G2399;
  assign G2409 = ~G2407 | ~G2408;
  assign G2420 = ~G2418 | ~G2419;
  assign G2436 = ~G2434 | ~G2435;
  assign G2454 = ~G2452 | ~G2453;
  assign G2470 = ~G5932 | ~G5935;
  assign G5936 = ~G5932;
  assign G5983 = ~G5977;
  assign G2589 = ~G2587 | ~G2588;
  assign G2600 = ~G2598 | ~G2599;
  assign G2618 = ~G2616 | ~G2617;
  assign G2643 = ~G2641 | ~G2642;
  assign G2655 = ~G2653 | ~G2654;
  assign G2676 = ~G2674 | ~G2675;
  assign G2701 = ~G2699 | ~G2700;
  assign G2734 = ~G2732 | ~G2733;
  assign G2740 = ~G6052 | ~G6055;
  assign G6056 = ~G6052;
  assign G3022 = G2956 & G2965 & G3018 & G2973;
  assign G3025 = G2956 & G2970;
  assign G3026 = G2977 & G2965 & G2956;
  assign G3027 = G2965 & G2979 & G2973 & G2956;
  assign G3029 = G2982 & G2992 & G3001 & G3021 & G3009;
  assign G3030 = G2982 & G2998;
  assign G3031 = G3006 & G2992 & G2982;
  assign G3032 = G2992 & G3013 & G3001 & G2982;
  assign G3033 = G2992 & G3015 & G2982 & G3009 & G3001;
  assign G3052 = ~G3050 | ~G3051;
  assign G3062 = ~G3060 | ~G3061;
  assign G3071 = ~G3069 | ~G3070;
  assign G3082 = ~G3080 | ~G3081;
  assign G3093 = ~G3091 | ~G3092;
  assign G3102 = ~G3100 | ~G3101;
  assign G3110 = ~G3108 | ~G3109;
  assign G3119 = ~G3117 | ~G3118;
  assign G3122 = ~G3120 | ~G3121;
  assign G3228 = G3176 & G3186 & G3195 & G3215 & G3203;
  assign G3231 = G3176 & G3192;
  assign G3232 = G3200 & G3186 & G3176;
  assign G3233 = G3186 & G3207 & G3195 & G3176;
  assign G3234 = G3186 & G3209 & G3176 & G3203 & G3195;
  assign G3283 = ~G3281 | ~G3282;
  assign G3295 = ~G3293 | ~G3294;
  assign G3314 = ~G3312 | ~G3313;
  assign G3344 = ~G3342 | ~G3343;
  assign G3353 = ~G3351 | ~G3352;
  assign G3365 = ~G3363 | ~G3364;
  assign G3381 = ~G3379 | ~G3380;
  assign G3399 = ~G3397 | ~G3398;
  assign G3417 = ~G3415 | ~G3416;
  assign G6685 = ~G6679;
  assign G3508 = ~G3504;
  assign G3517 = ~G3513;
  assign G3527 = ~G3525 | ~G3526;
  assign G3536 = ~G3534 | ~G3535;
  assign G3545 = ~G3543 | ~G3544;
  assign G3550 = ~G3548 | ~G3549;
  assign G3559 = ~G3557 | ~G3558;
  assign G3568 = ~G3566 | ~G3567;
  assign G3571 = G3522;
  assign G3575 = G3522;
  assign G3845 = ~G3843 | ~G3844;
  assign G3856 = ~G3854 | ~G3855;
  assign G3874 = ~G3872 | ~G3873;
  assign G3899 = ~G3897 | ~G3898;
  assign G3911 = ~G3909 | ~G3910;
  assign G3932 = ~G3930 | ~G3931;
  assign G3957 = ~G3955 | ~G3956;
  assign G3989 = ~G3987 | ~G3988;
  assign G3997 = ~G3995 | ~G3996;
  assign G4180 = ~G4178 | ~G4179;
  assign G4189 = ~G4187 | ~G4188;
  assign G4198 = ~G4196 | ~G4197;
  assign G4207 = ~G4203;
  assign G4216 = ~G4212;
  assign G4221 = ~G4219 | ~G4220;
  assign G4230 = ~G4226;
  assign G4239 = ~G4235;
  assign G4263 = G4244;
  assign G4267 = G4244;
  assign G4291 = ~G4289 | ~G4290;
  assign G4300 = ~G4298 | ~G4299;
  assign G4308 = ~G4306 | ~G4307;
  assign G4317 = ~G4315 | ~G4316;
  assign G4327 = ~G4325 | ~G4326;
  assign G4336 = ~G4334 | ~G4335;
  assign G4344 = ~G4342 | ~G4343;
  assign G4352 = ~G4350 | ~G4351;
  assign G4355 = ~G4353 | ~G4354;
  assign G4535 = ~G4531;
  assign G4544 = ~G4540;
  assign G4558 = ~G4554;
  assign G4563 = ~G4561 | ~G4562;
  assign G4572 = ~G4570 | ~G4571;
  assign G4577 = ~G4575 | ~G4576;
  assign G4586 = ~G4584 | ~G4585;
  assign G4595 = ~G4593 | ~G4594;
  assign G4598 = G4549;
  assign G4602 = G4549;
  assign G4716 = G1921;
  assign G4724 = G1859;
  assign G4732 = G1869;
  assign G4740 = G1885;
  assign G4748 = G1903;
  assign G4756 = G1093;
  assign G4764 = G1026;
  assign G4772 = G1038;
  assign G4780 = G1055;
  assign G4788 = G1074;
  assign G4939 = ~G4937 | ~G4938;
  assign G4980 = ~G4978 | ~G4979;
  assign G5044 = G895;
  assign G5054 = G853;
  assign G5064 = G792;
  assign G5074 = G827;
  assign G5084 = G805;
  assign G5094 = G805;
  assign G5132 = G895;
  assign G5142 = G853;
  assign G5152 = G792;
  assign G5162 = G827;
  assign G5365 = ~G5359;
  assign G5366 = ~G5362;
  assign G5488 = G1687;
  assign G5498 = G1573;
  assign G5508 = G1546;
  assign G5518 = G1556;
  assign G5546 = G1687;
  assign G5556 = G1573;
  assign G5566 = G1546;
  assign G5576 = G1556;
  assign G5614 = G1695;
  assign G5624 = G1655;
  assign G5634 = G1598;
  assign G5644 = G1630;
  assign G5654 = G1609;
  assign G5664 = G1609;
  assign G5702 = G1695;
  assign G5712 = G1655;
  assign G5722 = G1598;
  assign G5732 = G1630;
  assign G5820 = G1795;
  assign G5828 = G1795;
  assign G5836 = G1805;
  assign G5844 = G1805;
  assign G5852 = G1822;
  assign G5860 = G1822;
  assign G6121 = ~G6115;
  assign G6179 = ~G6173;
  assign G6261 = G2724;
  assign G7359 = ~G7353;
  assign G7360 = ~G7356;
  assign G7343 = ~G7337;
  assign G7344 = ~G7340;
  assign G6809 = ~G6763 | ~G6764;
  assign G6812 = ~G6753 | ~G6754;
  assign G6819 = ~G6807 | ~G6808;
  assign G6822 = ~G6797 | ~G6798;
  assign G6989 = ~G6983;
  assign G7135 = ~G7129;
  assign G7345 = ~G7291 | ~G7292;
  assign G7348 = ~G7281 | ~G7282;
  assign G7601 = ~G7595;
  assign G7602 = ~G7598;
  assign G7603 = ~G7549 | ~G7550;
  assign G7606 = ~G7539 | ~G7540;
  assign G7611 = ~G7593 | ~G7594;
  assign G7614 = ~G7583 | ~G7584;
  assign G929 = G928 | G927 | G926 | G802 | G925;
  assign G950 = G868 | G949;
  assign G1129 = G1128 | G1127 | G1126 | G1035 | G1125;
  assign G1708 = G1707 | G1706 | G1553 | G1705;
  assign G1715 = G1584 | G1714;
  assign G1726 = G1725 | G1724 | G1723 | G1606 | G1722;
  assign G1746 = G1669 | G1745;
  assign G1941 = G1940 | G1939 | G1802 | G1938;
  assign G1957 = G1956 | G1955 | G1954 | G1866 | G1953;
  assign G2471 = ~G5929 | ~G5936;
  assign G2741 = ~G6049 | ~G6056;
  assign G3028 = G3027 | G3026 | G2962 | G3025;
  assign G3034 = G3033 | G3032 | G3031 | G2989 | G3030;
  assign G3235 = G3234 | G3233 | G3232 | G3183 | G3231;
  assign G5014 = G946 | G945 | G845 | G944;
  assign G5034 = G940 | G939 | G938 | G821 | G937;
  assign G5102 = ~G948 & ~G845 & ~G947;
  assign G5122 = ~G943 & ~G942 & ~G821 & ~G941;
  assign G5367 = ~G5362 | ~G5365;
  assign G5368 = ~G5359 | ~G5366;
  assign G5478 = G1711 | G1710 | G1567 | G1709;
  assign G5536 = ~G1713 & ~G1567 & ~G1712;
  assign G5584 = G1742 | G1741 | G1647 | G1740;
  assign G5604 = G1736 | G1735 | G1734 | G1624 | G1733;
  assign G5672 = ~G1744 & ~G1647 & ~G1743;
  assign G5692 = ~G1739 & ~G1738 & ~G1624 & ~G1737;
  assign G5817 = G1944 | G1943 | G1816 | G1942;
  assign G5825 = ~G1946 & ~G1816 & ~G1945;
  assign G5833 = G1948 | G1834 | G1947;
  assign G5841 = ~G1834 & ~G1949;
  assign G6340 = ~G7356 | ~G7359;
  assign G6341 = ~G7353 | ~G7360;
  assign G6350 = ~G7340 | ~G7343;
  assign G6351 = ~G7337 | ~G7344;
  assign G7436 = ~G7598 | ~G7601;
  assign G7437 = ~G7595 | ~G7602;
  assign G4720 = ~G4716;
  assign G4728 = ~G4724;
  assign G4736 = ~G4732;
  assign G4744 = ~G4740;
  assign G4752 = ~G4748;
  assign G4760 = ~G4756;
  assign G4768 = ~G4764;
  assign G4776 = ~G4772;
  assign G4784 = ~G4780;
  assign G4792 = ~G4788;
  assign G3350 = ~G3344;
  assign G2406 = ~G2400;
  assign G924 = ~G920;
  assign G5088 = ~G5084;
  assign G5098 = ~G5094;
  assign G997 = G902 & G920;
  assign G1146 = G1108 & G1122;
  assign G1287 = ~G1284;
  assign G1291 = ~G1288;
  assign G1295 = ~G1292;
  assign G1299 = ~G1296;
  assign G1303 = ~G1300;
  assign G1307 = ~G1304;
  assign G1309 = G1284 & G1226 & G1217;
  assign G1312 = G1288 & G1230 & G1221;
  assign G1315 = G1292 & G1249 & G1240;
  assign G1318 = G1296 & G1253 & G1244;
  assign G1321 = G1300 & G1272 & G1263;
  assign G1324 = G1304 & G1276 & G1267;
  assign G1721 = ~G1718;
  assign G5522 = ~G5518;
  assign G5580 = ~G5576;
  assign G5658 = ~G5654;
  assign G5668 = ~G5664;
  assign G1788 = G1702 & G1718;
  assign G1974 = G1935 & G1950;
  assign G5824 = ~G5820;
  assign G5832 = ~G5828;
  assign G5840 = ~G5836;
  assign G5848 = ~G5844;
  assign G1999 = ~G5852 | ~G5855;
  assign G5856 = ~G5852;
  assign G2003 = ~G5860 | ~G5863;
  assign G5864 = ~G5860;
  assign G2472 = ~G2470 | ~G2471;
  assign G2487 = G2343 & G2372 & G2354 & G2400;
  assign G2492 = G2343 & G2366;
  assign G2493 = G2384 & G2354 & G2343;
  assign G2494 = G2354 & G2391 & G2372 & G2343;
  assign G2500 = G2354 & G2384;
  assign G2501 = G2354 & G2372 & G2391;
  assign G2502 = G2354 & G2400 & G2372;
  assign G2503 = G2354 & G2384;
  assign G2504 = G2354 & G2391 & G2372;
  assign G2505 = G2372 & G2391;
  assign G2506 = G2400 & G2372;
  assign G2507 = G2372 & G2391;
  assign G2511 = G2409 & G2431;
  assign G2512 = G2448 & G2420 & G2409;
  assign G2513 = G2420 & G2465 & G2436 & G2409;
  assign G2514 = G2420 & G2481 & G2409 & G2454 & G2436;
  assign G2518 = G2420 & G2448;
  assign G2519 = G2420 & G2436 & G2465;
  assign G2520 = G2420 & G2481 & G2454 & G2436;
  assign G2523 = G2465 & G2436;
  assign G2524 = G2481 & G2454 & G2436;
  assign G2527 = G2454 & G2481;
  assign G2742 = ~G2740 | ~G2741;
  assign G2749 = G2589 & G2600 & G2734 & G2618;
  assign G2754 = G2589 & G2612;
  assign G2755 = G2629 & G2600 & G2589;
  assign G2756 = G2600 & G2635 & G2618 & G2589;
  assign G2762 = G2600 & G2629;
  assign G2763 = G2600 & G2618 & G2635;
  assign G2764 = G2600 & G2734 & G2618;
  assign G2765 = G2600 & G2629;
  assign G2766 = G2600 & G2618 & G2635;
  assign G2767 = G2618 & G2635;
  assign G2776 = G2643 & G2670;
  assign G2777 = G2693 & G2655 & G2643;
  assign G2778 = G2655 & G2715 & G2676 & G2643;
  assign G2779 = G2655 & G2724 & G2643 & G2701 & G2676;
  assign G2788 = G2655 & G2693;
  assign G2789 = G2655 & G2676 & G2715;
  assign G2790 = G2655 & G2724 & G2701 & G2676;
  assign G2792 = G2655 & G2693;
  assign G2793 = G2655 & G2676 & G2715;
  assign G2794 = G2655 & G2724 & G2701 & G2676;
  assign G2795 = G2676 & G2715;
  assign G2796 = G2724 & G2701 & G2676;
  assign G2798 = G2676 & G2715;
  assign G2799 = G2724 & G2701 & G2676;
  assign G2800 = G2701 & G2724;
  assign G2804 = G2734 & G2618;
  assign G3035 = G3022 & G3029;
  assign G3045 = G3022 & G3034;
  assign G3123 = G3052 & G3062 & G3119 & G3071;
  assign G3128 = G3052 & G3068;
  assign G3129 = G3076 & G3062 & G3052;
  assign G3130 = G3062 & G3079 & G3071 & G3052;
  assign G3136 = G3082 & G3093 & G3102 & G3122 & G3110;
  assign G3139 = G3082 & G3099;
  assign G3140 = G3107 & G3093 & G3082;
  assign G3141 = G3093 & G3114 & G3102 & G3082;
  assign G3142 = G3093 & G3116 & G3082 & G3110 & G3102;
  assign G3249 = G3216 & G3228;
  assign G3431 = G3283 & G3314 & G3295 & G3344;
  assign G3434 = G3283 & G3308;
  assign G3435 = G3327 & G3295 & G3283;
  assign G3436 = G3295 & G3335 & G3314 & G3283;
  assign G3438 = G3295 & G3327;
  assign G3439 = G3295 & G3314 & G3335;
  assign G3440 = G3295 & G3344 & G3314;
  assign G3441 = G3295 & G3327;
  assign G3442 = G3295 & G3335 & G3314;
  assign G3443 = G3314 & G3335;
  assign G3444 = G3344 & G3314;
  assign G3445 = G3314 & G3335;
  assign G3446 = G3399 & G3353 & G3381 & G3365 & G3417;
  assign G3449 = G3353 & G3376;
  assign G3450 = G3393 & G3365 & G3353;
  assign G3451 = G3365 & G3410 & G3381 & G3353;
  assign G3452 = G3365 & G3425 & G3353 & G3399 & G3381;
  assign G3456 = G3365 & G3393;
  assign G3457 = G3365 & G3381 & G3410;
  assign G3458 = G3365 & G3425 & G3399 & G3381;
  assign G3460 = G3410 & G3381;
  assign G3461 = G3425 & G3399 & G3381;
  assign G3463 = G3399 & G3425;
  assign G3531 = ~G3527;
  assign G3540 = ~G3536;
  assign G3554 = ~G3550;
  assign G3563 = ~G3559;
  assign G3574 = ~G3571;
  assign G3578 = ~G3575;
  assign G3579 = G3545;
  assign G3583 = G3545;
  assign G3587 = G3568;
  assign G3591 = G3568;
  assign G3596 = G3571 & G3513 & G3504;
  assign G3599 = G3575 & G3517 & G3508;
  assign G4004 = G3845 & G3856 & G3989 & G3874;
  assign G4007 = G3845 & G3868;
  assign G4008 = G3885 & G3856 & G3845;
  assign G4009 = G3856 & G3891 & G3874 & G3845;
  assign G4011 = G3856 & G3885;
  assign G4012 = G3856 & G3874 & G3891;
  assign G4013 = G3856 & G3989 & G3874;
  assign G4014 = G3856 & G3885;
  assign G4015 = G3856 & G3874 & G3891;
  assign G4016 = G3874 & G3891;
  assign G4020 = G3899 & G3911 & G3932 & G3997 & G3957;
  assign G4024 = G3899 & G3926;
  assign G4025 = G3949 & G3911 & G3899;
  assign G4026 = G3911 & G3971 & G3932 & G3899;
  assign G4027 = G3911 & G3979 & G3899 & G3957 & G3932;
  assign G4035 = G3911 & G3949;
  assign G4036 = G3911 & G3932 & G3971;
  assign G4037 = G3911 & G3979 & G3957 & G3932;
  assign G4038 = G3957 & G3911 & G3997 & G3932;
  assign G4039 = G3911 & G3949;
  assign G4040 = G3911 & G3932 & G3971;
  assign G4041 = G3911 & G3979 & G3957 & G3932;
  assign G4042 = G3932 & G3971;
  assign G4043 = G3979 & G3957 & G3932;
  assign G4044 = G3957 & G3997 & G3932;
  assign G4045 = G3932 & G3971;
  assign G4046 = G3979 & G3957 & G3932;
  assign G4047 = G3957 & G3979;
  assign G4051 = G3989 & G3874;
  assign G4052 = G3997 & G3957;
  assign G4184 = ~G4180;
  assign G4193 = ~G4189;
  assign G4247 = G4198;
  assign G4251 = G4198;
  assign G4255 = G4221;
  assign G4259 = G4221;
  assign G4266 = ~G4263;
  assign G4270 = ~G4267;
  assign G4284 = G4263 & G4235 & G4226;
  assign G4287 = G4267 & G4239 & G4230;
  assign G4356 = G4291 & G4300 & G4352 & G4308;
  assign G4361 = G4291 & G4305;
  assign G4362 = G4312 & G4300 & G4291;
  assign G4363 = G4300 & G4314 & G4308 & G4291;
  assign G4369 = G4317 & G4327 & G4336 & G4355 & G4344;
  assign G4372 = G4317 & G4333;
  assign G4373 = G4341 & G4327 & G4317;
  assign G4374 = G4327 & G4348 & G4336 & G4317;
  assign G4375 = G4327 & G4349 & G4317 & G4344 & G4336;
  assign G4567 = ~G4563;
  assign G4581 = ~G4577;
  assign G4590 = ~G4586;
  assign G4601 = ~G4598;
  assign G4605 = ~G4602;
  assign G4606 = G4572;
  assign G4610 = G4572;
  assign G4614 = G4595;
  assign G4618 = G4595;
  assign G4623 = G4598 & G4540 & G4531;
  assign G4626 = G4602 & G4544 & G4535;
  assign G4796 = G3417;
  assign G4804 = G3353;
  assign G4812 = G3365;
  assign G4820 = G3381;
  assign G4828 = G3399;
  assign G4844 = G2409;
  assign G4852 = G2420;
  assign G4860 = G2436;
  assign G4868 = G2454;
  assign G4945 = ~G4939;
  assign G4948 = ~G4939 | ~G4946;
  assign G4986 = ~G4980;
  assign G4989 = ~G4980 | ~G4987;
  assign G5048 = ~G5044;
  assign G5058 = ~G5054;
  assign G5068 = ~G5064;
  assign G5078 = ~G5074;
  assign G5166 = ~G5162;
  assign G5136 = ~G5132;
  assign G5146 = ~G5142;
  assign G5156 = ~G5152;
  assign G5388 = ~G5367 | ~G5368;
  assign G5492 = ~G5488;
  assign G5502 = ~G5498;
  assign G5512 = ~G5508;
  assign G5550 = ~G5546;
  assign G5560 = ~G5556;
  assign G5570 = ~G5566;
  assign G5618 = ~G5614;
  assign G5628 = ~G5624;
  assign G5638 = ~G5634;
  assign G5648 = ~G5644;
  assign G5736 = ~G5732;
  assign G5706 = ~G5702;
  assign G5716 = ~G5712;
  assign G5726 = ~G5722;
  assign G5940 = G2343;
  assign G5948 = G2343;
  assign G5956 = G2354;
  assign G5964 = G2354;
  assign G5972 = G2372;
  assign G5980 = G2372;
  assign G6080 = G2734;
  assign G6090 = G2618;
  assign G6100 = G2589;
  assign G6110 = G2600;
  assign G6138 = G2734;
  assign G6148 = G2618;
  assign G6158 = G2589;
  assign G6168 = G2600;
  assign G6216 = G2701;
  assign G6226 = G2643;
  assign G6236 = G2676;
  assign G6246 = G2655;
  assign G6256 = G2655;
  assign G6267 = ~G6261;
  assign G6304 = G2701;
  assign G6314 = G2643;
  assign G6324 = G2676;
  assign G6342 = ~G6340 | ~G6341;
  assign G6352 = ~G6350 | ~G6351;
  assign G7351 = ~G7345;
  assign G7352 = ~G7348;
  assign G6642 = G3283;
  assign G6650 = G3283;
  assign G6658 = G3295;
  assign G6666 = G3295;
  assign G6674 = G3314;
  assign G6682 = G3314;
  assign G6815 = ~G6809;
  assign G6816 = ~G6812;
  assign G6825 = ~G6819;
  assign G6826 = ~G6822;
  assign G6948 = G3989;
  assign G6958 = G3874;
  assign G6968 = G3845;
  assign G6978 = G3856;
  assign G7006 = G3989;
  assign G7016 = G3874;
  assign G7026 = G3845;
  assign G7036 = G3856;
  assign G7074 = G3997;
  assign G7084 = G3957;
  assign G7094 = G3899;
  assign G7104 = G3932;
  assign G7114 = G3911;
  assign G7124 = G3911;
  assign G7162 = G3997;
  assign G7172 = G3957;
  assign G7182 = G3899;
  assign G7192 = G3932;
  assign G7438 = ~G7436 | ~G7437;
  assign G7617 = ~G7611;
  assign G7618 = ~G7614;
  assign G7609 = ~G7603;
  assign G7610 = ~G7606;
  assign G1151 = G1129 & G1108;
  assign G1002 = G902 & G929;
  assign G933 = ~G929;
  assign G1308 = G1287 & G1221 & G1226;
  assign G1311 = G1291 & G1217 & G1230;
  assign G1314 = G1295 & G1244 & G1249;
  assign G1317 = G1299 & G1240 & G1253;
  assign G1320 = G1303 & G1267 & G1272;
  assign G1323 = G1307 & G1263 & G1276;
  assign G1730 = ~G1726;
  assign G1789 = G1702 & G1726;
  assign G1981 = G1957 & G1935;
  assign G5823 = ~G5817;
  assign G1986 = ~G5817 | ~G5824;
  assign G5831 = ~G5825;
  assign G1989 = ~G5825 | ~G5832;
  assign G5839 = ~G5833;
  assign G1993 = ~G5833 | ~G5840;
  assign G5847 = ~G5841;
  assign G1996 = ~G5841 | ~G5848;
  assign G2000 = ~G5849 | ~G5856;
  assign G2004 = ~G5857 | ~G5864;
  assign G2495 = G2494 | G2493 | G2351 | G2492;
  assign G2515 = G2514 | G2513 | G2512 | G2417 | G2511;
  assign G2757 = G2756 | G2755 | G2597 | G2754;
  assign G2768 = G2629 | G2767;
  assign G2780 = G2779 | G2778 | G2777 | G2652 | G2776;
  assign G2801 = G2715 | G2800;
  assign G3046 = G3028 | G3045;
  assign G3131 = G3130 | G3129 | G3059 | G3128;
  assign G3143 = G3142 | G3141 | G3140 | G3090 | G3139;
  assign G3238 = ~G3235;
  assign G3258 = G3216 & G3235;
  assign G3437 = G3436 | G3435 | G3292 | G3434;
  assign G3453 = G3452 | G3451 | G3450 | G3362 | G3449;
  assign G3595 = G3574 & G3508 & G3513;
  assign G3598 = G3578 & G3504 & G3517;
  assign G4010 = G4009 | G4008 | G3853 | G4007;
  assign G4017 = G3885 | G4016;
  assign G4028 = G4027 | G4026 | G4025 | G3908 | G4024;
  assign G4048 = G3971 | G4047;
  assign G4283 = G4266 & G4230 & G4235;
  assign G4286 = G4270 & G4226 & G4239;
  assign G4364 = G4363 | G4362 | G4297 | G4361;
  assign G4376 = G4375 | G4374 | G4373 | G4324 | G4372;
  assign G4622 = G4601 & G4535 & G4540;
  assign G4625 = G4605 & G4531 & G4544;
  assign G4947 = ~G4942 | ~G4945;
  assign G4988 = ~G4983 | ~G4986;
  assign G5018 = ~G5014;
  assign G5019 = ~G5014 | ~G5017;
  assign G5024 = G950 | G956;
  assign G5038 = ~G5034;
  assign G5106 = ~G5102;
  assign G5107 = ~G5102 | ~G5105;
  assign G5112 = ~G950;
  assign G5126 = ~G5122;
  assign G5468 = G1715 | G1749;
  assign G5482 = ~G5478;
  assign G5526 = ~G1715;
  assign G5540 = ~G5536;
  assign G5588 = ~G5584;
  assign G5589 = ~G5584 | ~G5587;
  assign G5594 = G1746 | G1750;
  assign G5608 = ~G5604;
  assign G5676 = ~G5672;
  assign G5677 = ~G5672 | ~G5675;
  assign G5682 = ~G1746;
  assign G5696 = ~G5692;
  assign G5937 = G2502 | G2501 | G2366 | G2500;
  assign G5945 = ~G2504 & ~G2366 & ~G2503;
  assign G5953 = G2506 | G2384 | G2505;
  assign G5961 = ~G2384 & ~G2507;
  assign G6070 = G2764 | G2763 | G2612 | G2762;
  assign G6128 = ~G2766 & ~G2612 & ~G2765;
  assign G6264 = ~G2799 & ~G2693 & ~G2798;
  assign G6284 = ~G2794 & ~G2793 & ~G2670 & ~G2792;
  assign G6360 = ~G7348 | ~G7351;
  assign G6361 = ~G7345 | ~G7352;
  assign G6639 = G3440 | G3439 | G3308 | G3438;
  assign G6647 = ~G3442 & ~G3308 & ~G3441;
  assign G6655 = G3444 | G3327 | G3443;
  assign G6663 = ~G3327 & ~G3445;
  assign G6817 = ~G6812 | ~G6815;
  assign G6818 = ~G6809 | ~G6816;
  assign G6827 = ~G6822 | ~G6825;
  assign G6828 = ~G6819 | ~G6826;
  assign G6938 = G4013 | G4012 | G3868 | G4011;
  assign G6996 = ~G4015 & ~G3868 & ~G4014;
  assign G7044 = G4044 | G4043 | G3949 | G4042;
  assign G7064 = G4038 | G4037 | G4036 | G3926 | G4035;
  assign G7132 = ~G4046 & ~G3949 & ~G4045;
  assign G7152 = ~G4041 & ~G4040 & ~G3926 & ~G4039;
  assign G7446 = ~G7614 | ~G7617;
  assign G7447 = ~G7611 | ~G7618;
  assign G7456 = ~G7606 | ~G7609;
  assign G7457 = ~G7603 | ~G7610;
  assign G241 = G1117 | G1151;
  assign G265 = G908 | G1002;
  assign G2005 = ~G2003 | ~G2004;
  assign G4800 = ~G4796;
  assign G4808 = ~G4804;
  assign G4816 = ~G4812;
  assign G4824 = ~G4820;
  assign G4832 = ~G4828;
  assign G4848 = ~G4844;
  assign G4856 = ~G4852;
  assign G4864 = ~G4860;
  assign G4872 = ~G4868;
  assign G1310 = ~G1308 & ~G1309;
  assign G1313 = ~G1311 & ~G1312;
  assign G1316 = ~G1314 & ~G1315;
  assign G1319 = ~G1317 & ~G1318;
  assign G1322 = ~G1320 & ~G1321;
  assign G1325 = ~G1323 & ~G1324;
  assign G5392 = ~G5388;
  assign G1790 = G1708 | G1789;
  assign G1982 = G1941 | G1981;
  assign G1985 = ~G5820 | ~G5823;
  assign G1988 = ~G5828 | ~G5831;
  assign G1992 = ~G5836 | ~G5839;
  assign G1995 = ~G5844 | ~G5847;
  assign G2001 = ~G1999 | ~G2000;
  assign G2491 = ~G2487;
  assign G2508 = G2454 & G2409 & G2436 & G2420 & G2472;
  assign G2522 = G2420 & G2454 & G2436 & G4526 & G2472;
  assign G2526 = G2454 & G2436 & G4526 & G2472;
  assign G2529 = G2454 & G4526 & G2472;
  assign G2531 = G4526 & G2472;
  assign G5944 = ~G5940;
  assign G5952 = ~G5948;
  assign G5960 = ~G5956;
  assign G5968 = ~G5964;
  assign G2555 = ~G5972 | ~G5975;
  assign G5976 = ~G5972;
  assign G2559 = ~G5980 | ~G5983;
  assign G5984 = ~G5980;
  assign G2753 = ~G2749;
  assign G2771 = G2643 & G2655 & G2676 & G2742 & G2701;
  assign G2791 = G2701 & G2655 & G2742 & G2676;
  assign G2797 = G2701 & G2742 & G2676;
  assign G2807 = G2742 & G2701;
  assign G6114 = ~G6110;
  assign G6172 = ~G6168;
  assign G6250 = ~G6246;
  assign G6260 = ~G6256;
  assign G6346 = ~G6342;
  assign G6356 = ~G6352;
  assign G3127 = ~G3123;
  assign G3156 = G3123 & G3136;
  assign G3259 = G3223 | G3258;
  assign G3466 = G3431 & G3446;
  assign G6646 = ~G6642;
  assign G6654 = ~G6650;
  assign G6662 = ~G6658;
  assign G6670 = ~G6666;
  assign G3483 = ~G6674 | ~G6677;
  assign G6678 = ~G6674;
  assign G3487 = ~G6682 | ~G6685;
  assign G6686 = ~G6682;
  assign G3582 = ~G3579;
  assign G3586 = ~G3583;
  assign G3590 = ~G3587;
  assign G3594 = ~G3591;
  assign G3597 = ~G3595 & ~G3596;
  assign G3600 = ~G3598 & ~G3599;
  assign G3602 = G3579 & G3536 & G3527;
  assign G3605 = G3583 & G3540 & G3531;
  assign G3608 = G3587 & G3559 & G3550;
  assign G3611 = G3591 & G3563 & G3554;
  assign G4023 = ~G4020;
  assign G6982 = ~G6978;
  assign G7040 = ~G7036;
  assign G7118 = ~G7114;
  assign G7128 = ~G7124;
  assign G4089 = G4004 & G4020;
  assign G4250 = ~G4247;
  assign G4254 = ~G4251;
  assign G4258 = ~G4255;
  assign G4262 = ~G4259;
  assign G4272 = G4247 & G4189 & G4180;
  assign G4275 = G4251 & G4193 & G4184;
  assign G4278 = G4255 & G4212 & G4203;
  assign G4281 = G4259 & G4216 & G4207;
  assign G4285 = ~G4283 & ~G4284;
  assign G4288 = ~G4286 & ~G4287;
  assign G4360 = ~G4356;
  assign G4380 = ~G4369 | ~G89;
  assign G4386 = G4356 & G4369;
  assign G7442 = ~G7438;
  assign G4609 = ~G4606;
  assign G4613 = ~G4610;
  assign G4617 = ~G4614;
  assign G4621 = ~G4618;
  assign G4624 = ~G4622 & ~G4623;
  assign G4627 = ~G4625 & ~G4626;
  assign G4629 = G4606 & G4563 & G4554;
  assign G4632 = G4610 & G4567 & G4558;
  assign G4635 = G4614 & G4586 & G4577;
  assign G4638 = G4618 & G4590 & G4581;
  assign G4836 = G2472;
  assign G4949 = ~G4947 | ~G4948;
  assign G4990 = ~G4988 | ~G4989;
  assign G5020 = ~G5011 | ~G5018;
  assign G5108 = ~G5099 | ~G5106;
  assign G5590 = ~G5581 | ~G5588;
  assign G5678 = ~G5669 | ~G5676;
  assign G6084 = ~G6080;
  assign G6094 = ~G6090;
  assign G6104 = ~G6100;
  assign G6142 = ~G6138;
  assign G6152 = ~G6148;
  assign G6162 = ~G6158;
  assign G6206 = G2742;
  assign G6220 = ~G6216;
  assign G6230 = ~G6226;
  assign G6240 = ~G6236;
  assign G6328 = ~G6324;
  assign G6294 = G2742;
  assign G6308 = ~G6304;
  assign G6318 = ~G6314;
  assign G6362 = ~G6360 | ~G6361;
  assign G6840 = ~G6817 | ~G6818;
  assign G6848 = ~G6827 | ~G6828;
  assign G6952 = ~G6948;
  assign G6962 = ~G6958;
  assign G6972 = ~G6968;
  assign G7010 = ~G7006;
  assign G7020 = ~G7016;
  assign G7030 = ~G7026;
  assign G7078 = ~G7074;
  assign G7088 = ~G7084;
  assign G7098 = ~G7094;
  assign G7108 = ~G7104;
  assign G7196 = ~G7192;
  assign G7166 = ~G7162;
  assign G7176 = ~G7172;
  assign G7186 = ~G7182;
  assign G7448 = ~G7446 | ~G7447;
  assign G7458 = ~G7456 | ~G7457;
  assign G254 = G3046 & G3249;
  assign G260 = G3046 & G3249;
  assign G1987 = ~G1985 | ~G1986;
  assign G1994 = ~G1992 | ~G1993;
  assign G2002 = ~G2001;
  assign G962 = G933 & G924;
  assign G1751 = G1730 & G1721;
  assign G1990 = ~G1988 | ~G1989;
  assign G1997 = ~G1995 | ~G1996;
  assign G2499 = ~G2495;
  assign G2536 = G2515 & G2487;
  assign G5943 = ~G5937;
  assign G2542 = ~G5937 | ~G5944;
  assign G5951 = ~G5945;
  assign G2545 = ~G5945 | ~G5952;
  assign G5959 = ~G5953;
  assign G2549 = ~G5953 | ~G5960;
  assign G5967 = ~G5961;
  assign G2552 = ~G5961 | ~G5968;
  assign G2556 = ~G5969 | ~G5976;
  assign G2560 = ~G5977 | ~G5984;
  assign G2761 = ~G2757;
  assign G2784 = ~G2780;
  assign G2853 = G2749 & G2780;
  assign G3135 = ~G3131;
  assign G3146 = ~G3143;
  assign G3163 = G3123 & G3143;
  assign G3467 = G3453 & G3431;
  assign G6645 = ~G6639;
  assign G3470 = ~G6639 | ~G6646;
  assign G6653 = ~G6647;
  assign G3473 = ~G6647 | ~G6654;
  assign G6661 = ~G6655;
  assign G3477 = ~G6655 | ~G6662;
  assign G6669 = ~G6663;
  assign G3480 = ~G6663 | ~G6670;
  assign G3484 = ~G6671 | ~G6678;
  assign G3488 = ~G6679 | ~G6686;
  assign G3601 = G3582 & G3531 & G3536;
  assign G3604 = G3586 & G3527 & G3540;
  assign G3607 = G3590 & G3554 & G3559;
  assign G3610 = G3594 & G3550 & G3563;
  assign G4032 = ~G4028;
  assign G4090 = G4004 & G4028;
  assign G4271 = G4250 & G4184 & G4189;
  assign G4274 = G4254 & G4180 & G4193;
  assign G4277 = G4258 & G4207 & G4212;
  assign G4280 = G4262 & G4203 & G4216;
  assign G4368 = ~G4364;
  assign G4379 = ~G4376;
  assign G4387 = G4356 & G4376;
  assign G4628 = G4609 & G4558 & G4563;
  assign G4631 = G4613 & G4554 & G4567;
  assign G4634 = G4617 & G4581 & G4586;
  assign G4637 = G4621 & G4577 & G4590;
  assign G4841 = G2522 | G2520 | G2519 | G2431 | G2518;
  assign G4849 = G2526 | G2524 | G2448 | G2523;
  assign G4857 = G2529 | G2465 | G2527;
  assign G4865 = G2481 | G2531;
  assign G5021 = ~G5019 | ~G5020;
  assign G5028 = ~G5024;
  assign G5109 = ~G5107 | ~G5108;
  assign G5116 = ~G5112;
  assign G5369 = ~G1313 | ~G1310;
  assign G5377 = ~G1319 | ~G1316;
  assign G5385 = ~G1325 | ~G1322;
  assign G5472 = ~G5468;
  assign G5473 = ~G5468 | ~G5471;
  assign G5530 = ~G5526;
  assign G5531 = ~G5526 | ~G5529;
  assign G5591 = ~G5589 | ~G5590;
  assign G5598 = ~G5594;
  assign G5679 = ~G5677 | ~G5678;
  assign G5686 = ~G5682;
  assign G6060 = G2768 | G2804;
  assign G6074 = ~G6070;
  assign G6118 = ~G2768;
  assign G6132 = ~G6128;
  assign G6176 = G2797 | G2796 | G2693 | G2795;
  assign G6186 = G2801 | G2807;
  assign G6196 = G2791 | G2790 | G2789 | G2670 | G2788;
  assign G6268 = ~G6264;
  assign G6269 = ~G6264 | ~G6267;
  assign G6274 = ~G2801;
  assign G6288 = ~G6284;
  assign G6337 = ~G4288 | ~G4285;
  assign G6829 = ~G3600 | ~G3597;
  assign G6928 = G4017 | G4051;
  assign G6942 = ~G6938;
  assign G6986 = ~G4017;
  assign G7000 = ~G6996;
  assign G7048 = ~G7044;
  assign G7049 = ~G7044 | ~G7047;
  assign G7054 = G4048 | G4052;
  assign G7068 = ~G7064;
  assign G7136 = ~G7132;
  assign G7137 = ~G7132 | ~G7135;
  assign G7142 = ~G4048;
  assign G7156 = ~G7152;
  assign G7433 = ~G4627 | ~G4624;
  assign G242 = G1982 & G1146;
  assign G3151 = ~G3135 | ~G3127;
  assign G257 = G3249 & G3035 & G3156 & G89 & G4386;
  assign G263 = G3249 & G3035 & G3156 & G89 & G4386;
  assign G266 = G1790 & G997;
  assign G1991 = ~G1990;
  assign G1998 = ~G1997;
  assign G3489 = ~G3487 | ~G3488;
  assign G371 = ~G4836 | ~G4839;
  assign G4840 = ~G4836;
  assign G2561 = ~G2559 | ~G2560;
  assign G2532 = G2487 & G2508;
  assign G2537 = G2495 | G2536;
  assign G2541 = ~G5940 | ~G5943;
  assign G2544 = ~G5948 | ~G5951;
  assign G2548 = ~G5956 | ~G5959;
  assign G2551 = ~G5964 | ~G5967;
  assign G2557 = ~G2555 | ~G2556;
  assign G2563 = G2508 & G4526;
  assign G2577 = ~G2499 | ~G2491;
  assign G2775 = ~G2771;
  assign G2806 = ~G2771 | ~G4526;
  assign G2808 = ~G2761 | ~G2753;
  assign G2852 = G2749 & G2771;
  assign G2854 = G2757 | G2853;
  assign G6366 = ~G6362;
  assign G4381 = ~G4368 | ~G4360;
  assign G3164 = G3131 | G3163;
  assign G3241 = G3035 & G3156 & G89 & G4386;
  assign G3468 = G3437 | G3467;
  assign G3469 = ~G6642 | ~G6645;
  assign G3472 = ~G6650 | ~G6653;
  assign G3476 = ~G6658 | ~G6661;
  assign G3479 = ~G6666 | ~G6669;
  assign G3485 = ~G3483 | ~G3484;
  assign G3603 = ~G3601 & ~G3602;
  assign G3606 = ~G3604 & ~G3605;
  assign G3609 = ~G3607 & ~G3608;
  assign G3612 = ~G3610 & ~G3611;
  assign G6844 = ~G6840;
  assign G6852 = ~G6848;
  assign G4091 = G4010 | G4090;
  assign G4273 = ~G4271 & ~G4272;
  assign G4276 = ~G4274 & ~G4275;
  assign G4279 = ~G4277 & ~G4278;
  assign G4282 = ~G4280 & ~G4281;
  assign G4382 = G4379 & G4380;
  assign G4388 = G4364 | G4387;
  assign G7452 = ~G7448;
  assign G7462 = ~G7458;
  assign G4630 = ~G4628 & ~G4629;
  assign G4633 = ~G4631 & ~G4632;
  assign G4636 = ~G4634 & ~G4635;
  assign G4639 = ~G4637 & ~G4638;
  assign G4955 = ~G4949;
  assign G4958 = ~G4949 | ~G4956;
  assign G4996 = ~G4990;
  assign G4999 = ~G4990 | ~G4997;
  assign G5474 = ~G5465 | ~G5472;
  assign G5532 = ~G5523 | ~G5530;
  assign G6210 = ~G6206;
  assign G6270 = ~G6261 | ~G6268;
  assign G6298 = ~G6294;
  assign G7050 = ~G7041 | ~G7048;
  assign G7138 = ~G7129 | ~G7136;
  assign G3471 = ~G3469 | ~G3470;
  assign G3478 = ~G3476 | ~G3477;
  assign G3486 = ~G3485;
  assign G372 = ~G4833 | ~G4840;
  assign G2543 = ~G2541 | ~G2542;
  assign G2550 = ~G2548 | ~G2549;
  assign G2558 = ~G2557;
  assign G4847 = ~G4841;
  assign G387 = ~G4841 | ~G4848;
  assign G4855 = ~G4849;
  assign G390 = ~G4849 | ~G4856;
  assign G4863 = ~G4857;
  assign G393 = ~G4857 | ~G4864;
  assign G4871 = ~G4865;
  assign G396 = ~G4865 | ~G4872;
  assign G965 = ~G962;
  assign G5375 = ~G5369;
  assign G1327 = ~G5369 | ~G5376;
  assign G5383 = ~G5377;
  assign G1330 = ~G5377 | ~G5384;
  assign G5391 = ~G5385;
  assign G1333 = ~G5385 | ~G5392;
  assign G1754 = ~G1751;
  assign G2546 = ~G2544 | ~G2545;
  assign G2553 = ~G2551 | ~G2552;
  assign G2564 = G2515 | G2563;
  assign G2809 = G2784 & G2806;
  assign G2813 = G2784 & G2775;
  assign G6345 = ~G6337;
  assign G2860 = ~G6337 | ~G6346;
  assign G3474 = ~G3472 | ~G3473;
  assign G3481 = ~G3479 | ~G3480;
  assign G6835 = ~G6829;
  assign G3614 = ~G6829 | ~G6836;
  assign G4053 = G4032 & G4023;
  assign G7441 = ~G7433;
  assign G4516 = ~G7433 | ~G7442;
  assign G4957 = ~G4952 | ~G4955;
  assign G4998 = ~G4993 | ~G4996;
  assign G5027 = ~G5021;
  assign G5030 = ~G5021 | ~G5028;
  assign G5115 = ~G5109;
  assign G5118 = ~G5109 | ~G5116;
  assign G5475 = ~G5473 | ~G5474;
  assign G5533 = ~G5531 | ~G5532;
  assign G5597 = ~G5591;
  assign G5600 = ~G5591 | ~G5598;
  assign G5685 = ~G5679;
  assign G5688 = ~G5679 | ~G5686;
  assign G6064 = ~G6060;
  assign G6065 = ~G6060 | ~G6063;
  assign G6122 = ~G6118;
  assign G6123 = ~G6118 | ~G6121;
  assign G6180 = ~G6176;
  assign G6181 = ~G6176 | ~G6179;
  assign G6190 = ~G6186;
  assign G6200 = ~G6196;
  assign G6271 = ~G6269 | ~G6270;
  assign G6278 = ~G6274;
  assign G6347 = ~G4276 | ~G4273;
  assign G6357 = ~G4282 | ~G4279;
  assign G6837 = ~G3606 | ~G3603;
  assign G6845 = ~G3612 | ~G3609;
  assign G6932 = ~G6928;
  assign G6933 = ~G6928 | ~G6931;
  assign G6990 = ~G6986;
  assign G6991 = ~G6986 | ~G6989;
  assign G7051 = ~G7049 | ~G7050;
  assign G7058 = ~G7054;
  assign G7139 = ~G7137 | ~G7138;
  assign G7146 = ~G7142;
  assign G7443 = ~G4639 | ~G4636;
  assign G7453 = ~G4633 | ~G4630;
  assign G243 = G1146 & G3468 & G1974;
  assign G244 = G1146 & G1974 & G2537 & G3466;
  assign G245 = G1146 & G1974 & G3466 & G4526 & G2532;
  assign G255 = G3249 & G3164 & G3035;
  assign G256 = G3249 & G3035 & G4388 & G3156;
  assign G261 = G3249 & G3164 & G3035;
  assign G262 = G3249 & G3035 & G4388 & G3156;
  assign G267 = G997 & G4091 & G1788;
  assign G268 = G997 & G1788 & G2854 & G4089;
  assign G269 = G997 & G1788 & G4089 & G4526 & G2852;
  assign G3475 = ~G3474;
  assign G3482 = ~G3481;
  assign G373 = ~G371 | ~G372;
  assign G2547 = ~G2546;
  assign G2554 = ~G2553;
  assign G386 = ~G4844 | ~G4847;
  assign G389 = ~G4852 | ~G4855;
  assign G392 = ~G4860 | ~G4863;
  assign G395 = ~G4868 | ~G4871;
  assign G1326 = ~G5372 | ~G5375;
  assign G1329 = ~G5380 | ~G5383;
  assign G1332 = ~G5388 | ~G5391;
  assign G1436 = G4091 & G1788;
  assign G1440 = G1788 & G2854 & G4089;
  assign G1445 = G1788 & G4089 & G4526 & G2852;
  assign G1450 = G2854 & G4089;
  assign G1454 = G4089 & G4526 & G2852;
  assign G2859 = ~G6342 | ~G6345;
  assign G4385 = ~G4382;
  assign G3148 = G4382 & G4364;
  assign G3239 = G3164 & G3035;
  assign G3240 = G3035 & G4388 & G3156;
  assign G3265 = G3468 & G1974;
  assign G3267 = G1974 & G2537 & G3466;
  assign G3270 = G1974 & G3466 & G4526 & G2532;
  assign G3274 = G2537 & G3466;
  assign G3277 = G3466 & G4526 & G2532;
  assign G3613 = ~G6832 | ~G6835;
  assign G4515 = ~G7438 | ~G7441;
  assign G4959 = ~G4957 | ~G4958;
  assign G5000 = ~G4998 | ~G4999;
  assign G5029 = ~G5024 | ~G5027;
  assign G5117 = ~G5112 | ~G5115;
  assign G5599 = ~G5594 | ~G5597;
  assign G5687 = ~G5682 | ~G5685;
  assign G6066 = ~G6057 | ~G6064;
  assign G6124 = ~G6115 | ~G6122;
  assign G6182 = ~G6173 | ~G6180;
  assign G6934 = ~G6925 | ~G6932;
  assign G6992 = ~G6983 | ~G6990;
  assign G246 = G245 | G244 | G243 | G241 | G242;
  assign G258 = G257 | G256 | G255 | G3259 | G254;
  assign G264 = G263 | G262 | G261 | G3259 | G260;
  assign G270 = G269 | G268 | G267 | G265 | G266;
  assign G375 = G2564 & G2543;
  assign G378 = G2564 & G2550;
  assign G381 = G2564 & G2558;
  assign G384 = G2564 & G2406;
  assign G388 = ~G386 | ~G387;
  assign G391 = ~G389 | ~G390;
  assign G394 = ~G392 | ~G393;
  assign G397 = ~G395 | ~G396;
  assign G1328 = ~G1326 | ~G1327;
  assign G1331 = ~G1329 | ~G1330;
  assign G1334 = ~G1332 | ~G1333;
  assign G1447 = G1445 | G1440 | G1790 | G1436;
  assign G1766 = G1454 | G4091 | G1450;
  assign G2571 = ~G2564;
  assign G2579 = G2577 & G2564;
  assign G2812 = ~G2809;
  assign G2816 = ~G2813;
  assign G2851 = G2809 & G2757;
  assign G2861 = ~G2859 | ~G2860;
  assign G6355 = ~G6347;
  assign G2863 = ~G6347 | ~G6356;
  assign G6365 = ~G6357;
  assign G2866 = ~G6357 | ~G6366;
  assign G3147 = G4381 & G4385;
  assign G3242 = G3241 | G3240 | G3046 | G3239;
  assign G3271 = G3270 | G3267 | G1982 | G3265;
  assign G3279 = G3277 | G3468 | G3274;
  assign G3615 = ~G3613 | ~G3614;
  assign G6843 = ~G6837;
  assign G3617 = ~G6837 | ~G6844;
  assign G6851 = ~G6845;
  assign G3620 = ~G6845 | ~G6852;
  assign G4056 = ~G4053;
  assign G4517 = ~G4515 | ~G4516;
  assign G7451 = ~G7443;
  assign G4519 = ~G7443 | ~G7452;
  assign G7461 = ~G7453;
  assign G4522 = ~G7453 | ~G7462;
  assign G5031 = ~G5029 | ~G5030;
  assign G5119 = ~G5117 | ~G5118;
  assign G5481 = ~G5475;
  assign G5484 = ~G5475 | ~G5482;
  assign G5539 = ~G5533;
  assign G5542 = ~G5533 | ~G5540;
  assign G5601 = ~G5599 | ~G5600;
  assign G5689 = ~G5687 | ~G5688;
  assign G6067 = ~G6065 | ~G6066;
  assign G6125 = ~G6123 | ~G6124;
  assign G6183 = ~G6181 | ~G6182;
  assign G6277 = ~G6271;
  assign G6280 = ~G6271 | ~G6278;
  assign G6935 = ~G6933 | ~G6934;
  assign G6993 = ~G6991 | ~G6992;
  assign G7057 = ~G7051;
  assign G7060 = ~G7051 | ~G7058;
  assign G7145 = ~G7139;
  assign G7148 = ~G7139 | ~G7146;
  assign G4968 = ~G4959 | ~G4966;
  assign G5009 = ~G5000 | ~G5007;
  assign G2850 = G2808 & G2812;
  assign G2862 = ~G6352 | ~G6355;
  assign G2865 = ~G6362 | ~G6365;
  assign G3149 = G3147 | G3148;
  assign G3243 = ~G3228 | ~G3242;
  assign G3616 = ~G6840 | ~G6843;
  assign G3619 = ~G6848 | ~G6851;
  assign G4518 = ~G7448 | ~G7451;
  assign G4521 = ~G7458 | ~G7461;
  assign G4965 = ~G4959;
  assign G5006 = ~G5000;
  assign G5483 = ~G5478 | ~G5481;
  assign G5541 = ~G5536 | ~G5539;
  assign G6279 = ~G6274 | ~G6277;
  assign G7059 = ~G7054 | ~G7057;
  assign G7147 = ~G7142 | ~G7145;
  assign G374 = G2547 & G2571;
  assign G377 = G2554 & G2571;
  assign G380 = G2561 & G2571;
  assign G383 = G2400 & G2571;
  assign G955 = ~G920 | ~G1447;
  assign G4967 = ~G4962 | ~G4965;
  assign G5008 = ~G5003 | ~G5006;
  assign G975 = G1447;
  assign G1136 = G1038 & G1074 & G1055 & G3271 & G1093;
  assign G1140 = G1074 & G1055 & G3271 & G1093;
  assign G1143 = G1074 & G3271 & G1093;
  assign G1145 = G3271 & G1093;
  assign G1160 = G1122 & G3271;
  assign G1771 = ~G1766;
  assign G1964 = G1869 & G1903 & G1885 & G3279 & G1921;
  assign G1968 = G1903 & G1885 & G3279 & G1921;
  assign G1971 = G1903 & G3279 & G1921;
  assign G1973 = G3279 & G1921;
  assign G2007 = G1950 & G3279;
  assign G2578 = G2495 & G2571;
  assign G2864 = ~G2862 | ~G2863;
  assign G2867 = ~G2865 | ~G2866;
  assign G3150 = ~G3136 | ~G3149;
  assign G3245 = G3238 & G3243;
  assign G3618 = ~G3616 | ~G3617;
  assign G3621 = ~G3619 | ~G3620;
  assign G4067 = G2850 | G2851;
  assign G4520 = ~G4518 | ~G4519;
  assign G4523 = ~G4521 | ~G4522;
  assign G4713 = G3279;
  assign G4753 = G3271;
  assign G5037 = ~G5031;
  assign G5040 = ~G5031 | ~G5038;
  assign G5125 = ~G5119;
  assign G5128 = ~G5119 | ~G5126;
  assign G5485 = ~G5483 | ~G5484;
  assign G5543 = ~G5541 | ~G5542;
  assign G5607 = ~G5601;
  assign G5610 = ~G5601 | ~G5608;
  assign G5695 = ~G5689;
  assign G5698 = ~G5689 | ~G5696;
  assign G6073 = ~G6067;
  assign G6076 = ~G6067 | ~G6074;
  assign G6131 = ~G6125;
  assign G6134 = ~G6125 | ~G6132;
  assign G6189 = ~G6183;
  assign G6192 = ~G6183 | ~G6190;
  assign G6281 = ~G6279 | ~G6280;
  assign G6941 = ~G6935;
  assign G6944 = ~G6935 | ~G6942;
  assign G6999 = ~G6993;
  assign G7002 = ~G6993 | ~G7000;
  assign G7061 = ~G7059 | ~G7060;
  assign G7149 = ~G7147 | ~G7148;
  assign G376 = G374 | G375;
  assign G379 = G377 | G378;
  assign G382 = G380 | G381;
  assign G385 = G383 | G384;
  assign G958 = G933 & G955;
  assign G967 = ~G4967 | ~G4968;
  assign G971 = ~G5008 | ~G5009;
  assign G1161 = G1129 | G1160;
  assign G2008 = G1957 | G2007;
  assign G2580 = G2578 | G2579;
  assign G2868 = G2867 & G2864 & G1331 & G2861;
  assign G3152 = G3146 & G3150;
  assign G4443 = G3621 & G3618 & G1328 & G1334;
  assign G4524 = G4523 & G4520 & G3615 & G4517;
  assign G4721 = G1964 | G1962 | G1961 | G1880 | G1960;
  assign G4729 = G1968 | G1966 | G1897 | G1965;
  assign G4737 = G1971 | G1914 | G1969;
  assign G4745 = G1929 | G1973;
  assign G4761 = G1136 | G1134 | G1133 | G1050 | G1132;
  assign G4769 = G1140 | G1138 | G1068 | G1137;
  assign G4777 = G1143 | G1086 | G1141;
  assign G4785 = G1102 | G1145;
  assign G5039 = ~G5034 | ~G5037;
  assign G5127 = ~G5122 | ~G5125;
  assign G5609 = ~G5604 | ~G5607;
  assign G5697 = ~G5692 | ~G5695;
  assign G6075 = ~G6070 | ~G6073;
  assign G6133 = ~G6128 | ~G6131;
  assign G6191 = ~G6186 | ~G6189;
  assign G6943 = ~G6938 | ~G6941;
  assign G7001 = ~G6996 | ~G6999;
  assign G3248 = ~G3245;
  assign G248 = G3245 & G3223;
  assign G4719 = ~G4713;
  assign G294 = ~G4713 | ~G4720;
  assign G4759 = ~G4753;
  assign G323 = ~G4753 | ~G4760;
  assign G980 = ~G975;
  assign G4072 = ~G4067;
  assign G5041 = ~G5039 | ~G5040;
  assign G5129 = ~G5127 | ~G5128;
  assign G5491 = ~G5485;
  assign G5494 = ~G5485 | ~G5492;
  assign G5549 = ~G5543;
  assign G5552 = ~G5543 | ~G5550;
  assign G5611 = ~G5609 | ~G5610;
  assign G5699 = ~G5697 | ~G5698;
  assign G6077 = ~G6075 | ~G6076;
  assign G6135 = ~G6133 | ~G6134;
  assign G6193 = ~G6191 | ~G6192;
  assign G6287 = ~G6281;
  assign G6290 = ~G6281 | ~G6288;
  assign G6945 = ~G6943 | ~G6944;
  assign G7003 = ~G7001 | ~G7002;
  assign G7067 = ~G7061;
  assign G7070 = ~G7061 | ~G7068;
  assign G7155 = ~G7149;
  assign G7158 = ~G7149 | ~G7156;
  assign G247 = G3244 & G3248;
  assign G3155 = ~G3152;
  assign G251 = G3152 & G3131;
  assign G272 = G1176 & G1161;
  assign G961 = ~G958;
  assign G275 = G958 & G908;
  assign G293 = ~G4716 | ~G4719;
  assign G297 = G2008 & G1987;
  assign G300 = G2008 & G1994;
  assign G303 = G2008 & G2002;
  assign G306 = G2008 & G1856;
  assign G4727 = ~G4721;
  assign G309 = ~G4721 | ~G4728;
  assign G4735 = ~G4729;
  assign G312 = ~G4729 | ~G4736;
  assign G4743 = ~G4737;
  assign G315 = ~G4737 | ~G4744;
  assign G4751 = ~G4745;
  assign G318 = ~G4745 | ~G4752;
  assign G322 = ~G4756 | ~G4759;
  assign G4767 = ~G4761;
  assign G326 = ~G4761 | ~G4768;
  assign G4775 = ~G4769;
  assign G329 = ~G4769 | ~G4776;
  assign G4783 = ~G4777;
  assign G332 = ~G4777 | ~G4784;
  assign G4791 = ~G4785;
  assign G335 = ~G4785 | ~G4792;
  assign G412 = ~G4443;
  assign G414 = ~G4524;
  assign G416 = ~G2868;
  assign G2881 = G2868 & G4443 & G4524;
  assign G993 = G975 & G971 & G962;
  assign G994 = G975 & G967 & G965;
  assign G1166 = ~G1161;
  assign G1171 = G1161 & G1155;
  assign G1174 = G1161 & G1023;
  assign G2014 = ~G2008;
  assign G3459 = G3365 & G3399 & G3381 & G2580 & G3417;
  assign G3462 = G3399 & G3381 & G2580 & G3417;
  assign G3464 = G3399 & G2580 & G3417;
  assign G3465 = G2580 & G3417;
  assign G3490 = G3446 & G2580;
  assign G4793 = G2580;
  assign G5493 = ~G5488 | ~G5491;
  assign G5551 = ~G5546 | ~G5549;
  assign G6289 = ~G6284 | ~G6287;
  assign G7069 = ~G7064 | ~G7067;
  assign G7157 = ~G7152 | ~G7155;
  assign G249 = G247 | G248;
  assign G250 = G3151 & G3155;
  assign G274 = G957 & G961;
  assign G295 = ~G293 | ~G294;
  assign G308 = ~G4724 | ~G4727;
  assign G311 = ~G4732 | ~G4735;
  assign G314 = ~G4740 | ~G4743;
  assign G317 = ~G4748 | ~G4751;
  assign G324 = ~G322 | ~G323;
  assign G325 = ~G4764 | ~G4767;
  assign G328 = ~G4772 | ~G4775;
  assign G331 = ~G4780 | ~G4783;
  assign G334 = ~G4788 | ~G4791;
  assign G417 = G2881 & G2876 & G2878;
  assign G991 = G980 & G971 & G933;
  assign G992 = G980 & G967 & G929;
  assign G3491 = G3453 | G3490;
  assign G4801 = G3459 | G3458 | G3457 | G3376 | G3456;
  assign G4809 = G3462 | G3461 | G3393 | G3460;
  assign G4817 = G3464 | G3410 | G3463;
  assign G4825 = G3425 | G3465;
  assign G5047 = ~G5041;
  assign G5050 = ~G5041 | ~G5048;
  assign G5135 = ~G5129;
  assign G5138 = ~G5129 | ~G5136;
  assign G5495 = ~G5493 | ~G5494;
  assign G5553 = ~G5551 | ~G5552;
  assign G5617 = ~G5611;
  assign G5620 = ~G5611 | ~G5618;
  assign G5705 = ~G5699;
  assign G5708 = ~G5699 | ~G5706;
  assign G6083 = ~G6077;
  assign G6086 = ~G6077 | ~G6084;
  assign G6141 = ~G6135;
  assign G6144 = ~G6135 | ~G6142;
  assign G6199 = ~G6193;
  assign G6202 = ~G6193 | ~G6200;
  assign G6291 = ~G6289 | ~G6290;
  assign G6951 = ~G6945;
  assign G6954 = ~G6945 | ~G6952;
  assign G7009 = ~G7003;
  assign G7012 = ~G7003 | ~G7010;
  assign G7071 = ~G7069 | ~G7070;
  assign G7159 = ~G7157 | ~G7158;
  assign G252 = G250 | G251;
  assign G271 = G1117 & G1166;
  assign G276 = G274 | G275;
  assign G296 = G1991 & G2014;
  assign G299 = G1998 & G2014;
  assign G302 = G2005 & G2014;
  assign G305 = G1850 & G2014;
  assign G310 = ~G308 | ~G309;
  assign G313 = ~G311 | ~G312;
  assign G316 = ~G314 | ~G315;
  assign G319 = ~G317 | ~G318;
  assign G327 = ~G325 | ~G326;
  assign G330 = ~G328 | ~G329;
  assign G333 = ~G331 | ~G332;
  assign G336 = ~G334 | ~G335;
  assign G4799 = ~G4793;
  assign G343 = ~G4793 | ~G4800;
  assign G418 = ~G417;
  assign G1170 = G1158 & G1166;
  assign G1173 = G1019 & G1166;
  assign G5049 = ~G5044 | ~G5047;
  assign G5137 = ~G5132 | ~G5135;
  assign G5167 = G994 | G993 | G991 | G992;
  assign G5619 = ~G5614 | ~G5617;
  assign G5707 = ~G5702 | ~G5705;
  assign G6085 = ~G6080 | ~G6083;
  assign G6143 = ~G6138 | ~G6141;
  assign G6201 = ~G6196 | ~G6199;
  assign G6953 = ~G6948 | ~G6951;
  assign G7011 = ~G7006 | ~G7009;
  assign G273 = G271 | G272;
  assign G298 = G296 | G297;
  assign G301 = G299 | G300;
  assign G304 = G302 | G303;
  assign G307 = G305 | G306;
  assign G342 = ~G4796 | ~G4799;
  assign G346 = G3491 & G3471;
  assign G349 = G3491 & G3478;
  assign G352 = G3491 & G3486;
  assign G355 = G3491 & G3350;
  assign G4807 = ~G4801;
  assign G358 = ~G4801 | ~G4808;
  assign G4815 = ~G4809;
  assign G361 = ~G4809 | ~G4816;
  assign G4823 = ~G4817;
  assign G364 = ~G4817 | ~G4824;
  assign G4831 = ~G4825;
  assign G367 = ~G4825 | ~G4832;
  assign G1172 = G1170 | G1171;
  assign G1175 = G1173 | G1174;
  assign G3497 = ~G3491;
  assign G5051 = ~G5049 | ~G5050;
  assign G5139 = ~G5137 | ~G5138;
  assign G5501 = ~G5495;
  assign G5504 = ~G5495 | ~G5502;
  assign G5559 = ~G5553;
  assign G5562 = ~G5553 | ~G5560;
  assign G5621 = ~G5619 | ~G5620;
  assign G5709 = ~G5707 | ~G5708;
  assign G6087 = ~G6085 | ~G6086;
  assign G6145 = ~G6143 | ~G6144;
  assign G6203 = ~G6201 | ~G6202;
  assign G6297 = ~G6291;
  assign G6300 = ~G6291 | ~G6298;
  assign G6955 = ~G6953 | ~G6954;
  assign G7013 = ~G7011 | ~G7012;
  assign G7077 = ~G7071;
  assign G7080 = ~G7071 | ~G7078;
  assign G7165 = ~G7159;
  assign G7168 = ~G7159 | ~G7166;
  assign G344 = ~G342 | ~G343;
  assign G357 = ~G4804 | ~G4807;
  assign G360 = ~G4812 | ~G4815;
  assign G363 = ~G4820 | ~G4823;
  assign G366 = ~G4828 | ~G4831;
  assign G5173 = ~G5167;
  assign G422 = G1172;
  assign G469 = G1172;
  assign G419 = G1175;
  assign G471 = G1175;
  assign G5503 = ~G5498 | ~G5501;
  assign G5561 = ~G5556 | ~G5559;
  assign G6299 = ~G6294 | ~G6297;
  assign G7079 = ~G7074 | ~G7077;
  assign G7167 = ~G7162 | ~G7165;
  assign G345 = G3475 & G3497;
  assign G348 = G3482 & G3497;
  assign G351 = G3489 & G3497;
  assign G354 = G3344 & G3497;
  assign G359 = ~G357 | ~G358;
  assign G362 = ~G360 | ~G361;
  assign G365 = ~G363 | ~G364;
  assign G368 = ~G366 | ~G367;
  assign G5057 = ~G5051;
  assign G5060 = ~G5051 | ~G5058;
  assign G5145 = ~G5139;
  assign G5148 = ~G5139 | ~G5146;
  assign G5505 = ~G5503 | ~G5504;
  assign G5563 = ~G5561 | ~G5562;
  assign G5627 = ~G5621;
  assign G5630 = ~G5621 | ~G5628;
  assign G5715 = ~G5709;
  assign G5718 = ~G5709 | ~G5716;
  assign G6093 = ~G6087;
  assign G6096 = ~G6087 | ~G6094;
  assign G6151 = ~G6145;
  assign G6154 = ~G6145 | ~G6152;
  assign G6209 = ~G6203;
  assign G6212 = ~G6203 | ~G6210;
  assign G6301 = ~G6299 | ~G6300;
  assign G6961 = ~G6955;
  assign G6964 = ~G6955 | ~G6962;
  assign G7019 = ~G7013;
  assign G7022 = ~G7013 | ~G7020;
  assign G7081 = ~G7079 | ~G7080;
  assign G7169 = ~G7167 | ~G7168;
  assign G347 = G345 | G346;
  assign G350 = G348 | G349;
  assign G353 = G351 | G352;
  assign G356 = G354 | G355;
  assign G5059 = ~G5054 | ~G5057;
  assign G5147 = ~G5142 | ~G5145;
  assign G5629 = ~G5624 | ~G5627;
  assign G5717 = ~G5712 | ~G5715;
  assign G6095 = ~G6090 | ~G6093;
  assign G6153 = ~G6148 | ~G6151;
  assign G6211 = ~G6206 | ~G6209;
  assign G6963 = ~G6958 | ~G6961;
  assign G7021 = ~G7016 | ~G7019;
  assign G5061 = ~G5059 | ~G5060;
  assign G5149 = ~G5147 | ~G5148;
  assign G5511 = ~G5505;
  assign G5514 = ~G5505 | ~G5512;
  assign G5569 = ~G5563;
  assign G5572 = ~G5563 | ~G5570;
  assign G5631 = ~G5629 | ~G5630;
  assign G5719 = ~G5717 | ~G5718;
  assign G6097 = ~G6095 | ~G6096;
  assign G6155 = ~G6153 | ~G6154;
  assign G6213 = ~G6211 | ~G6212;
  assign G6307 = ~G6301;
  assign G6310 = ~G6301 | ~G6308;
  assign G6965 = ~G6963 | ~G6964;
  assign G7023 = ~G7021 | ~G7022;
  assign G7087 = ~G7081;
  assign G7090 = ~G7081 | ~G7088;
  assign G7175 = ~G7169;
  assign G7178 = ~G7169 | ~G7176;
  assign G5513 = ~G5508 | ~G5511;
  assign G5571 = ~G5566 | ~G5569;
  assign G6309 = ~G6304 | ~G6307;
  assign G7089 = ~G7084 | ~G7087;
  assign G7177 = ~G7172 | ~G7175;
  assign G5067 = ~G5061;
  assign G5070 = ~G5061 | ~G5068;
  assign G5155 = ~G5149;
  assign G5158 = ~G5149 | ~G5156;
  assign G5515 = ~G5513 | ~G5514;
  assign G5573 = ~G5571 | ~G5572;
  assign G5637 = ~G5631;
  assign G5640 = ~G5631 | ~G5638;
  assign G5725 = ~G5719;
  assign G5728 = ~G5719 | ~G5726;
  assign G6103 = ~G6097;
  assign G6106 = ~G6097 | ~G6104;
  assign G6161 = ~G6155;
  assign G6164 = ~G6155 | ~G6162;
  assign G6219 = ~G6213;
  assign G6222 = ~G6213 | ~G6220;
  assign G6311 = ~G6309 | ~G6310;
  assign G6971 = ~G6965;
  assign G6974 = ~G6965 | ~G6972;
  assign G7029 = ~G7023;
  assign G7032 = ~G7023 | ~G7030;
  assign G7091 = ~G7089 | ~G7090;
  assign G7179 = ~G7177 | ~G7178;
  assign G5069 = ~G5064 | ~G5067;
  assign G5157 = ~G5152 | ~G5155;
  assign G5639 = ~G5634 | ~G5637;
  assign G5727 = ~G5722 | ~G5725;
  assign G6105 = ~G6100 | ~G6103;
  assign G6163 = ~G6158 | ~G6161;
  assign G6221 = ~G6216 | ~G6219;
  assign G6973 = ~G6968 | ~G6971;
  assign G7031 = ~G7026 | ~G7029;
  assign G5521 = ~G5515;
  assign G1756 = ~G5515 | ~G5522;
  assign G5579 = ~G5573;
  assign G1761 = ~G5573 | ~G5580;
  assign G5071 = ~G5069 | ~G5070;
  assign G5159 = ~G5157 | ~G5158;
  assign G5641 = ~G5639 | ~G5640;
  assign G5729 = ~G5727 | ~G5728;
  assign G6107 = ~G6105 | ~G6106;
  assign G6165 = ~G6163 | ~G6164;
  assign G6223 = ~G6221 | ~G6222;
  assign G6317 = ~G6311;
  assign G6320 = ~G6311 | ~G6318;
  assign G6975 = ~G6973 | ~G6974;
  assign G7033 = ~G7031 | ~G7032;
  assign G7097 = ~G7091;
  assign G7100 = ~G7091 | ~G7098;
  assign G7185 = ~G7179;
  assign G7188 = ~G7179 | ~G7186;
  assign G1755 = ~G5518 | ~G5521;
  assign G1760 = ~G5576 | ~G5579;
  assign G6319 = ~G6314 | ~G6317;
  assign G7099 = ~G7094 | ~G7097;
  assign G7187 = ~G7182 | ~G7185;
  assign G1757 = ~G1755 | ~G1756;
  assign G1762 = ~G1760 | ~G1761;
  assign G6113 = ~G6107;
  assign G2818 = ~G6107 | ~G6114;
  assign G6171 = ~G6165;
  assign G2823 = ~G6165 | ~G6172;
  assign G6981 = ~G6975;
  assign G4058 = ~G6975 | ~G6982;
  assign G7039 = ~G7033;
  assign G4063 = ~G7033 | ~G7040;
  assign G5077 = ~G5071;
  assign G5080 = ~G5071 | ~G5078;
  assign G5165 = ~G5159;
  assign G5090 = ~G5159 | ~G5166;
  assign G5647 = ~G5641;
  assign G5650 = ~G5641 | ~G5648;
  assign G5735 = ~G5729;
  assign G5660 = ~G5729 | ~G5736;
  assign G6229 = ~G6223;
  assign G6232 = ~G6223 | ~G6230;
  assign G6321 = ~G6319 | ~G6320;
  assign G7101 = ~G7099 | ~G7100;
  assign G7189 = ~G7187 | ~G7188;
  assign G2817 = ~G6110 | ~G6113;
  assign G2822 = ~G6168 | ~G6171;
  assign G4057 = ~G6978 | ~G6981;
  assign G4062 = ~G7036 | ~G7039;
  assign G5079 = ~G5074 | ~G5077;
  assign G5089 = ~G5162 | ~G5165;
  assign G5649 = ~G5644 | ~G5647;
  assign G5659 = ~G5732 | ~G5735;
  assign G6231 = ~G6226 | ~G6229;
  assign G1782 = G1771 & G1762 & G1730;
  assign G1783 = G1771 & G1757 & G1726;
  assign G1784 = G1766 & G1762 & G1751;
  assign G1785 = G1766 & G1757 & G1754;
  assign G2819 = ~G2817 | ~G2818;
  assign G2824 = ~G2822 | ~G2823;
  assign G4059 = ~G4057 | ~G4058;
  assign G4064 = ~G4062 | ~G4063;
  assign G5081 = ~G5079 | ~G5080;
  assign G5091 = ~G5089 | ~G5090;
  assign G5651 = ~G5649 | ~G5650;
  assign G5661 = ~G5659 | ~G5660;
  assign G6233 = ~G6231 | ~G6232;
  assign G6327 = ~G6321;
  assign G6252 = ~G6321 | ~G6328;
  assign G7107 = ~G7101;
  assign G7110 = ~G7101 | ~G7108;
  assign G7195 = ~G7189;
  assign G7120 = ~G7189 | ~G7196;
  assign G5737 = G1785 | G1784 | G1782 | G1783;
  assign G6251 = ~G6324 | ~G6327;
  assign G7109 = ~G7104 | ~G7107;
  assign G7119 = ~G7192 | ~G7195;
  assign G5087 = ~G5081;
  assign G985 = ~G5081 | ~G5088;
  assign G5097 = ~G5091;
  assign G988 = ~G5091 | ~G5098;
  assign G5657 = ~G5651;
  assign G1776 = ~G5651 | ~G5658;
  assign G5667 = ~G5661;
  assign G1779 = ~G5661 | ~G5668;
  assign G2844 = G2833 & G2824 & G2784;
  assign G2845 = G2833 & G2819 & G2780;
  assign G2846 = G2828 & G2824 & G2813;
  assign G2847 = G2828 & G2819 & G2816;
  assign G4083 = G4072 & G4064 & G4032;
  assign G4084 = G4072 & G4059 & G4028;
  assign G4085 = G4067 & G4064 & G4053;
  assign G4086 = G4067 & G4059 & G4056;
  assign G6239 = ~G6233;
  assign G6242 = ~G6233 | ~G6240;
  assign G6253 = ~G6251 | ~G6252;
  assign G7111 = ~G7109 | ~G7110;
  assign G7121 = ~G7119 | ~G7120;
  assign G984 = ~G5084 | ~G5087;
  assign G987 = ~G5094 | ~G5097;
  assign G1775 = ~G5654 | ~G5657;
  assign G1778 = ~G5664 | ~G5667;
  assign G5743 = ~G5737;
  assign G6241 = ~G6236 | ~G6239;
  assign G6329 = G2847 | G2846 | G2844 | G2845;
  assign G7197 = G4086 | G4085 | G4083 | G4084;
  assign G986 = ~G984 | ~G985;
  assign G989 = ~G987 | ~G988;
  assign G1777 = ~G1775 | ~G1776;
  assign G1780 = ~G1778 | ~G1779;
  assign G6259 = ~G6253;
  assign G2841 = ~G6253 | ~G6260;
  assign G7117 = ~G7111;
  assign G4077 = ~G7111 | ~G7118;
  assign G7127 = ~G7121;
  assign G4080 = ~G7121 | ~G7128;
  assign G6243 = ~G6241 | ~G6242;
  assign G990 = ~G989;
  assign G996 = G975 & G986;
  assign G1781 = ~G1780;
  assign G1787 = G1766 & G1777;
  assign G2840 = ~G6256 | ~G6259;
  assign G6335 = ~G6329;
  assign G4076 = ~G7114 | ~G7117;
  assign G4079 = ~G7124 | ~G7127;
  assign G7203 = ~G7197;
  assign G995 = G990 & G980;
  assign G1786 = G1781 & G1771;
  assign G6249 = ~G6243;
  assign G2838 = ~G6243 | ~G6250;
  assign G2842 = ~G2840 | ~G2841;
  assign G4078 = ~G4076 | ~G4077;
  assign G4081 = ~G4079 | ~G4080;
  assign G2837 = ~G6246 | ~G6249;
  assign G2843 = ~G2842;
  assign G4082 = ~G4081;
  assign G4088 = G4067 & G4078;
  assign G5170 = G995 | G996;
  assign G5740 = G1786 | G1787;
  assign G2839 = ~G2837 | ~G2838;
  assign G2848 = G2843 & G2833;
  assign G4087 = G4082 & G4072;
  assign G1791 = ~G5740 | ~G5743;
  assign G1003 = ~G5170 | ~G5173;
  assign G5174 = ~G5170;
  assign G5744 = ~G5740;
  assign G2849 = G2828 & G2839;
  assign G7200 = G4087 | G4088;
  assign G1792 = ~G5737 | ~G5744;
  assign G1004 = ~G5167 | ~G5174;
  assign G6332 = G2848 | G2849;
  assign G320 = ~G1791 | ~G1792;
  assign G337 = ~G1003 | ~G1004;
  assign G4092 = ~G7200 | ~G7203;
  assign G7204 = ~G7200;
  assign G321 = ~G320;
  assign G338 = ~G337;
  assign G4093 = ~G7197 | ~G7204;
  assign G2855 = ~G6332 | ~G6335;
  assign G6336 = ~G6332;
  assign G369 = ~G4092 | ~G4093;
  assign G2856 = ~G6329 | ~G6336;
  assign G370 = ~G369;
  assign G398 = ~G2855 | ~G2856;
  assign G399 = ~G398;
endmodule


