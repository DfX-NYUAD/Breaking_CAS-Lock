// Benchmark "b21_C_lock" written by ABC on Thu May 13 23:37:50 2021

module b21_C_lock ( 
    keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
    keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
    keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
    keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
    keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
    keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
    keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
    keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
    keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
    keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
    keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
    keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
    keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
    keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
    keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
    keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
    keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
    keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
    keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
    keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
    keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
    keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
    keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
    keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
    keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
    keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
    keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
    keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
    keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
    keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
    keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
    keyinput_156, keyinput_157, keyinput_158, keyinput_159, SI_31_, SI_30_,
    SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
    SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_,
    SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_,
    SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
    P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
    P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
    P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
    P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
    P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
    P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
    P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
    P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
    P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
    P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
    P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
    P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
    P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
    P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
    P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
    P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
    P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
    P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
    P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
    P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
    P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
    P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
    P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
    P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
    P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
    P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
    P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
    P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
    P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
    P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
    P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
    P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
    P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
    P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
    P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
    P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
    P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
    P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
    P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
    P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
    P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
    P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
    P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
    P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
    P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
    P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
    P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
    P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
    P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
    P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
    P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
    P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
    P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
    P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
    P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
    P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
    P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
    P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
    P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
    P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN,
    P1_U3240  );
  input  keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4,
    keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9,
    keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14,
    keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19,
    keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24,
    keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29,
    keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34,
    keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39,
    keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44,
    keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49,
    keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54,
    keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59,
    keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64,
    keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69,
    keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74,
    keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79,
    keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84,
    keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89,
    keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94,
    keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99,
    keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104,
    keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109,
    keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114,
    keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119,
    keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124,
    keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129,
    keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134,
    keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139,
    keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144,
    keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149,
    keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154,
    keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159,
    SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_,
    SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_,
    SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_,
    SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN,
    P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
    P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
    P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
    P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
    P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
    P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
    P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
    P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
    P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN,
    P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
    P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
    P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
    P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
    P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
    P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
    P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
    P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
    P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
    P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
    P1_IR_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
    P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
    P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
    P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN;
  output P1_U3240;
  wire n14461, n9338, n7293, n8118, n7294, n7642, n11962, n11767, n12016,
    n12123, n12384, n8432, n14621, n8411, n14937, n7300, n9339, n7696,
    n7533, n7796, n7422, n7479, n14700, n7494, n14752, n7646, n7647,
    n14758, n9601, n7706, n14976, n14942, n8304, n10535, n10531, n7435,
    n7438, n7877, n7867, n7883, n7898, n7500, n14654, n14690, n7490, n7491,
    n7492, n7493, n7484, n7485, n7483, n7504, n7505, n14751, n14812, n7425,
    n7423, n14786, n14701, n14913, n14777, n14803, n14770, n14888, n14631,
    n11843, n7849, n7535, n7813, n7811, n8153, n7600, n7601, n7310, n7693,
    n7694, n14925, n14884, n13776, n14863, n14958, n7445, n8302, n8278,
    n7427, n7429, n7638, n8048, n8236, n7630, n7807, n7804, n7446, n7949,
    n7831, n12873, n10170, n12680, n14897, n8389, n10992, n14797, n14994,
    n14193, n14980, n13833, n14644, n14974, n8890, n7967, n10530, n7532,
    n8375, n14612, n13400, n8266, n15007, n14939, n8151, n7499, n14662,
    n7489, n7498, n14723, n14750, n14804, n7440, n7432, n7433, n7434,
    n7439, n7436, n7437, n7430, n7428, n7707, n7534, n7851, n7850, n7822,
    n7821, n7453, n7511, n7512, n7645, n7631, n7424, n7506, n7634, n7641,
    n7720, n7856, n7905, n7923, n7944, n7962, n7643, n7644, n7996, n8030,
    n8223, n8203, n14914, n14449, n14998, n14743, n14972, n11906, n7531,
    n8394, n7895, n7448, n8248, n7695, n7853, n7854, n8230, n7697, n7817,
    n7816, n7819, n8189, n11299, n14132, n10706, n7603, n10225, n7480,
    n12364, n12365, n9549, n7692, n10772, n9590, n9579, n11766, n14905,
    n7447, n10691, n10267, n10166, n8307, n14419, n14336, n7648, n8270,
    n14978, n13212, n14962, n12820, n12184, n12156, n14025, n14230, n13608,
    n13200, n13175, n12804, n12638, n7866, n8355, n8337, n7443, n8335,
    n8320, n8291, n7637, n8019, n7421, n8214, n8216, n8096, n7442, n11330,
    n13821, n7452, n13523, n13223, n12982, n12626, n7502, n7501, n8080,
    n14940, n13683, n13387, n14462, n9332, n13698, n13408, n13139, n13085,
    n7649, n12896, n12733, n9265, n15005, n7632, n7507, n7301, n7305,
    n7308, n7309, n7311, n14744, n7314, n7319, n7322, n7878, n7327, n7330,
    n7335, n7336, n7338, n7345, n7346, n7347, n14628, n7352, n7358, n7359,
    n7360, n7366, n7367, n7369, n7370, n15000, n7657, n7513, n7374, n7377,
    n7381, n8105, n14634, n7386, n7848, n7389, n7391, n7394, n7396, n7397,
    n7398, n7399, n7400, n7405, n8170, n7426, n8003, n7431, n9343, n7441,
    n7444, n10536, n7913, n7449, n7450, n7451, n7508, n7510, n11182, n7454,
    n7477, n7478, n14795, n7481, n7482, n14946, n7486, n14693, n7487,
    n7488, n14699, n7495, n7496, n7497, n7868, n10886, n7652, n7503,
    n14739, n14736, n12008, n14727, n14657, n7629, n7509, n7865, n11097,
    n11997, n7951, n7608, n8004, n7628, n8171, n8245, n7633, n7635, n7636,
    n7931, n7639, n7640, n7986, n7650, n7651, P1_U3240_Lock, n7653, n7654,
    n7655, n7789, n7656, n8060, n14788, n8410, n11768, n14694, n14724,
    n14653, n14703, n14696, n7855, n7852, n7726, n7769, n8324, n8294,
    n8256, n7982, n8039, n8416, n7771, n9328, n8362, n8282, n7887, n8012,
    n11378, n11963, n14616, n9996, n7728, n7727, n8319, n8321, n7730,
    n7729, n7731, n7847, n8303, n7733, n7732, n7734, n7845, n8292, n7736,
    n7735, n7737, n7843, n8279, n7739, n7738, n7740, n8267, n7742, n7741,
    n7743, n7841, n7884, n7745, n7744, n7746, n7840, n7896, n7748, n7747,
    n7749, n7838, n7914, n7751, n7750, n7752, n7837, n8246, n7754, n7753,
    n7755, n7836, n7932, n7757, n7756, n7833, n7835, n7759, n7758, n7830,
    n7832, n7761, n7760, n7762, n7829, n7987, n7764, n7763, n7826, n7828,
    n7766, n7765, n7767, n7825, n8020, n7768, n7824, n7770, n8046, n7772,
    n7775, n7773, n7774, n7776, n7783, n11084, n8688, n7777, n7781, n8068,
    n7778, n7779, n7780, n7782, n11127, n7785, n7784, n7787, n7786, n8095,
    n7788, n8116, n10996, n7791, n7790, n7793, n7792, n8114, n7795, n7794,
    n8132, n11078, n7798, n7797, n7800, n7799, n8130, n7802, n7801, n8152,
    n7803, n7805, n9183, n7806, n7808, n7809, n11196, n7810, n7812, n8197,
    n7814, n7815, n7818, n8213, n7820, n8234, n7823, n8002, n7827, n7968,
    n7948, n7834, n7839, n7842, n7844, n7846, n13315, n9307, n7858, n7857,
    n7860, n7859, n7861, n9330, n8059, n7863, n8188, n8049, n9308, n7862,
    n7864, n8165, n8164, n8181, n10172, n7869, n7872, n7870, n7871, n7873,
    n7874, n8109, n7882, n8220, n7876, n8069, n7875, n7880, n9345, n8180,
    n7879, n7881, n11341, n10031, n14805, n14761, n14813, n14992, n12549,
    n7886, n9266, n7885, n14222, n7888, n7894, n7890, n7889, n7892, n7891,
    n7893, n13861, n14881, n12493, n8977, n7904, n7897, n7902, n7899,
    n7900, n7901, n7903, n14126, n7906, n7912, n8380, n7908, n7907, n7910,
    n7909, n7911, n13944, n14638, n12280, n8959, n7922, n7915, n7920,
    n7916, n7917, n8249, n8251, n7918, n14098, n14092, n7919, n7921,
    n14068, n7930, n7925, n7924, n7928, n7926, n7927, n7929, n13862,
    n14729, n14982, n11893, n8922, n7938, n7933, n7936, n8229, n7934,
    n13639, n13630, n7935, n7937, n7940, n7939, n7943, n7941, n7942, n7946,
    n13816, n7945, n13591, n7947, n14714, n14821, n11782, n8905, n7956,
    n7950, n7954, n7952, n13152, n13143, n7953, n7955, n7958, n7957, n7961,
    n7959, n7960, n7964, n13486, n7963, n13661, n7965, n14823, n14855,
    n7966, n7977, n7969, n7975, n7970, n7989, n7971, n7972, n7973, n12852,
    n12399, n7974, n7976, n7979, n7978, n7981, n7980, n7984, n13551, n7983,
    n13221, n7985, n14706, n14858, n14853, n11592, n8851, n7993, n7988,
    n7991, n12400, n12393, n7990, n7992, n7995, n7994, n8001, n7999,
    n13321, n7997, n7998, n8000, n8037, n8038, n11538, n8009, n11530,
    n8007, n8005, n11949, n11939, n8006, n8008, n8011, n8010, n8017, n8015,
    n13194, n8013, n8014, n8016, n8018, n14702, n14698, n11374, n8027,
    n11366, n8025, n8021, n8022, n8052, n8051, n8054, n8023, n11615,
    n11622, n8024, n8026, n8029, n8028, n8035, n8033, n13206, n8031, n8032,
    n8034, n8490, n8036, n14645, n14852, n13331, n8041, n12872, n8040,
    n8045, n8043, n8042, n8044, n8047, n11377, n8058, n8050, n8056, n8053,
    n11515, n11384, n8055, n8057, n14868, n8061, n11001, n8067, n8062,
    n8065, n8063, n8064, n8066, n11152, n11022, n8071, n8070, n8075, n8073,
    n8072, n8074, n8088, n8086, n8077, n8076, n8081, n8079, n8078, n8085,
    n9562, n8084, n8082, n10942, n8083, n12357, n8087, n8103, n8090, n8089,
    n8094, n8092, n8091, n8093, n8097, n11125, n8100, n8098, n11025,
    n11393, n8099, n8102, n9161, n8101, n12017, n8104, n8472, n14831,
    n8107, n8106, n8113, n8111, n8108, n8110, n8112, n8115, n10984, n8121,
    n8117, n8119, n8134, n8133, n11052, n10985, n8120, n8124, n8122, n8123,
    n14871, n11920, n12178, n14917, n14944, n11971, n8125, n8127, n8126,
    n12227, n8128, n8129, n8131, n11076, n8138, n8135, n8136, n11051,
    n11441, n8137, n8140, n9156, n8139, n12236, n14832, n8142, n8141,
    n8150, n8148, n8144, n8143, n8145, n12261, n8146, n8147, n8149, n9171,
    n8159, n8154, n8156, n8155, n8157, n11140, n11060, n8158, n8161, n9172,
    n8160, n14833, n11919, n12269, n14672, n14947, n8163, n8162, n8169,
    n8166, n12216, n8167, n8168, n9182, n8174, n8172, n11112, n11105,
    n8173, n8176, n9177, n8175, n14671, n12197, n12221, n14673, n14953,
    n14835, n8179, n8178, n8186, n8184, n12815, n8182, n8183, n8185, n8187,
    n8196, n8190, n8191, n8194, n8193, n8192, n8209, n11260, n11252, n8195,
    n8200, n8198, n8199, n14650, n9197, n12771, n14676, n8202, n8201,
    n8208, n8206, n12521, n8204, n8205, n8207, n8482, n11293, n8212, n8210,
    n11275, n11294, n8211, n8218, n8215, n11302, n8217, n12556, n14666,
    n12377, n14840, n8222, n8221, n8227, n8225, n12679, n8224, n8226,
    n8228, n8233, n8231, n11311, n11336, n8232, n8238, n8235, n11329,
    n8237, n14825, n14683, n14692, n14846, n8491, n14646, n12977, n8242,
    n8241, n8493, n14967, n14851, n12128, n8941, n8255, n8247, n8253,
    n8250, n13888, n13638, n8252, n8254, n13832, n8263, n8258, n8257,
    n8261, n8259, n8260, n8262, n13757, n8264, n14715, n14822, n14639,
    n14637, n14878, n12736, n8269, n12730, n8268, n14003, n9794, n8276,
    n8272, n8271, n8274, n8273, n8275, n13942, n14633, n12899, n8281,
    n12893, n8280, n14188, n9862, n8288, n8284, n8283, n8286, n8285, n8287,
    n11166, n8289, n14816, n14632, n14988, n13083, n8293, n14259, n10087,
    n8300, n8296, n8295, n8298, n8297, n8299, n11272, n14740, n14748,
    n13186, n8306, n13136, n8305, n14414, n10148, n8313, n8309, n8308,
    n8311, n8310, n8312, n11323, n8314, n8315, n14424, n14990, n8318,
    n8317, n8334, n8336, n13456, n8323, n13403, n8322, n8342, n10227,
    n8330, n8326, n8325, n8328, n8327, n8329, n11326, n8331, n14806, n8333,
    n8332, n8354, n8356, n8338, n8340, n9313, n8339, n8341, n8363, n10295,
    n8348, n8344, n8343, n8346, n8345, n8347, n11527, n10032, n8351, n8358,
    n8357, n8360, n8359, n8373, n8374, n9317, n8361, n8379, n10708, n8369,
    n8365, n8364, n8367, n8366, n8368, n11635, n10698, n14622, n14802,
    n8372, n8371, n9344, n9342, n8376, n9322, n8378, n9333, n8377, n8540,
    n8386, n8382, n8381, n8384, n8383, n8385, n11570, n8387, n8392, n8533,
    n8390, n15009, n14903, n8391, n8393, n8395, n9779, n13222, n14614,
    n8400, n8399, n8403, n8401, n8402, n14798, n8434, n8421, n8412, n8413,
    n8414, n8415, n8431, n8430, n8420, n8422, n8423, n8424, n9791, n8433,
    n13082, n8435, n9785, n14611, n11671, n10752, n11670, n14943, n12748,
    n12747, n13171, n13939, n13081, n9341, n9340, n10532, n14450, n12015,
    n10534, n10533, n10541, n10538, n10537, n10539, n10540, n14463, n11188,
    n11187, n11191, n11189, n11190, n14780, n14950, n14916, n14951, n14839,
    n14960, n12749, n14964, n14689, n14902, n14966, n14968, n13934, n14984,
    n14451, n14465, n14464, n14613, n14615, n14620, n15012, n14794, n14618,
    n14617, n14619, n14896, n14934, n14799, n15004, n14792, n14783, n14625,
    n14623, n14624, n14771, n14630, n14626, n14627, n14629, n14776, n14738,
    n14880, n14636, n14817, n14635, n14746, n14735, n14730, n14641, n14731,
    n14640, n14728, n14642, n14643, n14713, n14849, n14697, n14648, n14647,
    n14649, n14651, n14842, n14652, n14665, n14663, n14656, n14829, n14655,
    n14661, n14659, n14675, n14658, n14660, n14664, n14669, n14667, n14670,
    n14668, n14682, n14680, n14674, n14827, n14677, n14826, n14678, n14679,
    n14681, n14686, n14684, n14685, n14687, n14688, n14695, n14691, n14711,
    n14705, n14704, n14707, n14709, n14708, n14710, n14712, n14824, n14718,
    n14717, n14876, n14716, n14720, n14719, n14721, n14722, n14726, n14725,
    n14745, n14875, n14732, n14733, n14734, n14737, n14742, n14741, n14983,
    n14747, n14749, n14820, n14754, n14753, n14757, n14755, n14756, n14768,
    n14763, n14759, n14760, n14762, n14766, n14764, n14765, n14767, n14769,
    n14774, n14889, n14772, n14773, n14775, n14779, n14778, n14941, n14781,
    n14787, n14782, n14785, n14784, n14791, n14789, n14790, n14793, n14796,
    n14901, n14801, n14800, n14895, n14893, n14814, n14809, n14807, n14808,
    n14810, n14811, n14907, n14815, n14926, n14818, n14819, n14912, n14862,
    n14866, n14860, n14828, n14864, n14830, n14837, n14834, n14836, n14838,
    n14844, n14841, n14843, n14845, n14847, n14848, n14850, n14854, n14870,
    n14856, n14857, n14859, n14861, n14874, n14865, n14867, n14869, n14908,
    n14872, n14873, n14879, n14877, n14909, n14883, n14882, n14885, n14886,
    n14887, n14923, n14890, n14891, n14892, n14894, n14899, n14936, n14898,
    n14900, n14904, n14932, n14906, n14930, n14910, n14911, n14921, n14915,
    n14919, n14918, n14920, n14922, n14924, n14928, n14927, n14929, n14931,
    n14933, n14935, n14938, n15002, n14996, n14945, n14949, n14948, n14956,
    n14952, n14954, n14955, n14957, n14959, n14961, n14963, n14965, n14970,
    n14969, n14971, n14973, n14975, n14977, n14979, n14981, n14986, n14985,
    n14987, n14989, n14991, n14993, n14995, n14997, n14999, n15001, n15003,
    n15006, n15008, n15010, n15011, input_0, input_1, AND_1, input_2, OR_2,
    input_3, AND_3, input_4, OR_4, input_5, AND_5, input_6, AND_6, input_7,
    OR_7, input_8, AND_8, input_9, OR_9, input_10, AND_10, input_11, OR_11,
    input_12, AND_12, input_13, OR_13, input_14, AND_14, input_15, OR_15,
    input_16, OR_16, input_17, OR_17, input_18, AND_18, input_19, OR_19,
    input_20, OR_20, input_21, OR_21, input_22, AND_22, input_23, OR_23,
    input_24, OR_24, input_25, AND_25, input_26, AND_26, input_27, OR_27,
    input_28, OR_28, input_29, AND_29, input_30, AND_30, input_31, AND_31,
    input_32, OR_32, input_33, AND_33, input_34, AND_34, input_35, OR_35,
    input_36, AND_36, input_37, OR_37, input_38, OR_38, input_39, AND_39,
    input_40, AND_40, input_41, AND_41, input_42, OR_42, input_43, OR_43,
    input_44, AND_44, input_45, OR_45, input_46, OR_46, input_47, OR_47,
    input_48, OR_48, input_49, AND_49, input_50, AND_50, input_51, OR_51,
    input_52, OR_52, input_53, AND_53, input_54, OR_54, input_55, OR_55,
    input_56, AND_56, input_57, OR_57, input_58, AND_58, input_59, OR_59,
    input_60, OR_60, input_61, AND_61, input_62, OR_62, input_63, AND_63,
    input_64, AND_64, input_65, AND_65, input_66, OR_66, input_67, AND_67,
    input_68, AND_68, input_69, OR_69, input_70, OR_70, input_71, AND_71,
    input_72, AND_72, input_73, AND_73, input_74, OR_74, input_75, AND_75,
    input_76, AND_76, input_77, OR_77, input_78, AND_78, input_79, AND_79,
    input_80, input_81, AND_81, input_82, OR_82, input_83, AND_83,
    input_84, OR_84, input_85, AND_85, input_86, AND_86, input_87, OR_87,
    input_88, AND_88, input_89, OR_89, input_90, AND_90, input_91, OR_91,
    input_92, AND_92, input_93, OR_93, input_94, AND_94, input_95, OR_95,
    input_96, OR_96, input_97, OR_97, input_98, AND_98, input_99, OR_99,
    input_100, OR_100, input_101, OR_101, input_102, AND_102, input_103,
    OR_103, input_104, OR_104, input_105, AND_105, input_106, AND_106,
    input_107, OR_107, input_108, OR_108, input_109, AND_109, input_110,
    AND_110, input_111, AND_111, input_112, OR_112, input_113, AND_113,
    input_114, AND_114, input_115, OR_115, input_116, AND_116, input_117,
    OR_117, input_118, OR_118, input_119, AND_119, input_120, AND_120,
    input_121, AND_121, input_122, OR_122, input_123, OR_123, input_124,
    AND_124, input_125, OR_125, input_126, OR_126, input_127, OR_127,
    input_128, OR_128, input_129, AND_129, input_130, AND_130, input_131,
    OR_131, input_132, OR_132, input_133, AND_133, input_134, OR_134,
    input_135, OR_135, input_136, AND_136, input_137, OR_137, input_138,
    AND_138, input_139, OR_139, input_140, OR_140, input_141, AND_141,
    input_142, OR_142, input_143, AND_143, input_144, AND_144, input_145,
    AND_145, input_146, OR_146, input_147, AND_147, input_148, AND_148,
    input_149, OR_149, input_150, OR_150, input_151, AND_151, input_152,
    AND_152, input_153, AND_153, input_154, OR_154, input_155, AND_155,
    input_156, AND_156, input_157, OR_157, input_158, AND_158, input_159,
    AND_159, AND_159_INV, CASOP;
  assign n14461 = ~n8059;
  assign n9338 = ~n7796;
  assign n7293 = ~n7300 | ~n7381;
  assign n8118 = ~P1_IR_REG_1__SCAN_IN & ~P1_IR_REG_0__SCAN_IN;
  assign n7294 = ~n8069;
  assign n7642 = ~n7640 | ~n7643;
  assign n11962 = ~n7501 | ~n7502;
  assign n11767 = n8081 | n8080;
  assign n12016 = ~n11997;
  assign n12123 = ~n12236;
  assign n12384 = n8102 | n8101;
  assign n8432 = n8431 & n8430;
  assign n14621 = ~n8395 ^ n8394;
  assign n8411 = n8410 | P1_IR_REG_21__SCAN_IN;
  assign n14937 = ~n7900 ^ P1_IR_REG_19__SCAN_IN;
  assign n7300 = ~n7898;
  assign n9339 = ~n9338;
  assign n7696 = n7852 & n7533;
  assign n7533 = n7534 & n7535;
  assign n7796 = ~n7424 | ~n7422;
  assign n7422 = ~n7423 | ~n7506;
  assign n7479 = n7695 & n7696;
  assign n14700 = n14699 & n14783;
  assign n7494 = ~n14853;
  assign n14752 = n14742 | n14741;
  assign n7646 = ~n8234 & ~n7647;
  assign n7647 = ~n7819;
  assign n14758 = n14419 | n8314;
  assign n9601 = ~n11962;
  assign n7706 = n7707 & n8394;
  assign n14976 = n14714 & n14821;
  assign n14942 = n14622 & n14802;
  assign n8304 = ~n8049;
  assign n10535 = ~n7796;
  assign n10531 = ~n7438 | ~n7435;
  assign n7435 = ~n7436 & ~n7399;
  assign n7438 = ~n8375 | ~n7439;
  assign n7877 = ~n7867 ^ P1_IR_REG_30__SCAN_IN;
  assign n7867 = ~n10886 | ~P1_IR_REG_31__SCAN_IN;
  assign n7883 = ~n7840 | ~n7839;
  assign n7898 = ~n7479 | ~n7358;
  assign n7500 = ~n7865;
  assign n14654 = ~n14944 & ~n14831;
  assign n14690 = n14682 & n14681;
  assign n7490 = ~n14691;
  assign n7491 = ~n7493 & ~n7492;
  assign n7492 = ~n14692;
  assign n7493 = n14691 & n14689;
  assign n7484 = ~n14712 | ~n7485;
  assign n7485 = n14713 & n7346;
  assign n7483 = n14719 & n7345;
  assign n7504 = ~n14745 | ~n7505;
  assign n7505 = ~n14878;
  assign n14751 = ~n14888 & ~n14750;
  assign n14812 = n14449 & n8387;
  assign n7425 = ~P1_ADDR_REG_19__SCAN_IN & ~P1_RD_REG_SCAN_IN;
  assign n7423 = P2_ADDR_REG_19__SCAN_IN & P1_ADDR_REG_19__SCAN_IN;
  assign n14786 = n7477 & n7370;
  assign n14701 = n13387 | n13523;
  assign n14913 = ~n11766 & ~n11997;
  assign n14777 = ~n14812;
  assign n14803 = n14449 | n8387;
  assign n14770 = ~n10267 & ~n10032;
  assign n14888 = n14419 & n8314;
  assign n14631 = n14025 | n13942;
  assign n11843 = n7486 & n14863;
  assign n7849 = ~P1_IR_REG_8__SCAN_IN;
  assign n7535 = ~P1_IR_REG_6__SCAN_IN & ~P1_IR_REG_7__SCAN_IN;
  assign n7813 = ~n7811 | ~n7810;
  assign n7811 = n9339 | n11196;
  assign n8153 = ~n7600 | ~n8118;
  assign n7600 = n7601 & n8133;
  assign n7601 = ~P1_IR_REG_2__SCAN_IN & ~P1_IR_REG_4__SCAN_IN;
  assign n7310 = n8061 & n11001;
  assign n7693 = n7878 | n7694;
  assign n7694 = ~P1_REG0_REG_6__SCAN_IN;
  assign n14925 = n10225 | n8331;
  assign n14884 = ~n14336 & ~n11272;
  assign n13776 = n7922 & n7921;
  assign n14863 = ~n11962 | ~n12123;
  assign n14958 = n14650 & n14676;
  assign n7445 = ~n8321;
  assign n8302 = ~n7845 | ~n7844;
  assign n8278 = ~n7429 | ~n7427;
  assign n7427 = ~n7428 & ~n7394;
  assign n7429 = ~n7883 | ~n7430;
  assign n7638 = n7932 & n7639;
  assign n8048 = ~n7509 | ~n7338;
  assign n8236 = ~n8216 | ~n7819;
  assign n7630 = n7631 & n7809;
  assign n7807 = n9339 | n9183;
  assign n7804 = ~n7803 | ~n7446;
  assign n7446 = ~n9338 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n7949 = ~n7832 & ~n7831;
  assign n7831 = n7642 & n7391;
  assign n12873 = ~n12804;
  assign n10170 = ~n10166;
  assign n12680 = ~n12638;
  assign n14897 = n14621 | n14937;
  assign n8389 = ~n7300 | ~n7720;
  assign n10992 = ~n8045 & ~n8044;
  assign n14797 = ~n14465 | ~n14464;
  assign n14994 = n14925 & n14806;
  assign n14193 = ~n8281 | ~n8280;
  assign n14980 = n14715 & n14822;
  assign n13833 = ~n8255 | ~n8254;
  assign n14644 = ~n14976;
  assign n14974 = n7966 | n14823;
  assign n8890 = ~n7967 ^ n7968;
  assign n7967 = ~n7642 | ~n7829;
  assign n10530 = n10532 ^ n10531;
  assign n7532 = ~n7865 | ~P1_IR_REG_31__SCAN_IN;
  assign n8375 = ~n8358 | ~n8357;
  assign n14612 = ~n7861 ^ P1_IR_REG_27__SCAN_IN;
  assign n13400 = ~n8424 ^ P1_IR_REG_26__SCAN_IN;
  assign n8266 = ~n7431 | ~n7841;
  assign n15007 = ~n8533;
  assign n14939 = ~n15009;
  assign n8151 = ~n7804 ^ SI_5_;
  assign n7499 = n7866 & n7870;
  assign n14662 = ~n14661 & ~n14660;
  assign n7489 = ~n7327 & ~n14792;
  assign n7498 = ~n14703;
  assign n14723 = ~n7484 | ~n7483;
  assign n14750 = n7650 & n14783;
  assign n14804 = ~n14623 & ~n14628;
  assign n7440 = ~n7441 | ~n9342;
  assign n7432 = ~n7433 | ~n8267;
  assign n7433 = ~n7434 | ~n7841;
  assign n7434 = ~n7884;
  assign n7439 = ~n7440;
  assign n7436 = ~n7440 & ~n7437;
  assign n7437 = ~n8374;
  assign n7430 = ~n7432;
  assign n7428 = ~n7432 & ~n7841;
  assign n7707 = ~P1_IR_REG_20__SCAN_IN;
  assign n7534 = n7849 & n7848;
  assign n7851 = ~P1_IR_REG_9__SCAN_IN & ~P1_IR_REG_10__SCAN_IN;
  assign n7850 = ~P1_IR_REG_11__SCAN_IN;
  assign n7822 = ~n7821 | ~n7820;
  assign n7821 = n10536 | n11330;
  assign n7453 = ~n7454;
  assign n7511 = n7646 & n7512;
  assign n7512 = n8197 | n7513;
  assign n7645 = ~n7646 | ~n8213;
  assign n7631 = n7805 | n8170;
  assign n7424 = ~n7425 | ~n7726;
  assign n7506 = ~P2_RD_REG_SCAN_IN;
  assign n7634 = n7638 | n7635;
  assign n7641 = ~n7968;
  assign n7720 = n8248 & n7856;
  assign n7856 = ~P1_IR_REG_19__SCAN_IN;
  assign n7905 = n7923 & P1_REG3_REG_18__SCAN_IN;
  assign n7923 = n8256 & P1_REG3_REG_17__SCAN_IN;
  assign n7944 = n7962 & P1_REG3_REG_15__SCAN_IN;
  assign n7962 = n7982 & P1_REG3_REG_14__SCAN_IN;
  assign n7643 = ~n7828 & ~n7644;
  assign n7644 = ~n7987;
  assign n7996 = n8012 & P1_REG3_REG_12__SCAN_IN;
  assign n8030 = n8039 & P1_REG3_REG_10__SCAN_IN;
  assign n8223 = n8203 & P1_REG3_REG_8__SCAN_IN;
  assign n8203 = n8181 & P1_REG3_REG_7__SCAN_IN;
  assign n14914 = ~n11963 | ~n12017;
  assign n14449 = ~n8378 | ~n8377;
  assign n14998 = ~n14628 & ~n14770;
  assign n14743 = n14631 & n14633;
  assign n14972 = ~n14858 & ~n14853;
  assign n11906 = n8161 | n8160;
  assign n7531 = ~n7301 & ~P1_IR_REG_27__SCAN_IN;
  assign n8394 = ~P1_IR_REG_22__SCAN_IN;
  assign n7895 = ~n7448 | ~n7838;
  assign n7448 = ~n7913 | ~n7914;
  assign n8248 = ~P1_IR_REG_17__SCAN_IN;
  assign n7695 = ~n8153;
  assign n7853 = ~P1_IR_REG_14__SCAN_IN;
  assign n7854 = ~P1_IR_REG_12__SCAN_IN & ~P1_IR_REG_13__SCAN_IN;
  assign n8230 = ~n7697 & ~n8153;
  assign n7697 = ~n7386 | ~n7848;
  assign n7817 = ~n7816 | ~n7815;
  assign n7816 = n10536 | n11299;
  assign n7819 = n7817 | SI_8_;
  assign n8189 = ~n7695 | ~n7848;
  assign n11299 = ~P1_DATAO_REG_8__SCAN_IN;
  assign n14132 = n7904 & n7903;
  assign n10706 = n8362 & n8361;
  assign n7603 = ~n7310 & ~n7330;
  assign n10225 = ~n8323 | ~n8322;
  assign n7480 = n7347 & n14793;
  assign n12364 = ~n8227 & ~n8226;
  assign n12365 = ~n8186 & ~n8185;
  assign n9549 = ~n8169 & ~n7692;
  assign n7692 = ~n8168 | ~n7693;
  assign n10772 = ~n8150 & ~n8149;
  assign n9590 = ~n8113 & ~n8112;
  assign n9579 = ~n8094 & ~n8093;
  assign n11766 = ~n8075 & ~n8074;
  assign n14905 = ~n7447 | ~n14451;
  assign n7447 = ~n7305 | ~n14461;
  assign n10691 = ~n10706;
  assign n10267 = ~n8340 | ~n8339;
  assign n10166 = ~n7863 | ~n7862;
  assign n8307 = n8294 & P1_REG3_REG_23__SCAN_IN;
  assign n14419 = ~n8306 | ~n8305;
  assign n14336 = n7648 & n8293;
  assign n7648 = ~n13085 | ~n14461;
  assign n8270 = n7887 & P1_REG3_REG_20__SCAN_IN;
  assign n14978 = n13939 | n14638;
  assign n13212 = n8027 & n8026;
  assign n14962 = n14666 & n14840;
  assign n12820 = ~n8200 | ~n8199;
  assign n12184 = n8176 | n8175;
  assign n12156 = n8124 | n8123;
  assign n14025 = n8269 & n8268;
  assign n14230 = n7886 & n7885;
  assign n13608 = ~n7956 | ~n7955;
  assign n13200 = n8009 & n8008;
  assign n13175 = ~n13212;
  assign n12804 = n8058 & n8057;
  assign n12638 = n8238 & n8237;
  assign n7866 = ~P1_IR_REG_28__SCAN_IN;
  assign n8355 = ~n8338 | ~n8337;
  assign n8337 = ~n7444 | ~n7443;
  assign n7443 = n8336 & n7400;
  assign n8335 = n7444 & n7400;
  assign n8320 = ~n7846 | ~n7847;
  assign n8291 = ~n7843 | ~n7842;
  assign n7637 = ~n7834;
  assign n8019 = ~n7421 | ~n7824;
  assign n7421 = ~n8048 | ~n8046;
  assign n8214 = ~n7510 | ~n7814;
  assign n8216 = n8214 | n8213;
  assign n8096 = ~n7656 | ~n7783;
  assign n7442 = ~n8375 & ~n8374;
  assign n11330 = ~P1_DATAO_REG_9__SCAN_IN;
  assign n13821 = ~n7938 | ~n7937;
  assign n7452 = n15011 & n14902;
  assign n13523 = n8001 | n8000;
  assign n13223 = n8017 | n8016;
  assign n12982 = n8035 | n8034;
  assign n12626 = n8208 | n8207;
  assign n7502 = ~n8180 | ~P1_REG0_REG_4__SCAN_IN;
  assign n7501 = n7377 & n8129;
  assign n8080 = ~n8079 | ~n8078;
  assign n14940 = ~n14905;
  assign n13683 = ~n7977 | ~n7976;
  assign n13387 = n7993 & n7992;
  assign n14462 = ~n10541 ^ n10540;
  assign n9332 = ~n10886 | ~n7873;
  assign n13698 = ~n8375 ^ n8374;
  assign n13408 = ~n13456;
  assign n13139 = ~n13186;
  assign n13085 = ~n8291 ^ n7649;
  assign n7649 = ~n8292;
  assign n12896 = ~n12899;
  assign n12733 = ~n12736;
  assign n9265 = ~n12549;
  assign n15005 = ~n14937;
  assign n7632 = ~n8152 | ~n7507;
  assign n7507 = ~n8151;
  assign n7301 = ~n7308 | ~n7336;
  assign n7305 = n10530 ^ SI_30_;
  assign n7308 = n7720 & n7706;
  assign n7309 = n8356 ^ n8355;
  assign n7311 = ~n13776 | ~n13862;
  assign n14744 = ~n14748 & ~n14884;
  assign n7314 = n7359 & n7608;
  assign n7319 = n14832 & n14871;
  assign n7322 = n7452 & n7450;
  assign n7878 = ~n8180;
  assign n7327 = n7491 & n7490;
  assign n7330 = ~n9330 & ~n11022;
  assign n7335 = n8188 | n8068;
  assign n7336 = n7860 & n7859;
  assign n7338 = n7645 & n7823;
  assign n7345 = n14821 | n14783;
  assign n7346 = n14855 | n14792;
  assign n7347 = n14896 | n14792;
  assign n14628 = n10267 & n10032;
  assign n7352 = n14747 | n14884;
  assign n7358 = n7314 & n7855;
  assign n7359 = n7854 & n7853;
  assign n7360 = ~n14983 & ~n14881;
  assign n7366 = n14791 & n7482;
  assign n7367 = n7898 | n7301;
  assign n7369 = n14706 & n14701;
  assign n7370 = ~n14779 & ~n14778;
  assign n15000 = ~n14777 | ~n14803;
  assign n7657 = ~n15000;
  assign n7513 = ~n7814;
  assign n7374 = n14863 & n7319;
  assign n7377 = n8127 & n8126;
  assign n7381 = n7720 & n7707;
  assign n8105 = n7877 | n9332;
  assign n14634 = n14193 | n8289;
  assign n7386 = n7535 & n7849;
  assign n7848 = ~P1_IR_REG_5__SCAN_IN;
  assign n7389 = n7634 & n8246;
  assign n7391 = n7641 & n7829;
  assign n7394 = SI_21_ & n7740;
  assign n7396 = n7479 & n7314;
  assign n7397 = n7445 & n7847;
  assign n7398 = n7695 & n7359;
  assign n7399 = SI_29_ & n9344;
  assign n7400 = SI_25_ | n8319;
  assign n7405 = n14620 & n14619;
  assign n8170 = ~n7808 ^ SI_6_;
  assign n7426 = ~n8019 & ~n8020;
  assign n8003 = ~n7426 & ~n7825;
  assign n7431 = ~n7883 | ~n7884;
  assign n9343 = ~n7442 & ~n8376;
  assign n7441 = ~n8376;
  assign n7444 = ~n7846 | ~n7397;
  assign n10536 = ~n9338;
  assign n7913 = ~n7449 | ~n7837;
  assign n7449 = ~n7636 | ~n7389;
  assign n7450 = ~n7451 | ~n14939;
  assign n7451 = ~n14938 ^ n14937;
  assign n7508 = ~n7453 | ~n7814;
  assign n7510 = ~n7454 | ~n8197;
  assign n11182 = ~n7454 ^ n8198;
  assign n7454 = ~n7628 | ~n7630;
  assign n7477 = ~n7478 | ~n7657;
  assign n7478 = ~n14775 | ~n14776;
  assign n14795 = ~n7481 | ~n7480;
  assign n7481 = ~n7366 | ~n14790;
  assign n7482 = ~n15004;
  assign n14946 = ~n14863 | ~n14832;
  assign n7486 = ~n8125 | ~n7374;
  assign n14693 = ~n7487 | ~n7489;
  assign n7487 = ~n7488 | ~n7491;
  assign n7488 = ~n14690;
  assign n14699 = ~n7495 | ~n7494;
  assign n7495 = ~n7496 | ~n7369;
  assign n7496 = ~n7497 | ~n14645;
  assign n7497 = ~n7498 | ~n14851;
  assign n7868 = ~n7500 | ~n7866;
  assign n10886 = ~n7500 | ~n7499;
  assign n7652 = ~n7503 | ~n7352;
  assign n7503 = ~n7360 | ~n7504;
  assign n14739 = ~n14738 & ~n14737;
  assign n14736 = ~n14735 & ~n14734;
  assign n12008 = ~n8088 | ~n8087;
  assign n14727 = ~n14726 & ~n14725;
  assign n14657 = ~n14656 & ~n14655;
  assign n7629 = ~n8170 & ~n8151;
  assign n7509 = ~n7508 | ~n7511;
  assign n7865 = ~n7531 | ~n7300;
  assign n11097 = ~n7532 ^ P1_IR_REG_28__SCAN_IN;
  assign n11997 = ~n7603 | ~n7335;
  assign n7951 = ~n7398 | ~n7696;
  assign n7608 = ~P1_IR_REG_15__SCAN_IN;
  assign n8004 = ~n7696 | ~n7695;
  assign n7628 = ~n7629 | ~n8152;
  assign n8171 = ~n7632 | ~n7805;
  assign n8245 = ~n7633 | ~n7836;
  assign n7633 = ~n7637 | ~n7638;
  assign n7635 = ~n7836;
  assign n7636 = ~n7834 | ~n7836;
  assign n7931 = ~n7834 & ~n7835;
  assign n7639 = ~n7835;
  assign n7640 = ~n7827;
  assign n7986 = ~n7827 & ~n7828;
  assign n7650 = ~n7651 | ~n14820;
  assign n7651 = ~n7652 | ~n14632;
  assign P1_U3240_Lock = ~n7654 | ~n7653;
  assign n7653 = ~n7322 & ~n7405;
  assign n7654 = ~n7655 | ~n14904;
  assign n7655 = ~n14901 | ~n14900;
  assign n7789 = ~n8095 | ~n8096;
  assign n7656 = ~n7782 | ~SI_1_;
  assign n8060 = ~n7783 | ~n7782;
  assign n14788 = ~n14785 | ~n14786;
  assign n8410 = ~n7300 | ~n7308;
  assign n11768 = ~n8085 | ~n12357;
  assign n14694 = n14966 & n14693;
  assign n14724 = n14723 & n14722;
  assign n14653 = ~n11843;
  assign n14703 = ~n14697 & ~n14696;
  assign n14696 = n14695 & n14694;
  assign n7855 = ~P1_IR_REG_16__SCAN_IN & ~P1_IR_REG_18__SCAN_IN;
  assign n7852 = n7851 & n7850;
  assign n7726 = ~P2_ADDR_REG_19__SCAN_IN;
  assign n7769 = n10536 | n11378;
  assign n8324 = n8307 & P1_REG3_REG_24__SCAN_IN;
  assign n8294 = n8282 & P1_REG3_REG_22__SCAN_IN;
  assign n8256 = n7944 & P1_REG3_REG_16__SCAN_IN;
  assign n7982 = n7996 & P1_REG3_REG_13__SCAN_IN;
  assign n8039 = n8223 & P1_REG3_REG_9__SCAN_IN;
  assign n8416 = n8434 & n8421;
  assign n7771 = ~n7769 | ~n7768;
  assign n9328 = n14621 | n15007;
  assign n8362 = ~n13698 | ~n14461;
  assign n8282 = n8270 & P1_REG3_REG_21__SCAN_IN;
  assign n7887 = n7905 & P1_REG3_REG_19__SCAN_IN;
  assign n8012 = n8030 & P1_REG3_REG_11__SCAN_IN;
  assign n11378 = ~P1_DATAO_REG_10__SCAN_IN;
  assign n11963 = ~n9579;
  assign n14616 = n9791 & n8435;
  assign n9996 = ~n9322;
  assign n7728 = ~n10535 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n7727 = ~n9339 | ~P2_DATAO_REG_25__SCAN_IN;
  assign n8319 = ~n7728 | ~n7727;
  assign n8321 = ~SI_25_ ^ n8319;
  assign n7730 = ~n10535 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n7729 = ~n10536 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n7731 = ~n7730 | ~n7729;
  assign n7847 = ~SI_24_ | ~n7731;
  assign n8303 = SI_24_ ^ n7731;
  assign n7733 = ~n10535 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n7732 = ~n9339 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n7734 = ~n7733 | ~n7732;
  assign n7845 = ~SI_23_ | ~n7734;
  assign n8292 = SI_23_ ^ n7734;
  assign n7736 = ~n10535 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n7735 = ~n10536 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n7737 = ~n7736 | ~n7735;
  assign n7843 = ~SI_22_ | ~n7737;
  assign n8279 = SI_22_ ^ n7737;
  assign n7739 = ~n10535 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n7738 = ~n10536 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n7740 = ~n7739 | ~n7738;
  assign n8267 = SI_21_ ^ n7740;
  assign n7742 = ~n10535 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n7741 = ~n9339 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n7743 = ~n7742 | ~n7741;
  assign n7841 = ~SI_20_ | ~n7743;
  assign n7884 = SI_20_ ^ n7743;
  assign n7745 = ~n10535 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n7744 = ~n9339 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n7746 = ~n7745 | ~n7744;
  assign n7840 = ~SI_19_ | ~n7746;
  assign n7896 = SI_19_ ^ n7746;
  assign n7748 = ~n9338 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n7747 = ~n10536 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n7749 = ~n7748 | ~n7747;
  assign n7838 = ~SI_18_ | ~n7749;
  assign n7914 = SI_18_ ^ n7749;
  assign n7751 = ~n9338 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n7750 = ~n10536 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n7752 = ~n7751 | ~n7750;
  assign n7837 = ~SI_17_ | ~n7752;
  assign n8246 = SI_17_ ^ n7752;
  assign n7754 = ~n9338 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n7753 = ~n10536 | ~P2_DATAO_REG_16__SCAN_IN;
  assign n7755 = ~n7754 | ~n7753;
  assign n7836 = ~SI_16_ | ~n7755;
  assign n7932 = SI_16_ ^ n7755;
  assign n7757 = ~n9338 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n7756 = ~n10536 | ~P2_DATAO_REG_15__SCAN_IN;
  assign n7833 = ~n7757 | ~n7756;
  assign n7835 = ~SI_15_ & ~n7833;
  assign n7759 = ~n9338 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n7758 = ~n9339 | ~P2_DATAO_REG_14__SCAN_IN;
  assign n7830 = ~n7759 | ~n7758;
  assign n7832 = ~SI_14_ & ~n7830;
  assign n7761 = ~n10535 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n7760 = ~n10536 | ~P2_DATAO_REG_13__SCAN_IN;
  assign n7762 = ~n7761 | ~n7760;
  assign n7829 = ~SI_13_ | ~n7762;
  assign n7987 = SI_13_ ^ n7762;
  assign n7764 = ~n10535 | ~P1_DATAO_REG_12__SCAN_IN;
  assign n7763 = ~n9339 | ~P2_DATAO_REG_12__SCAN_IN;
  assign n7826 = ~n7764 | ~n7763;
  assign n7828 = ~SI_12_ & ~n7826;
  assign n7766 = ~n10535 | ~P1_DATAO_REG_11__SCAN_IN;
  assign n7765 = ~n9339 | ~P2_DATAO_REG_11__SCAN_IN;
  assign n7767 = ~n7766 | ~n7765;
  assign n7825 = ~SI_11_ & ~n7767;
  assign n8020 = ~SI_11_ ^ n7767;
  assign n7768 = ~n9339 | ~P2_DATAO_REG_10__SCAN_IN;
  assign n7824 = ~SI_10_ | ~n7771;
  assign n7770 = ~SI_10_;
  assign n8046 = ~n7771 ^ n7770;
  assign n7772 = ~P1_DATAO_REG_0__SCAN_IN | ~P1_DATAO_REG_1__SCAN_IN;
  assign n7775 = n7796 | n7772;
  assign n7773 = P2_DATAO_REG_0__SCAN_IN & P2_DATAO_REG_1__SCAN_IN;
  assign n7774 = ~n7796 | ~n7773;
  assign n7776 = ~n7775 | ~n7774;
  assign n7783 = ~n7776 | ~SI_0_;
  assign n11084 = ~P1_DATAO_REG_1__SCAN_IN;
  assign n8688 = ~P1_DATAO_REG_0__SCAN_IN | ~SI_0_;
  assign n7777 = n11084 & n8688;
  assign n7781 = n7796 | n7777;
  assign n8068 = ~P2_DATAO_REG_1__SCAN_IN;
  assign n7778 = ~P2_DATAO_REG_0__SCAN_IN | ~SI_0_;
  assign n7779 = ~n8068 | ~n7778;
  assign n7780 = ~n7796 | ~n7779;
  assign n7782 = ~n7781 | ~n7780;
  assign n11127 = ~P1_DATAO_REG_2__SCAN_IN;
  assign n7785 = n7796 | n11127;
  assign n7784 = ~n7796 | ~P2_DATAO_REG_2__SCAN_IN;
  assign n7787 = ~n7785 | ~n7784;
  assign n7786 = ~SI_2_;
  assign n8095 = ~n7787 ^ n7786;
  assign n7788 = ~n7787 | ~SI_2_;
  assign n8116 = ~n7789 | ~n7788;
  assign n10996 = ~P1_DATAO_REG_3__SCAN_IN;
  assign n7791 = n7796 | n10996;
  assign n7790 = ~n7796 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n7793 = ~n7791 | ~n7790;
  assign n7792 = ~SI_3_;
  assign n8114 = ~n7793 ^ n7792;
  assign n7795 = ~n8116 | ~n8114;
  assign n7794 = ~n7793 | ~SI_3_;
  assign n8132 = ~n7795 | ~n7794;
  assign n11078 = ~P1_DATAO_REG_4__SCAN_IN;
  assign n7798 = n7796 | n11078;
  assign n7797 = ~n7796 | ~P2_DATAO_REG_4__SCAN_IN;
  assign n7800 = ~n7798 | ~n7797;
  assign n7799 = ~SI_4_;
  assign n8130 = ~n7800 ^ n7799;
  assign n7802 = ~n8132 | ~n8130;
  assign n7801 = ~n7800 | ~SI_4_;
  assign n8152 = ~n7802 | ~n7801;
  assign n7803 = ~n9339 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n7805 = ~n7804 | ~SI_5_;
  assign n9183 = ~P1_DATAO_REG_6__SCAN_IN;
  assign n7806 = ~n10536 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n7808 = ~n7807 | ~n7806;
  assign n7809 = ~n7808 | ~SI_6_;
  assign n11196 = ~P1_DATAO_REG_7__SCAN_IN;
  assign n7810 = ~n9339 | ~P2_DATAO_REG_7__SCAN_IN;
  assign n7812 = ~SI_7_;
  assign n8197 = ~n7813 ^ n7812;
  assign n7814 = ~n7813 | ~SI_7_;
  assign n7815 = ~n9339 | ~P2_DATAO_REG_8__SCAN_IN;
  assign n7818 = ~n7817 | ~SI_8_;
  assign n8213 = ~n7819 | ~n7818;
  assign n7820 = ~n10536 | ~P2_DATAO_REG_9__SCAN_IN;
  assign n8234 = ~n7822 ^ SI_9_;
  assign n7823 = ~n7822 | ~SI_9_;
  assign n8002 = ~SI_12_ ^ n7826;
  assign n7827 = ~n8003 & ~n8002;
  assign n7968 = ~SI_14_ ^ n7830;
  assign n7948 = ~SI_15_ ^ n7833;
  assign n7834 = ~n7949 & ~n7948;
  assign n7839 = ~n7896 | ~n7895;
  assign n7842 = ~n8279 | ~n8278;
  assign n7844 = ~n8292 | ~n8291;
  assign n7846 = ~n8303 | ~n8302;
  assign n13315 = n8321 ^ n8320;
  assign n9307 = ~n13315;
  assign n7858 = ~P1_IR_REG_21__SCAN_IN & ~P1_IR_REG_24__SCAN_IN;
  assign n7857 = ~P1_IR_REG_26__SCAN_IN;
  assign n7860 = n7858 & n7857;
  assign n7859 = ~P1_IR_REG_23__SCAN_IN & ~P1_IR_REG_25__SCAN_IN;
  assign n7861 = ~n7367 | ~P1_IR_REG_31__SCAN_IN;
  assign n9330 = n11097 | n14612;
  assign n8059 = ~n9330 | ~n9339;
  assign n7863 = ~n9307 | ~n14461;
  assign n8188 = ~n9330 | ~n9338;
  assign n8049 = ~n8188;
  assign n9308 = ~P2_DATAO_REG_25__SCAN_IN;
  assign n7862 = n8304 | n9308;
  assign n7864 = P1_REG3_REG_4__SCAN_IN & P1_REG3_REG_5__SCAN_IN;
  assign n8165 = ~n7864 | ~P1_REG3_REG_3__SCAN_IN;
  assign n8164 = ~P1_REG3_REG_6__SCAN_IN;
  assign n8181 = ~n8165 & ~n8164;
  assign n10172 = P1_REG3_REG_25__SCAN_IN ^ n8324;
  assign n7869 = ~n7868 | ~P1_IR_REG_31__SCAN_IN;
  assign n7872 = ~n7869 | ~P1_IR_REG_29__SCAN_IN;
  assign n7870 = ~P1_IR_REG_29__SCAN_IN;
  assign n7871 = ~n7870 | ~P1_IR_REG_31__SCAN_IN;
  assign n7873 = ~n7872 | ~n7871;
  assign n7874 = ~n9332;
  assign n8109 = n7877 & n7874;
  assign n7882 = ~n10172 | ~n8109;
  assign n8220 = ~n8105;
  assign n7876 = ~n8220 | ~P1_REG1_REG_25__SCAN_IN;
  assign n8069 = ~n7877 | ~n9332;
  assign n7875 = ~n7294 | ~P1_REG2_REG_25__SCAN_IN;
  assign n7880 = ~n7876 | ~n7875;
  assign n9345 = ~n7877;
  assign n8180 = n9345 & n9332;
  assign n7879 = n8180 & P1_REG0_REG_25__SCAN_IN;
  assign n7881 = ~n7880 & ~n7879;
  assign n11341 = ~n7882 | ~n7881;
  assign n10031 = ~n11341;
  assign n14805 = ~n10166 | ~n10031;
  assign n14761 = ~n14805;
  assign n14813 = ~n10170 | ~n11341;
  assign n14992 = ~n14813 | ~n14805;
  assign n12549 = ~n7884 ^ n7883;
  assign n7886 = ~n9265 | ~n14461;
  assign n9266 = ~P2_DATAO_REG_20__SCAN_IN;
  assign n7885 = n8304 | n9266;
  assign n14222 = ~P1_REG3_REG_20__SCAN_IN ^ n7887;
  assign n7888 = ~n14222;
  assign n7894 = ~n7888 | ~n8109;
  assign n7890 = ~n8380 | ~P1_REG1_REG_20__SCAN_IN;
  assign n7889 = ~n7294 | ~P1_REG2_REG_20__SCAN_IN;
  assign n7892 = ~n7890 | ~n7889;
  assign n7891 = n8180 & P1_REG0_REG_20__SCAN_IN;
  assign n7893 = ~n7892 & ~n7891;
  assign n13861 = ~n7894 | ~n7893;
  assign n14881 = ~n14230 & ~n13861;
  assign n12493 = ~n7896 ^ n7895;
  assign n8977 = ~n12493;
  assign n7904 = ~n8977 | ~n14461;
  assign n7897 = ~P2_DATAO_REG_19__SCAN_IN;
  assign n7902 = n8304 | n7897;
  assign n7899 = n7898 | P1_IR_REG_17__SCAN_IN;
  assign n7900 = ~n7899 | ~P1_IR_REG_31__SCAN_IN;
  assign n7901 = n9330 | n15005;
  assign n7903 = n7902 & n7901;
  assign n14126 = ~P1_REG3_REG_19__SCAN_IN ^ n7905;
  assign n7906 = ~n14126;
  assign n7912 = ~n7906 | ~n8109;
  assign n8380 = ~n8105;
  assign n7908 = ~n8380 | ~P1_REG1_REG_19__SCAN_IN;
  assign n7907 = ~n7294 | ~P1_REG2_REG_19__SCAN_IN;
  assign n7910 = ~n7908 | ~n7907;
  assign n7909 = n8180 & P1_REG0_REG_19__SCAN_IN;
  assign n7911 = ~n7910 & ~n7909;
  assign n13944 = ~n7912 | ~n7911;
  assign n14638 = ~n14132 & ~n13944;
  assign n12280 = ~n7914 ^ n7913;
  assign n8959 = ~n12280;
  assign n7922 = ~n8959 | ~n14461;
  assign n7915 = ~P2_DATAO_REG_18__SCAN_IN;
  assign n7920 = n8188 | n7915;
  assign n7916 = ~P1_IR_REG_16__SCAN_IN;
  assign n7917 = ~n7396 | ~n7916;
  assign n8249 = ~n7917 | ~P1_IR_REG_31__SCAN_IN;
  assign n8251 = ~n8249 | ~n8248;
  assign n7918 = ~n8251 | ~P1_IR_REG_31__SCAN_IN;
  assign n14098 = ~n7918 ^ P1_IR_REG_18__SCAN_IN;
  assign n14092 = ~n14098;
  assign n7919 = n9330 | n14092;
  assign n7921 = n7920 & n7919;
  assign n14068 = P1_REG3_REG_18__SCAN_IN ^ n7923;
  assign n7930 = ~n14068 | ~n8109;
  assign n7925 = ~n7294 | ~P1_REG2_REG_18__SCAN_IN;
  assign n7924 = ~n8180 | ~P1_REG0_REG_18__SCAN_IN;
  assign n7928 = ~n7925 | ~n7924;
  assign n7926 = ~P1_REG1_REG_18__SCAN_IN;
  assign n7927 = ~n8105 & ~n7926;
  assign n7929 = ~n7928 & ~n7927;
  assign n13862 = ~n7930 | ~n7929;
  assign n14729 = n13776 | n13862;
  assign n14982 = ~n7311 | ~n14729;
  assign n11893 = ~n7932 ^ n7931;
  assign n8922 = ~n11893;
  assign n7938 = ~n8922 | ~n14461;
  assign n7933 = ~P2_DATAO_REG_16__SCAN_IN;
  assign n7936 = n8304 | n7933;
  assign n8229 = ~P1_IR_REG_31__SCAN_IN;
  assign n7934 = n7396 | n8229;
  assign n13639 = ~n7934 ^ P1_IR_REG_16__SCAN_IN;
  assign n13630 = ~n13639;
  assign n7935 = n9330 | n13630;
  assign n7937 = n7936 & n7935;
  assign n7940 = ~n8180 | ~P1_REG0_REG_16__SCAN_IN;
  assign n7939 = ~n7294 | ~P1_REG2_REG_16__SCAN_IN;
  assign n7943 = ~n7940 | ~n7939;
  assign n7941 = ~P1_REG1_REG_16__SCAN_IN;
  assign n7942 = ~n8105 & ~n7941;
  assign n7946 = ~n7943 & ~n7942;
  assign n13816 = P1_REG3_REG_16__SCAN_IN ^ n7944;
  assign n7945 = ~n13816 | ~n8109;
  assign n13591 = ~n7946 | ~n7945;
  assign n7947 = ~n13591;
  assign n14714 = n13821 | n7947;
  assign n14821 = ~n13821 | ~n7947;
  assign n11782 = n7949 ^ n7948;
  assign n8905 = ~n11782;
  assign n7956 = ~n8905 | ~n14461;
  assign n7950 = ~P2_DATAO_REG_15__SCAN_IN;
  assign n7954 = n8304 | n7950;
  assign n7952 = ~n7951 | ~P1_IR_REG_31__SCAN_IN;
  assign n13152 = ~n7952 ^ P1_IR_REG_15__SCAN_IN;
  assign n13143 = ~n13152;
  assign n7953 = n9330 | n13143;
  assign n7955 = n7954 & n7953;
  assign n7958 = ~n7294 | ~P1_REG2_REG_15__SCAN_IN;
  assign n7957 = ~n8180 | ~P1_REG0_REG_15__SCAN_IN;
  assign n7961 = ~n7958 | ~n7957;
  assign n7959 = ~P1_REG1_REG_15__SCAN_IN;
  assign n7960 = ~n8105 & ~n7959;
  assign n7964 = ~n7961 & ~n7960;
  assign n13486 = P1_REG3_REG_15__SCAN_IN ^ n7962;
  assign n7963 = ~n13486 | ~n8109;
  assign n13661 = ~n7964 | ~n7963;
  assign n7965 = ~n13661;
  assign n14823 = ~n13608 & ~n7965;
  assign n14855 = ~n13608 | ~n7965;
  assign n7966 = ~n14855;
  assign n7977 = ~n8890 | ~n14461;
  assign n7969 = ~P2_DATAO_REG_14__SCAN_IN;
  assign n7975 = n8304 | n7969;
  assign n7970 = n8004 | P1_IR_REG_12__SCAN_IN;
  assign n7989 = ~n7970 | ~P1_IR_REG_31__SCAN_IN;
  assign n7971 = ~P1_IR_REG_13__SCAN_IN;
  assign n7972 = ~n7989 | ~n7971;
  assign n7973 = ~n7972 | ~P1_IR_REG_31__SCAN_IN;
  assign n12852 = ~n7973 ^ P1_IR_REG_14__SCAN_IN;
  assign n12399 = ~n12852;
  assign n7974 = n9330 | n12399;
  assign n7976 = n7975 & n7974;
  assign n7979 = ~n8380 | ~P1_REG1_REG_14__SCAN_IN;
  assign n7978 = ~n8180 | ~P1_REG0_REG_14__SCAN_IN;
  assign n7981 = ~n7979 | ~n7978;
  assign n7980 = n7294 & P1_REG2_REG_14__SCAN_IN;
  assign n7984 = ~n7981 & ~n7980;
  assign n13551 = P1_REG3_REG_14__SCAN_IN ^ n7982;
  assign n7983 = ~n8109 | ~n13551;
  assign n13221 = ~n7984 | ~n7983;
  assign n7985 = ~n13221;
  assign n14706 = ~n13683 | ~n7985;
  assign n14858 = ~n14706;
  assign n14853 = ~n13683 & ~n7985;
  assign n11592 = ~n7987 ^ n7986;
  assign n8851 = ~n11592;
  assign n7993 = ~n8851 | ~n14461;
  assign n7988 = ~P2_DATAO_REG_13__SCAN_IN;
  assign n7991 = n8304 | n7988;
  assign n12400 = ~n7989 ^ P1_IR_REG_13__SCAN_IN;
  assign n12393 = ~n12400;
  assign n7990 = n9330 | n12393;
  assign n7992 = n7991 & n7990;
  assign n7995 = ~n8380 | ~P1_REG1_REG_13__SCAN_IN;
  assign n7994 = ~n7294 | ~P1_REG2_REG_13__SCAN_IN;
  assign n8001 = ~n7995 | ~n7994;
  assign n7999 = ~n8180 | ~P1_REG0_REG_13__SCAN_IN;
  assign n13321 = ~P1_REG3_REG_13__SCAN_IN ^ n7996;
  assign n7997 = ~n13321;
  assign n7998 = ~n8109 | ~n7997;
  assign n8000 = ~n7999 | ~n7998;
  assign n8037 = ~n14701;
  assign n8038 = ~n13387 | ~n13523;
  assign n11538 = ~n8003 ^ n8002;
  assign n8009 = ~n11538 | ~n14461;
  assign n11530 = ~P2_DATAO_REG_12__SCAN_IN;
  assign n8007 = n8304 | n11530;
  assign n8005 = ~n8004 | ~P1_IR_REG_31__SCAN_IN;
  assign n11949 = ~n8005 ^ P1_IR_REG_12__SCAN_IN;
  assign n11939 = ~n11949;
  assign n8006 = n9330 | n11939;
  assign n8008 = n8007 & n8006;
  assign n8011 = ~n8220 | ~P1_REG1_REG_12__SCAN_IN;
  assign n8010 = ~n7294 | ~P1_REG2_REG_12__SCAN_IN;
  assign n8017 = ~n8011 | ~n8010;
  assign n8015 = ~n8180 | ~P1_REG0_REG_12__SCAN_IN;
  assign n13194 = ~P1_REG3_REG_12__SCAN_IN ^ n8012;
  assign n8013 = ~n13194;
  assign n8014 = ~n8109 | ~n8013;
  assign n8016 = ~n8015 | ~n8014;
  assign n8018 = ~n13200 | ~n13223;
  assign n14702 = ~n8038 | ~n8018;
  assign n14698 = ~n13200 & ~n13223;
  assign n11374 = ~n8020 ^ n8019;
  assign n8027 = ~n11374 | ~n14461;
  assign n11366 = ~P2_DATAO_REG_11__SCAN_IN;
  assign n8025 = n8188 | n11366;
  assign n8021 = ~P1_IR_REG_9__SCAN_IN;
  assign n8022 = ~n8230 | ~n8021;
  assign n8052 = ~n8022 | ~P1_IR_REG_31__SCAN_IN;
  assign n8051 = ~P1_IR_REG_10__SCAN_IN;
  assign n8054 = ~n8052 | ~n8051;
  assign n8023 = ~n8054 | ~P1_IR_REG_31__SCAN_IN;
  assign n11615 = ~n8023 ^ P1_IR_REG_11__SCAN_IN;
  assign n11622 = ~n11615;
  assign n8024 = n9330 | n11622;
  assign n8026 = n8025 & n8024;
  assign n8029 = ~n8220 | ~P1_REG1_REG_11__SCAN_IN;
  assign n8028 = ~n7294 | ~P1_REG2_REG_11__SCAN_IN;
  assign n8035 = ~n8029 | ~n8028;
  assign n8033 = ~n8180 | ~P1_REG0_REG_11__SCAN_IN;
  assign n13206 = ~P1_REG3_REG_11__SCAN_IN ^ n8030;
  assign n8031 = ~n13206;
  assign n8032 = ~n8109 | ~n8031;
  assign n8034 = ~n8033 | ~n8032;
  assign n8490 = ~n13212 | ~n12982;
  assign n8036 = ~n14698 & ~n8490;
  assign n14645 = ~n14702 & ~n8036;
  assign n14852 = ~n8037 & ~n14645;
  assign n13331 = ~n14701 | ~n8038;
  assign n8041 = ~n8380 | ~P1_REG1_REG_10__SCAN_IN;
  assign n12872 = P1_REG3_REG_10__SCAN_IN ^ n8039;
  assign n8040 = ~n8109 | ~n12872;
  assign n8045 = ~n8041 | ~n8040;
  assign n8043 = ~n8180 | ~P1_REG0_REG_10__SCAN_IN;
  assign n8042 = ~n7294 | ~P1_REG2_REG_10__SCAN_IN;
  assign n8044 = ~n8043 | ~n8042;
  assign n8047 = ~n8046;
  assign n11377 = ~n8048 ^ n8047;
  assign n8058 = ~n11377 | ~n14461;
  assign n8050 = ~P2_DATAO_REG_10__SCAN_IN;
  assign n8056 = n8304 | n8050;
  assign n8053 = n8052 | n8051;
  assign n11515 = n8054 & n8053;
  assign n11384 = ~n11515;
  assign n8055 = n9330 | n11384;
  assign n8057 = n8056 & n8055;
  assign n14868 = ~n10992 & ~n12873;
  assign n8061 = ~n8059;
  assign n11001 = ~n8060 ^ SI_1_;
  assign n8067 = ~n8118;
  assign n8062 = ~P1_IR_REG_1__SCAN_IN;
  assign n8065 = ~n8062 | ~P1_IR_REG_31__SCAN_IN;
  assign n8063 = ~P1_IR_REG_31__SCAN_IN | ~P1_IR_REG_0__SCAN_IN;
  assign n8064 = ~n8063 | ~P1_IR_REG_1__SCAN_IN;
  assign n8066 = ~n8065 | ~n8064;
  assign n11152 = n8067 & n8066;
  assign n11022 = ~n11152;
  assign n8071 = ~n7294 | ~P1_REG2_REG_1__SCAN_IN;
  assign n8070 = ~n8380 | ~P1_REG1_REG_1__SCAN_IN;
  assign n8075 = ~n8071 | ~n8070;
  assign n8073 = ~n8180 | ~P1_REG0_REG_1__SCAN_IN;
  assign n8072 = ~n8109 | ~P1_REG3_REG_1__SCAN_IN;
  assign n8074 = ~n8073 | ~n8072;
  assign n8088 = ~n14913;
  assign n8086 = ~n11766 | ~n11997;
  assign n8077 = ~n8380 | ~P1_REG1_REG_0__SCAN_IN;
  assign n8076 = ~n8180 | ~P1_REG0_REG_0__SCAN_IN;
  assign n8081 = ~n8077 | ~n8076;
  assign n8079 = ~n7294 | ~P1_REG2_REG_0__SCAN_IN;
  assign n8078 = ~n8109 | ~P1_REG3_REG_0__SCAN_IN;
  assign n8085 = ~n11767;
  assign n9562 = ~P1_IR_REG_0__SCAN_IN;
  assign n8084 = n9330 | n9562;
  assign n8082 = ~n9339 | ~SI_0_;
  assign n10942 = ~n8082 ^ P2_DATAO_REG_0__SCAN_IN;
  assign n8083 = ~n9330 | ~n10942;
  assign n12357 = ~n8084 | ~n8083;
  assign n8087 = ~n8086 | ~n11768;
  assign n8103 = ~n12008;
  assign n8090 = ~n8220 | ~P1_REG1_REG_2__SCAN_IN;
  assign n8089 = ~n7294 | ~P1_REG2_REG_2__SCAN_IN;
  assign n8094 = ~n8090 | ~n8089;
  assign n8092 = ~n8180 | ~P1_REG0_REG_2__SCAN_IN;
  assign n8091 = ~n8109 | ~P1_REG3_REG_2__SCAN_IN;
  assign n8093 = ~n8092 | ~n8091;
  assign n8097 = ~n8095;
  assign n11125 = ~n8097 ^ n8096;
  assign n8100 = ~n8061 | ~n11125;
  assign n8098 = n8229 | n8118;
  assign n11025 = ~n8098 ^ P1_IR_REG_2__SCAN_IN;
  assign n11393 = ~n11025;
  assign n8099 = n9330 | n11393;
  assign n8102 = ~n8100 | ~n8099;
  assign n9161 = ~P2_DATAO_REG_2__SCAN_IN;
  assign n8101 = ~n8188 & ~n9161;
  assign n12017 = ~n12384;
  assign n8104 = ~n8103 | ~n14914;
  assign n8472 = ~n9579 | ~n12384;
  assign n14831 = ~n8104 | ~n8472;
  assign n8107 = ~n8220 | ~P1_REG1_REG_3__SCAN_IN;
  assign n8106 = ~n7294 | ~P1_REG2_REG_3__SCAN_IN;
  assign n8113 = ~n8107 | ~n8106;
  assign n8111 = ~n8180 | ~P1_REG0_REG_3__SCAN_IN;
  assign n8108 = ~P1_REG3_REG_3__SCAN_IN;
  assign n8110 = ~n8109 | ~n8108;
  assign n8112 = ~n8111 | ~n8110;
  assign n8115 = ~n8114;
  assign n10984 = ~n8116 ^ n8115;
  assign n8121 = ~n8061 | ~n10984;
  assign n8117 = ~P1_IR_REG_2__SCAN_IN;
  assign n8119 = ~n8118 | ~n8117;
  assign n8134 = ~n8119 | ~P1_IR_REG_31__SCAN_IN;
  assign n8133 = ~P1_IR_REG_3__SCAN_IN;
  assign n11052 = ~n8134 ^ P1_IR_REG_3__SCAN_IN;
  assign n10985 = ~n11052;
  assign n8120 = n9330 | n10985;
  assign n8124 = ~n8121 | ~n8120;
  assign n8122 = ~P2_DATAO_REG_3__SCAN_IN;
  assign n8123 = ~n8188 & ~n8122;
  assign n14871 = ~n9590 | ~n12156;
  assign n11920 = ~n9590;
  assign n12178 = ~n12156;
  assign n14917 = ~n11920 | ~n12178;
  assign n14944 = ~n14871 | ~n14917;
  assign n11971 = ~n14944;
  assign n8125 = ~n14831 | ~n11971;
  assign n8127 = ~n8380 | ~P1_REG1_REG_4__SCAN_IN;
  assign n8126 = ~n7294 | ~P1_REG2_REG_4__SCAN_IN;
  assign n12227 = ~P1_REG3_REG_3__SCAN_IN ^ P1_REG3_REG_4__SCAN_IN;
  assign n8128 = ~n12227;
  assign n8129 = ~n8109 | ~n8128;
  assign n8131 = ~n8130;
  assign n11076 = ~n8132 ^ n8131;
  assign n8138 = ~n8061 | ~n11076;
  assign n8135 = ~n8134 | ~n8133;
  assign n8136 = ~n8135 | ~P1_IR_REG_31__SCAN_IN;
  assign n11051 = ~n8136 ^ P1_IR_REG_4__SCAN_IN;
  assign n11441 = ~n11051;
  assign n8137 = n9330 | n11441;
  assign n8140 = ~n8138 | ~n8137;
  assign n9156 = ~P2_DATAO_REG_4__SCAN_IN;
  assign n8139 = ~n8188 & ~n9156;
  assign n12236 = n8140 | n8139;
  assign n14832 = ~n9601 | ~n12236;
  assign n8142 = ~n8220 | ~P1_REG1_REG_5__SCAN_IN;
  assign n8141 = ~n7294 | ~P1_REG2_REG_5__SCAN_IN;
  assign n8150 = ~n8142 | ~n8141;
  assign n8148 = ~n8180 | ~P1_REG0_REG_5__SCAN_IN;
  assign n8144 = ~P1_REG3_REG_5__SCAN_IN;
  assign n8143 = ~P1_REG3_REG_3__SCAN_IN | ~P1_REG3_REG_4__SCAN_IN;
  assign n8145 = ~n8144 | ~n8143;
  assign n12261 = ~n8165 | ~n8145;
  assign n8146 = ~n12261;
  assign n8147 = ~n8109 | ~n8146;
  assign n8149 = ~n8148 | ~n8147;
  assign n9171 = ~n8152 ^ n8151;
  assign n8159 = ~n8061 | ~n9171;
  assign n8154 = ~n8153 | ~P1_IR_REG_31__SCAN_IN;
  assign n8156 = ~n8154 | ~P1_IR_REG_5__SCAN_IN;
  assign n8155 = ~n7848 | ~P1_IR_REG_31__SCAN_IN;
  assign n8157 = ~n8156 | ~n8155;
  assign n11140 = n8189 & n8157;
  assign n11060 = ~n11140;
  assign n8158 = n9330 | n11060;
  assign n8161 = ~n8159 | ~n8158;
  assign n9172 = ~P2_DATAO_REG_5__SCAN_IN;
  assign n8160 = ~n8188 & ~n9172;
  assign n14833 = ~n10772 | ~n11906;
  assign n11919 = ~n10772;
  assign n12269 = ~n11906;
  assign n14672 = ~n11919 | ~n12269;
  assign n14947 = ~n14833 | ~n14672;
  assign n8163 = ~n8220 | ~P1_REG1_REG_6__SCAN_IN;
  assign n8162 = ~n7294 | ~P1_REG2_REG_6__SCAN_IN;
  assign n8169 = ~n8163 | ~n8162;
  assign n8166 = n8165 & n8164;
  assign n12216 = n8166 | n8181;
  assign n8167 = ~n12216;
  assign n8168 = ~n8109 | ~n8167;
  assign n9182 = ~n8171 ^ n8170;
  assign n8174 = ~n8061 | ~n9182;
  assign n8172 = ~n8189 | ~P1_IR_REG_31__SCAN_IN;
  assign n11112 = ~n8172 ^ P1_IR_REG_6__SCAN_IN;
  assign n11105 = ~n11112;
  assign n8173 = n9330 | n11105;
  assign n8176 = ~n8174 | ~n8173;
  assign n9177 = ~P2_DATAO_REG_6__SCAN_IN;
  assign n8175 = ~n8304 & ~n9177;
  assign n14671 = ~n9549 | ~n12184;
  assign n12197 = ~n9549;
  assign n12221 = ~n12184;
  assign n14673 = ~n12197 | ~n12221;
  assign n14953 = ~n14671 | ~n14673;
  assign n14835 = ~n14671;
  assign n8179 = ~n8380 | ~P1_REG1_REG_7__SCAN_IN;
  assign n8178 = ~n7294 | ~P1_REG2_REG_7__SCAN_IN;
  assign n8186 = ~n8179 | ~n8178;
  assign n8184 = ~n8180 | ~P1_REG0_REG_7__SCAN_IN;
  assign n12815 = ~n8181 ^ P1_REG3_REG_7__SCAN_IN;
  assign n8182 = ~n12815;
  assign n8183 = ~n8109 | ~n8182;
  assign n8185 = ~n8184 | ~n8183;
  assign n8187 = ~P2_DATAO_REG_7__SCAN_IN;
  assign n8196 = n8188 | n8187;
  assign n8190 = ~n8189 & ~P1_IR_REG_6__SCAN_IN;
  assign n8191 = ~n8190 & ~n8229;
  assign n8194 = ~n8191 | ~P1_IR_REG_7__SCAN_IN;
  assign n8193 = ~n8191;
  assign n8192 = ~P1_IR_REG_7__SCAN_IN;
  assign n8209 = ~n8193 | ~n8192;
  assign n11260 = n8194 & n8209;
  assign n11252 = ~n11260;
  assign n8195 = n9330 | n11252;
  assign n8200 = n8196 & n8195;
  assign n8198 = ~n8197;
  assign n8199 = ~n8061 | ~n11182;
  assign n14650 = ~n12365 | ~n12820;
  assign n9197 = ~n12365;
  assign n12771 = ~n12820;
  assign n14676 = ~n9197 | ~n12771;
  assign n8202 = ~n8220 | ~P1_REG1_REG_8__SCAN_IN;
  assign n8201 = ~n7294 | ~P1_REG2_REG_8__SCAN_IN;
  assign n8208 = ~n8202 | ~n8201;
  assign n8206 = ~n8180 | ~P1_REG0_REG_8__SCAN_IN;
  assign n12521 = ~P1_REG3_REG_8__SCAN_IN ^ n8203;
  assign n8204 = ~n12521;
  assign n8205 = ~n8109 | ~n8204;
  assign n8207 = ~n8206 | ~n8205;
  assign n8482 = ~n12626;
  assign n11293 = ~P2_DATAO_REG_8__SCAN_IN;
  assign n8212 = n8304 | n11293;
  assign n8210 = ~n8209 | ~P1_IR_REG_31__SCAN_IN;
  assign n11275 = ~n8210 ^ P1_IR_REG_8__SCAN_IN;
  assign n11294 = ~n11275;
  assign n8211 = n9330 | n11294;
  assign n8218 = n8212 & n8211;
  assign n8215 = ~n8214 | ~n8213;
  assign n11302 = ~n8216 | ~n8215;
  assign n8217 = ~n8061 | ~n11302;
  assign n12556 = ~n8218 | ~n8217;
  assign n14666 = ~n8482 | ~n12556;
  assign n12377 = ~n12556;
  assign n14840 = ~n12626 | ~n12377;
  assign n8222 = ~n8220 | ~P1_REG1_REG_9__SCAN_IN;
  assign n8221 = ~n7294 | ~P1_REG2_REG_9__SCAN_IN;
  assign n8227 = ~n8222 | ~n8221;
  assign n8225 = ~n8180 | ~P1_REG0_REG_9__SCAN_IN;
  assign n12679 = P1_REG3_REG_9__SCAN_IN ^ n8223;
  assign n8224 = ~n8109 | ~n12679;
  assign n8226 = ~n8225 | ~n8224;
  assign n8228 = ~P2_DATAO_REG_9__SCAN_IN;
  assign n8233 = n8304 | n8228;
  assign n8231 = n8230 | n8229;
  assign n11311 = ~n8231 ^ P1_IR_REG_9__SCAN_IN;
  assign n11336 = ~n11311;
  assign n8232 = n9330 | n11336;
  assign n8238 = n8233 & n8232;
  assign n8235 = ~n8234;
  assign n11329 = ~n8236 ^ n8235;
  assign n8237 = ~n8061 | ~n11329;
  assign n14825 = ~n12364 & ~n12680;
  assign n14683 = ~n12364 | ~n12680;
  assign n14692 = ~n10992 | ~n12873;
  assign n14846 = ~n14683 | ~n14692;
  assign n8491 = ~n12982;
  assign n14646 = ~n13175 | ~n8491;
  assign n12977 = ~n13200;
  assign n8242 = ~n12977 | ~n13223;
  assign n8241 = ~n13223;
  assign n8493 = ~n13200 | ~n8241;
  assign n14967 = ~n8242 | ~n8493;
  assign n14851 = ~n14698;
  assign n12128 = ~n8246 ^ n8245;
  assign n8941 = ~n12128;
  assign n8255 = ~n8941 | ~n14461;
  assign n8247 = ~P2_DATAO_REG_17__SCAN_IN;
  assign n8253 = n8188 | n8247;
  assign n8250 = n8249 | n8248;
  assign n13888 = n8251 & n8250;
  assign n13638 = ~n13888;
  assign n8252 = n9330 | n13638;
  assign n8254 = n8253 & n8252;
  assign n13832 = P1_REG3_REG_17__SCAN_IN ^ n8256;
  assign n8263 = ~n13832 | ~n8109;
  assign n8258 = ~n8180 | ~P1_REG0_REG_17__SCAN_IN;
  assign n8257 = ~n7294 | ~P1_REG2_REG_17__SCAN_IN;
  assign n8261 = ~n8258 | ~n8257;
  assign n8259 = ~P1_REG1_REG_17__SCAN_IN;
  assign n8260 = ~n8105 & ~n8259;
  assign n8262 = ~n8261 & ~n8260;
  assign n13757 = ~n8263 | ~n8262;
  assign n8264 = ~n13757;
  assign n14715 = n13833 | n8264;
  assign n14822 = ~n13833 | ~n8264;
  assign n14639 = ~n14132 | ~n13944;
  assign n14637 = ~n14230 | ~n13861;
  assign n14878 = ~n14639 | ~n14637;
  assign n12736 = ~n8267 ^ n8266;
  assign n8269 = ~n12733 | ~n14461;
  assign n12730 = ~P2_DATAO_REG_21__SCAN_IN;
  assign n8268 = n8188 | n12730;
  assign n14003 = ~P1_REG3_REG_21__SCAN_IN ^ n8270;
  assign n9794 = ~n14003;
  assign n8276 = ~n9794 | ~n8109;
  assign n8272 = ~n8380 | ~P1_REG1_REG_21__SCAN_IN;
  assign n8271 = ~n7294 | ~P1_REG2_REG_21__SCAN_IN;
  assign n8274 = ~n8272 | ~n8271;
  assign n8273 = n8180 & P1_REG0_REG_21__SCAN_IN;
  assign n8275 = ~n8274 & ~n8273;
  assign n13942 = ~n8276 | ~n8275;
  assign n14633 = ~n14025 | ~n13942;
  assign n12899 = ~n8279 ^ n8278;
  assign n8281 = ~n12896 | ~n14461;
  assign n12893 = ~P2_DATAO_REG_22__SCAN_IN;
  assign n8280 = n8304 | n12893;
  assign n14188 = ~P1_REG3_REG_22__SCAN_IN ^ n8282;
  assign n9862 = ~n14188;
  assign n8288 = ~n9862 | ~n8109;
  assign n8284 = ~n8380 | ~P1_REG1_REG_22__SCAN_IN;
  assign n8283 = ~n7294 | ~P1_REG2_REG_22__SCAN_IN;
  assign n8286 = ~n8284 | ~n8283;
  assign n8285 = n8180 & P1_REG0_REG_22__SCAN_IN;
  assign n8287 = ~n8286 & ~n8285;
  assign n11166 = ~n8288 | ~n8287;
  assign n8289 = ~n11166;
  assign n14816 = n14193 & n8289;
  assign n14632 = ~n14816;
  assign n14988 = ~n14632 | ~n14634;
  assign n13083 = ~P2_DATAO_REG_23__SCAN_IN;
  assign n8293 = n8304 | n13083;
  assign n14259 = ~P1_REG3_REG_23__SCAN_IN ^ n8294;
  assign n10087 = ~n14259;
  assign n8300 = ~n10087 | ~n8109;
  assign n8296 = ~n8380 | ~P1_REG1_REG_23__SCAN_IN;
  assign n8295 = ~n7294 | ~P1_REG2_REG_23__SCAN_IN;
  assign n8298 = ~n8296 | ~n8295;
  assign n8297 = n8180 & P1_REG0_REG_23__SCAN_IN;
  assign n8299 = ~n8298 & ~n8297;
  assign n11272 = ~n8300 | ~n8299;
  assign n14740 = ~n14336 | ~n11272;
  assign n14748 = ~n14740;
  assign n13186 = ~n8303 ^ n8302;
  assign n8306 = ~n13139 | ~n14461;
  assign n13136 = ~P2_DATAO_REG_24__SCAN_IN;
  assign n8305 = n8304 | n13136;
  assign n14414 = ~P1_REG3_REG_24__SCAN_IN ^ n8307;
  assign n10148 = ~n14414;
  assign n8313 = ~n10148 | ~n8109;
  assign n8309 = ~n8380 | ~P1_REG1_REG_24__SCAN_IN;
  assign n8308 = ~n7294 | ~P1_REG2_REG_24__SCAN_IN;
  assign n8311 = ~n8309 | ~n8308;
  assign n8310 = n8180 & P1_REG0_REG_24__SCAN_IN;
  assign n8312 = ~n8311 & ~n8310;
  assign n11323 = ~n8313 | ~n8312;
  assign n8314 = ~n11323;
  assign n8315 = ~n14888;
  assign n14424 = ~n8315 | ~n14758;
  assign n14990 = ~n14424;
  assign n8318 = ~n10535 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n8317 = ~n10536 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n8334 = ~n8318 | ~n8317;
  assign n8336 = SI_26_ ^ n8334;
  assign n13456 = ~n8336 ^ n8335;
  assign n8323 = ~n13408 | ~n14461;
  assign n13403 = ~P2_DATAO_REG_26__SCAN_IN;
  assign n8322 = n8188 | n13403;
  assign n8342 = ~n8324 | ~P1_REG3_REG_25__SCAN_IN;
  assign n10227 = ~n8342 ^ P1_REG3_REG_26__SCAN_IN;
  assign n8330 = ~n10227 | ~n8109;
  assign n8326 = ~n8380 | ~P1_REG1_REG_26__SCAN_IN;
  assign n8325 = ~n7294 | ~P1_REG2_REG_26__SCAN_IN;
  assign n8328 = ~n8326 | ~n8325;
  assign n8327 = n8180 & P1_REG0_REG_26__SCAN_IN;
  assign n8329 = ~n8328 & ~n8327;
  assign n11326 = ~n8330 | ~n8329;
  assign n8331 = ~n11326;
  assign n14806 = ~n10225 | ~n8331;
  assign n8333 = ~n10535 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n8332 = ~n10536 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n8354 = ~n8333 | ~n8332;
  assign n8356 = SI_27_ ^ n8354;
  assign n8338 = ~SI_26_ | ~n8334;
  assign n8340 = ~n7309 | ~n14461;
  assign n9313 = ~P2_DATAO_REG_27__SCAN_IN;
  assign n8339 = n8304 | n9313;
  assign n8341 = ~P1_REG3_REG_26__SCAN_IN;
  assign n8363 = ~n8342 & ~n8341;
  assign n10295 = P1_REG3_REG_27__SCAN_IN ^ n8363;
  assign n8348 = ~n10295 | ~n8109;
  assign n8344 = ~n8380 | ~P1_REG1_REG_27__SCAN_IN;
  assign n8343 = ~n7294 | ~P1_REG2_REG_27__SCAN_IN;
  assign n8346 = ~n8344 | ~n8343;
  assign n8345 = n8180 & P1_REG0_REG_27__SCAN_IN;
  assign n8347 = ~n8346 & ~n8345;
  assign n11527 = ~n8348 | ~n8347;
  assign n10032 = ~n11527;
  assign n8351 = ~n14770;
  assign n8358 = ~SI_27_ | ~n8354;
  assign n8357 = ~n8356 | ~n8355;
  assign n8360 = ~n10535 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n8359 = ~n9339 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n8373 = ~n8360 | ~n8359;
  assign n8374 = ~SI_28_ ^ n8373;
  assign n9317 = ~P2_DATAO_REG_28__SCAN_IN;
  assign n8361 = n8188 | n9317;
  assign n8379 = n8363 & P1_REG3_REG_27__SCAN_IN;
  assign n10708 = P1_REG3_REG_28__SCAN_IN ^ n8379;
  assign n8369 = ~n10708 | ~n8109;
  assign n8365 = ~n8380 | ~P1_REG1_REG_28__SCAN_IN;
  assign n8364 = ~n8180 | ~P1_REG0_REG_28__SCAN_IN;
  assign n8367 = ~n8365 | ~n8364;
  assign n8366 = n7294 & P1_REG2_REG_28__SCAN_IN;
  assign n8368 = ~n8367 & ~n8366;
  assign n11635 = ~n8369 | ~n8368;
  assign n10698 = ~n11635;
  assign n14622 = ~n10691 | ~n10698;
  assign n14802 = ~n10706 | ~n11635;
  assign n8372 = ~n10535 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n8371 = ~n9339 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n9344 = ~n8372 | ~n8371;
  assign n9342 = SI_29_ ^ n9344;
  assign n8376 = ~SI_28_ & ~n8373;
  assign n9322 = ~n9342 ^ n9343;
  assign n8378 = ~n9996 | ~n14461;
  assign n9333 = ~P2_DATAO_REG_29__SCAN_IN;
  assign n8377 = n8188 | n9333;
  assign n8540 = n8379 & P1_REG3_REG_28__SCAN_IN;
  assign n8386 = ~n8540 | ~n8109;
  assign n8382 = ~n8380 | ~P1_REG1_REG_29__SCAN_IN;
  assign n8381 = ~n7294 | ~P1_REG2_REG_29__SCAN_IN;
  assign n8384 = ~n8382 | ~n8381;
  assign n8383 = n8180 & P1_REG0_REG_29__SCAN_IN;
  assign n8385 = ~n8384 & ~n8383;
  assign n11570 = ~n8386 | ~n8385;
  assign n8387 = ~n11570;
  assign n8392 = ~n7293 | ~P1_IR_REG_31__SCAN_IN;
  assign n8533 = ~n8392 ^ P1_IR_REG_21__SCAN_IN;
  assign n8390 = ~n8389 | ~P1_IR_REG_31__SCAN_IN;
  assign n15009 = ~n8390 ^ P1_IR_REG_20__SCAN_IN;
  assign n14903 = n8533 & n15009;
  assign n8391 = ~P1_IR_REG_21__SCAN_IN;
  assign n8393 = ~n8392 | ~n8391;
  assign n8395 = ~n8393 | ~P1_IR_REG_31__SCAN_IN;
  assign n9779 = ~n9328;
  assign n13222 = n11097 & n9779;
  assign n14614 = ~n13222;
  assign n8400 = ~n7294 | ~P1_REG2_REG_30__SCAN_IN;
  assign n8399 = ~n8180 | ~P1_REG0_REG_30__SCAN_IN;
  assign n8403 = ~n8400 | ~n8399;
  assign n8401 = ~P1_REG1_REG_30__SCAN_IN;
  assign n8402 = ~n8105 & ~n8401;
  assign n14798 = n8403 | n8402;
  assign n8434 = ~n8411 | ~P1_IR_REG_31__SCAN_IN;
  assign n8421 = ~P1_IR_REG_31__SCAN_IN | ~P1_IR_REG_23__SCAN_IN;
  assign n8412 = ~P1_IR_REG_24__SCAN_IN;
  assign n8413 = n8421 & n8412;
  assign n8414 = ~n8434 | ~n8413;
  assign n8415 = ~n8414 | ~P1_IR_REG_31__SCAN_IN;
  assign n8431 = ~n8415 ^ P1_IR_REG_25__SCAN_IN;
  assign n8430 = ~n8416 ^ P1_IR_REG_24__SCAN_IN;
  assign n8420 = ~P1_IR_REG_24__SCAN_IN & ~P1_IR_REG_25__SCAN_IN;
  assign n8422 = n8421 & n8420;
  assign n8423 = ~n8434 | ~n8422;
  assign n8424 = ~n8423 | ~P1_IR_REG_31__SCAN_IN;
  assign n9791 = ~n13400 | ~n8432;
  assign n8433 = ~P1_IR_REG_23__SCAN_IN;
  assign n13082 = ~n8434 ^ n8433;
  assign n8435 = n13082 & P1_STATE_REG_SCAN_IN;
  assign n9785 = n15009 | n14937;
  assign n14611 = ~n9785;
  assign n11671 = ~n11766 | ~n12016;
  assign n10752 = ~n11766;
  assign n11670 = ~n10752 | ~n11997;
  assign n14943 = n8472 & n14914;
  assign n12748 = ~n10992 & ~n12804;
  assign n12747 = ~n10992 | ~n12804;
  assign n13171 = ~n14646 | ~n8490;
  assign n13939 = ~n14639;
  assign n13081 = ~P1_STATE_REG_SCAN_IN;
  assign n9341 = ~n9338 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n9340 = ~n9339 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n10532 = ~n9341 | ~n9340;
  assign n14450 = ~P2_DATAO_REG_30__SCAN_IN;
  assign n12015 = ~n12357;
  assign n10534 = ~n10530 | ~SI_30_;
  assign n10533 = ~n10532 | ~n10531;
  assign n10541 = ~n10534 | ~n10533;
  assign n10538 = ~n10535 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n10537 = ~n10536 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n10539 = ~n10538 | ~n10537;
  assign n10540 = ~n10539 ^ SI_31_;
  assign n14463 = ~P2_DATAO_REG_31__SCAN_IN;
  assign n11188 = ~n7294 | ~P1_REG2_REG_31__SCAN_IN;
  assign n11187 = ~n8180 | ~P1_REG0_REG_31__SCAN_IN;
  assign n11191 = ~n11188 | ~n11187;
  assign n11189 = ~P1_REG1_REG_31__SCAN_IN;
  assign n11190 = ~n8105 & ~n11189;
  assign n14780 = ~n11191 & ~n11190;
  assign n14950 = ~n11671 | ~n11670;
  assign n14916 = ~n11767 | ~n12015;
  assign n14951 = ~n11768 | ~n14916;
  assign n14839 = ~n14825;
  assign n14960 = ~n14683 | ~n14839;
  assign n12749 = ~n12747;
  assign n14964 = ~n12749 & ~n12748;
  assign n14689 = ~n14683;
  assign n14902 = ~n13082 & ~n13081;
  assign n14966 = ~n13171;
  assign n14968 = ~n13331;
  assign n13934 = ~n14881;
  assign n14984 = ~n13934 | ~n14637;
  assign n14451 = n8304 | n14450;
  assign n14465 = ~n14462 | ~n14461;
  assign n14464 = n8304 | n14463;
  assign n14613 = ~n14612 | ~n14611;
  assign n14615 = ~n14614 & ~n14613;
  assign n14620 = ~n14616 | ~n14615;
  assign n15012 = ~n14902;
  assign n14794 = ~n14621;
  assign n14618 = ~n15012 & ~n14794;
  assign n14617 = ~P1_B_REG_SCAN_IN;
  assign n14619 = ~n14618 & ~n14617;
  assign n14896 = ~n14797 | ~n14780;
  assign n14934 = ~n14797 & ~n14780;
  assign n14799 = ~n14934;
  assign n15004 = ~n14896 | ~n14799;
  assign n14792 = n14621 & n14937;
  assign n14783 = ~n14792;
  assign n14625 = ~n14802 ^ n14783;
  assign n14623 = ~n14622;
  assign n14624 = ~n14802 | ~n14804;
  assign n14771 = ~n14625 | ~n14624;
  assign n14630 = ~n14771;
  assign n14626 = ~n14770 | ~n14783;
  assign n14627 = ~n14942 | ~n14626;
  assign n14629 = ~n14628 & ~n14627;
  assign n14776 = n14630 | n14629;
  assign n14738 = ~n14634;
  assign n14880 = ~n14632 | ~n14631;
  assign n14636 = ~n14880 & ~n14783;
  assign n14817 = ~n14634 | ~n14633;
  assign n14635 = ~n14817 & ~n14792;
  assign n14746 = ~n14636 & ~n14635;
  assign n14735 = ~n14743 | ~n14637;
  assign n14730 = ~n14638;
  assign n14641 = ~n14730 | ~n14783;
  assign n14731 = n14639 & n14792;
  assign n14640 = ~n14731;
  assign n14728 = ~n14641 | ~n14640;
  assign n14642 = ~n14823;
  assign n14643 = ~n14642 & ~n14783;
  assign n14713 = ~n14644 & ~n14643;
  assign n14849 = ~n14701 | ~n14646;
  assign n14697 = n14849 & n14792;
  assign n14648 = n14833 & n14671;
  assign n14647 = ~n14673;
  assign n14649 = ~n14648 & ~n14647;
  assign n14651 = ~n14649 | ~n14958;
  assign n14842 = n14666 & n14650;
  assign n14652 = ~n14651 | ~n14842;
  assign n14665 = ~n14652 | ~n14792;
  assign n14663 = ~n14792 | ~n14653;
  assign n14656 = ~n14832;
  assign n14829 = ~n14863 | ~n14917;
  assign n14655 = ~n14654 & ~n14829;
  assign n14661 = ~n14792 & ~n14657;
  assign n14659 = ~n14953;
  assign n14675 = ~n14958;
  assign n14658 = ~n14947 & ~n14675;
  assign n14660 = ~n14659 | ~n14658;
  assign n14664 = ~n14663 | ~n14662;
  assign n14669 = ~n14665 | ~n14664;
  assign n14667 = ~n14666;
  assign n14670 = ~n14667 | ~n14783;
  assign n14668 = n14840 & n14670;
  assign n14682 = ~n14669 | ~n14668;
  assign n14680 = ~n14670;
  assign n14674 = ~n14673 | ~n14672;
  assign n14827 = ~n14671 | ~n14674;
  assign n14677 = ~n14827 & ~n14675;
  assign n14826 = ~n14840 | ~n14676;
  assign n14678 = n14677 | n14826;
  assign n14679 = ~n14678 | ~n14783;
  assign n14681 = n14680 | n14679;
  assign n14686 = ~n14690 | ~n14683;
  assign n14684 = ~n14868;
  assign n14685 = n14684 & n14839;
  assign n14687 = n14686 & n14685;
  assign n14688 = ~n14687 & ~n14783;
  assign n14695 = ~n14688 | ~n14692;
  assign n14691 = ~n14825 & ~n14964;
  assign n14711 = ~n14700 & ~n14974;
  assign n14705 = ~n14702 | ~n14701;
  assign n14704 = ~n14703 | ~n14851;
  assign n14707 = ~n14705 | ~n14704;
  assign n14709 = ~n14707 | ~n14706;
  assign n14708 = ~n14853 & ~n14783;
  assign n14710 = ~n14709 | ~n14708;
  assign n14712 = ~n14711 | ~n14710;
  assign n14824 = ~n14714;
  assign n14718 = ~n14824 | ~n14783;
  assign n14717 = ~n14822 & ~n14783;
  assign n14876 = n7311 & n14715;
  assign n14716 = ~n14876 & ~n14792;
  assign n14720 = ~n14717 & ~n14716;
  assign n14719 = n14718 & n14720;
  assign n14721 = ~n14720;
  assign n14722 = n14721 | n14980;
  assign n14726 = ~n14729 | ~n14724;
  assign n14725 = ~n7311 & ~n14783;
  assign n14745 = ~n14728 | ~n14727;
  assign n14875 = ~n14730 | ~n14729;
  assign n14732 = ~n14731 | ~n14875;
  assign n14733 = ~n14745 | ~n14732;
  assign n14734 = ~n14881 & ~n14733;
  assign n14737 = ~n14746 & ~n14736;
  assign n14742 = ~n14884 & ~n14739;
  assign n14741 = ~n14740 | ~n14792;
  assign n14983 = ~n14744 | ~n14743;
  assign n14747 = ~n14746;
  assign n14749 = ~n14758;
  assign n14820 = ~n14749 & ~n14748;
  assign n14754 = ~n14752 | ~n14751;
  assign n14753 = ~n14888 | ~n14783;
  assign n14757 = ~n14754 | ~n14753;
  assign n14755 = n14813 & n14805;
  assign n14756 = n14755 & n14806;
  assign n14768 = ~n14757 | ~n14756;
  assign n14763 = ~n14806;
  assign n14759 = ~n14813 | ~n14758;
  assign n14760 = ~n14759 | ~n14792;
  assign n14762 = n14761 | n14760;
  assign n14766 = n14763 | n14762;
  assign n14764 = ~n14806 | ~n14805;
  assign n14765 = ~n14764 | ~n14783;
  assign n14767 = n14766 & n14765;
  assign n14769 = ~n14768 | ~n14767;
  assign n14774 = ~n14925 | ~n14769;
  assign n14889 = ~n8351 | ~n14925;
  assign n14772 = ~n14889 | ~n14792;
  assign n14773 = n14772 & n14771;
  assign n14775 = ~n14774 | ~n14773;
  assign n14779 = ~n14803 & ~n14792;
  assign n14778 = ~n14777 & ~n14783;
  assign n14941 = ~n14798;
  assign n14781 = ~n14941 & ~n14780;
  assign n14787 = ~n14940 | ~n14781;
  assign n14782 = ~n14786 | ~n14787;
  assign n14785 = n14940 | n14781;
  assign n14784 = ~n14782 | ~n14785;
  assign n14791 = ~n14784 | ~n14783;
  assign n14789 = ~n14788 | ~n14787;
  assign n14790 = ~n14789 | ~n14792;
  assign n14793 = ~n14934 | ~n14792;
  assign n14796 = ~n14795 ^ n14794;
  assign n14901 = ~n14796 | ~n14897;
  assign n14801 = ~n14798 | ~n14797;
  assign n14800 = ~n14799 | ~n14940;
  assign n14895 = ~n14801 | ~n14800;
  assign n14893 = n14801 | n14905;
  assign n14814 = ~n14803 | ~n14802;
  assign n14809 = ~n14804;
  assign n14807 = n14806 & n14805;
  assign n14808 = ~n14807 & ~n14889;
  assign n14810 = ~n14809 & ~n14808;
  assign n14811 = ~n14814 & ~n14810;
  assign n14907 = ~n14812 & ~n14811;
  assign n14815 = ~n14813;
  assign n14926 = ~n14815 & ~n14814;
  assign n14818 = ~n14884 & ~n14816;
  assign n14819 = ~n14818 | ~n14817;
  assign n14912 = ~n14820 | ~n14819;
  assign n14862 = ~n14822 | ~n14821;
  assign n14866 = ~n14824 & ~n14823;
  assign n14860 = ~n14866;
  assign n14828 = ~n14826 & ~n14825;
  assign n14864 = n14828 & n14827;
  assign n14830 = ~n14829;
  assign n14837 = ~n14831 | ~n14830;
  assign n14834 = ~n14833 | ~n14832;
  assign n14836 = ~n14835 & ~n14834;
  assign n14838 = ~n14837 | ~n14836;
  assign n14844 = ~n14864 | ~n14838;
  assign n14841 = ~n14840 | ~n14839;
  assign n14843 = n14842 | n14841;
  assign n14845 = ~n14844 | ~n14843;
  assign n14847 = ~n14846 & ~n14845;
  assign n14848 = ~n14868 & ~n14847;
  assign n14850 = ~n14849 & ~n14848;
  assign n14854 = ~n14851 | ~n14850;
  assign n14870 = ~n14853 & ~n14852;
  assign n14856 = ~n14854 | ~n14870;
  assign n14857 = ~n14856 | ~n14855;
  assign n14859 = ~n14858 & ~n14857;
  assign n14861 = ~n14860 & ~n14859;
  assign n14874 = ~n14862 & ~n14861;
  assign n14865 = n14864 & n14863;
  assign n14867 = ~n14866 | ~n14865;
  assign n14869 = ~n14868 & ~n14867;
  assign n14908 = ~n14870 | ~n14869;
  assign n14872 = ~n14908 & ~n14871;
  assign n14873 = ~n14875 & ~n14872;
  assign n14879 = ~n14874 | ~n14873;
  assign n14877 = ~n14876 & ~n14875;
  assign n14909 = ~n14878 & ~n14877;
  assign n14883 = ~n14879 | ~n14909;
  assign n14882 = ~n14881 & ~n14880;
  assign n14885 = ~n14883 | ~n14882;
  assign n14886 = ~n14885 & ~n14884;
  assign n14887 = ~n14912 & ~n14886;
  assign n14923 = ~n14888 & ~n14887;
  assign n14890 = ~n14889 & ~n14923;
  assign n14891 = ~n14926 | ~n14890;
  assign n14892 = ~n14907 | ~n14891;
  assign n14894 = ~n14893 | ~n14892;
  assign n14899 = ~n14895 | ~n14894;
  assign n14936 = ~n14896;
  assign n14898 = ~n14936 & ~n14897;
  assign n14900 = ~n14899 | ~n14898;
  assign n14904 = n14903 & n14902;
  assign n14932 = ~n14941 & ~n14905;
  assign n14906 = ~n14941 | ~n14905;
  assign n14930 = ~n14907 | ~n14906;
  assign n14910 = ~n14908;
  assign n14911 = ~n14910 | ~n14909;
  assign n14921 = ~n14912 & ~n14911;
  assign n14915 = ~n14913 & ~n15007;
  assign n14919 = ~n14915 | ~n14914;
  assign n14918 = ~n14917 | ~n14916;
  assign n14920 = ~n14919 & ~n14918;
  assign n14922 = ~n14921 | ~n14920;
  assign n14924 = ~n14923 | ~n14922;
  assign n14928 = ~n14925 | ~n14924;
  assign n14927 = ~n14926 | ~n14998;
  assign n14929 = ~n14928 & ~n14927;
  assign n14931 = ~n14930 & ~n14929;
  assign n14933 = ~n14932 & ~n14931;
  assign n14935 = ~n14934 & ~n14933;
  assign n14938 = ~n14936 & ~n14935;
  assign n15002 = ~n14941 ^ n14940;
  assign n14996 = ~n14942;
  assign n14945 = ~n14943;
  assign n14949 = ~n14945 & ~n14944;
  assign n14948 = ~n14947 & ~n14946;
  assign n14956 = ~n14949 | ~n14948;
  assign n14952 = ~n14950;
  assign n14954 = ~n14952 & ~n14951;
  assign n14955 = ~n14954 | ~n14659;
  assign n14957 = ~n14956 & ~n14955;
  assign n14959 = ~n14958 | ~n14957;
  assign n14961 = ~n14960 & ~n14959;
  assign n14963 = ~n14962 | ~n14961;
  assign n14965 = ~n14964 & ~n14963;
  assign n14970 = ~n14966 | ~n14965;
  assign n14969 = ~n14968 | ~n14967;
  assign n14971 = ~n14970 & ~n14969;
  assign n14973 = ~n14972 | ~n14971;
  assign n14975 = ~n14974 & ~n14973;
  assign n14977 = ~n14976 | ~n14975;
  assign n14979 = ~n14978 & ~n14977;
  assign n14981 = ~n14980 | ~n14979;
  assign n14986 = ~n14982 & ~n14981;
  assign n14985 = ~n14984 & ~n14983;
  assign n14987 = ~n14986 | ~n14985;
  assign n14989 = ~n14988 & ~n14987;
  assign n14991 = ~n14990 | ~n14989;
  assign n14993 = ~n14992 & ~n14991;
  assign n14995 = ~n14994 | ~n14993;
  assign n14997 = ~n14996 & ~n14995;
  assign n14999 = ~n14998 | ~n14997;
  assign n15001 = ~n15000 & ~n14999;
  assign n15003 = ~n15002 | ~n15001;
  assign n15006 = ~n15004 & ~n15003;
  assign n15008 = ~n15006 ^ n15005;
  assign n15010 = ~n15008 | ~n15007;
  assign n15011 = ~n15010 | ~n15009;
  assign input_0 = keyinput_0 ^ SI_31_;
  assign input_1 = keyinput_1 ^ SI_30_;
  assign AND_1 = input_0 & input_1;
  assign input_2 = ~keyinput_2 ^ SI_29_;
  assign OR_2 = input_2 | AND_1;
  assign input_3 = keyinput_3 ^ SI_28_;
  assign AND_3 = input_3 & OR_2;
  assign input_4 = ~keyinput_4 ^ SI_27_;
  assign OR_4 = input_4 | AND_3;
  assign input_5 = ~keyinput_5 ^ SI_26_;
  assign AND_5 = input_5 & OR_4;
  assign input_6 = ~keyinput_6 ^ SI_25_;
  assign AND_6 = input_6 & AND_5;
  assign input_7 = keyinput_7 ^ SI_24_;
  assign OR_7 = input_7 | AND_6;
  assign input_8 = keyinput_8 ^ SI_23_;
  assign AND_8 = input_8 & OR_7;
  assign input_9 = ~keyinput_9 ^ SI_22_;
  assign OR_9 = input_9 | AND_8;
  assign input_10 = keyinput_10 ^ SI_21_;
  assign AND_10 = input_10 & OR_9;
  assign input_11 = keyinput_11 ^ SI_20_;
  assign OR_11 = input_11 | AND_10;
  assign input_12 = keyinput_12 ^ SI_19_;
  assign AND_12 = input_12 & OR_11;
  assign input_13 = keyinput_13 ^ SI_18_;
  assign OR_13 = input_13 | AND_12;
  assign input_14 = keyinput_14 ^ SI_17_;
  assign AND_14 = input_14 & OR_13;
  assign input_15 = ~keyinput_15 ^ SI_16_;
  assign OR_15 = input_15 | AND_14;
  assign input_16 = keyinput_16 ^ SI_15_;
  assign OR_16 = input_16 | OR_15;
  assign input_17 = keyinput_17 ^ SI_14_;
  assign OR_17 = input_17 | OR_16;
  assign input_18 = ~keyinput_18 ^ SI_13_;
  assign AND_18 = input_18 & OR_17;
  assign input_19 = keyinput_19 ^ SI_12_;
  assign OR_19 = input_19 | AND_18;
  assign input_20 = keyinput_20 ^ SI_11_;
  assign OR_20 = input_20 | OR_19;
  assign input_21 = keyinput_21 ^ SI_10_;
  assign OR_21 = input_21 | OR_20;
  assign input_22 = keyinput_22 ^ SI_9_;
  assign AND_22 = input_22 & OR_21;
  assign input_23 = keyinput_23 ^ SI_8_;
  assign OR_23 = input_23 | AND_22;
  assign input_24 = keyinput_24 ^ SI_7_;
  assign OR_24 = input_24 | OR_23;
  assign input_25 = keyinput_25 ^ SI_6_;
  assign AND_25 = input_25 & OR_24;
  assign input_26 = ~keyinput_26 ^ SI_5_;
  assign AND_26 = input_26 & AND_25;
  assign input_27 = keyinput_27 ^ SI_4_;
  assign OR_27 = input_27 | AND_26;
  assign input_28 = ~keyinput_28 ^ SI_3_;
  assign OR_28 = input_28 | OR_27;
  assign input_29 = keyinput_29 ^ SI_2_;
  assign AND_29 = input_29 & OR_28;
  assign input_30 = keyinput_30 ^ SI_1_;
  assign AND_30 = input_30 & AND_29;
  assign input_31 = keyinput_31 ^ SI_0_;
  assign AND_31 = input_31 & AND_30;
  assign input_32 = ~keyinput_32 ^ P2_RD_REG_SCAN_IN;
  assign OR_32 = input_32 | AND_31;
  assign input_33 = ~keyinput_33 ^ P2_DATAO_REG_31__SCAN_IN;
  assign AND_33 = input_33 & OR_32;
  assign input_34 = ~keyinput_34 ^ P2_DATAO_REG_30__SCAN_IN;
  assign AND_34 = input_34 & AND_33;
  assign input_35 = keyinput_35 ^ P2_DATAO_REG_29__SCAN_IN;
  assign OR_35 = input_35 | AND_34;
  assign input_36 = ~keyinput_36 ^ P2_DATAO_REG_28__SCAN_IN;
  assign AND_36 = input_36 & OR_35;
  assign input_37 = ~keyinput_37 ^ P2_DATAO_REG_27__SCAN_IN;
  assign OR_37 = input_37 | AND_36;
  assign input_38 = keyinput_38 ^ P2_DATAO_REG_26__SCAN_IN;
  assign OR_38 = input_38 | OR_37;
  assign input_39 = ~keyinput_39 ^ P2_DATAO_REG_25__SCAN_IN;
  assign AND_39 = input_39 & OR_38;
  assign input_40 = ~keyinput_40 ^ P2_DATAO_REG_24__SCAN_IN;
  assign AND_40 = input_40 & AND_39;
  assign input_41 = keyinput_41 ^ P2_DATAO_REG_23__SCAN_IN;
  assign AND_41 = input_41 & AND_40;
  assign input_42 = keyinput_42 ^ P2_DATAO_REG_22__SCAN_IN;
  assign OR_42 = input_42 | AND_41;
  assign input_43 = keyinput_43 ^ P2_DATAO_REG_21__SCAN_IN;
  assign OR_43 = input_43 | OR_42;
  assign input_44 = keyinput_44 ^ P2_DATAO_REG_20__SCAN_IN;
  assign AND_44 = input_44 & OR_43;
  assign input_45 = keyinput_45 ^ P2_DATAO_REG_19__SCAN_IN;
  assign OR_45 = input_45 | AND_44;
  assign input_46 = ~keyinput_46 ^ P2_DATAO_REG_18__SCAN_IN;
  assign OR_46 = input_46 | OR_45;
  assign input_47 = keyinput_47 ^ P2_DATAO_REG_17__SCAN_IN;
  assign OR_47 = input_47 | OR_46;
  assign input_48 = ~keyinput_48 ^ P2_DATAO_REG_16__SCAN_IN;
  assign OR_48 = input_48 | OR_47;
  assign input_49 = ~keyinput_49 ^ P2_DATAO_REG_15__SCAN_IN;
  assign AND_49 = input_49 & OR_48;
  assign input_50 = ~keyinput_50 ^ P2_DATAO_REG_14__SCAN_IN;
  assign AND_50 = input_50 & AND_49;
  assign input_51 = ~keyinput_51 ^ P2_DATAO_REG_13__SCAN_IN;
  assign OR_51 = input_51 | AND_50;
  assign input_52 = ~keyinput_52 ^ P2_DATAO_REG_12__SCAN_IN;
  assign OR_52 = input_52 | OR_51;
  assign input_53 = keyinput_53 ^ P2_DATAO_REG_11__SCAN_IN;
  assign AND_53 = input_53 & OR_52;
  assign input_54 = keyinput_54 ^ P2_DATAO_REG_10__SCAN_IN;
  assign OR_54 = input_54 | AND_53;
  assign input_55 = ~keyinput_55 ^ P2_DATAO_REG_9__SCAN_IN;
  assign OR_55 = input_55 | OR_54;
  assign input_56 = ~keyinput_56 ^ P2_DATAO_REG_8__SCAN_IN;
  assign AND_56 = input_56 & OR_55;
  assign input_57 = ~keyinput_57 ^ P2_DATAO_REG_7__SCAN_IN;
  assign OR_57 = input_57 | AND_56;
  assign input_58 = keyinput_58 ^ P2_DATAO_REG_6__SCAN_IN;
  assign AND_58 = input_58 & OR_57;
  assign input_59 = keyinput_59 ^ P1_IR_REG_0__SCAN_IN;
  assign OR_59 = input_59 | AND_58;
  assign input_60 = keyinput_60 ^ P1_IR_REG_1__SCAN_IN;
  assign OR_60 = input_60 | OR_59;
  assign input_61 = keyinput_61 ^ P1_IR_REG_2__SCAN_IN;
  assign AND_61 = input_61 & OR_60;
  assign input_62 = ~keyinput_62 ^ P1_IR_REG_3__SCAN_IN;
  assign OR_62 = input_62 | AND_61;
  assign input_63 = ~keyinput_63 ^ P1_IR_REG_4__SCAN_IN;
  assign AND_63 = input_63 & OR_62;
  assign input_64 = ~keyinput_64 ^ P1_IR_REG_5__SCAN_IN;
  assign AND_64 = input_64 & AND_63;
  assign input_65 = ~keyinput_65 ^ P1_IR_REG_6__SCAN_IN;
  assign AND_65 = input_65 & AND_64;
  assign input_66 = ~keyinput_66 ^ P1_IR_REG_7__SCAN_IN;
  assign OR_66 = input_66 | AND_65;
  assign input_67 = ~keyinput_67 ^ P1_IR_REG_8__SCAN_IN;
  assign AND_67 = input_67 & OR_66;
  assign input_68 = ~keyinput_68 ^ P1_IR_REG_9__SCAN_IN;
  assign AND_68 = input_68 & AND_67;
  assign input_69 = ~keyinput_69 ^ P1_IR_REG_10__SCAN_IN;
  assign OR_69 = input_69 | AND_68;
  assign input_70 = ~keyinput_70 ^ P1_IR_REG_11__SCAN_IN;
  assign OR_70 = input_70 | OR_69;
  assign input_71 = ~keyinput_71 ^ P1_IR_REG_12__SCAN_IN;
  assign AND_71 = input_71 & OR_70;
  assign input_72 = keyinput_72 ^ P1_IR_REG_13__SCAN_IN;
  assign AND_72 = input_72 & AND_71;
  assign input_73 = ~keyinput_73 ^ P1_IR_REG_14__SCAN_IN;
  assign AND_73 = input_73 & AND_72;
  assign input_74 = ~keyinput_74 ^ P1_IR_REG_15__SCAN_IN;
  assign OR_74 = input_74 | AND_73;
  assign input_75 = keyinput_75 ^ P1_IR_REG_16__SCAN_IN;
  assign AND_75 = input_75 & OR_74;
  assign input_76 = ~keyinput_76 ^ P1_IR_REG_17__SCAN_IN;
  assign AND_76 = input_76 & AND_75;
  assign input_77 = ~keyinput_77 ^ P1_IR_REG_18__SCAN_IN;
  assign OR_77 = input_77 | AND_76;
  assign input_78 = keyinput_78 ^ P1_IR_REG_19__SCAN_IN;
  assign AND_78 = input_78 & OR_77;
  assign input_79 = keyinput_79 ^ P1_IR_REG_20__SCAN_IN;
  assign AND_79 = input_79 & AND_78;
  assign input_80 = keyinput_80 ^ SI_31_;
  assign input_81 = keyinput_81 ^ SI_30_;
  assign AND_81 = input_80 & input_81;
  assign input_82 = keyinput_82 ^ SI_29_;
  assign OR_82 = input_82 | AND_81;
  assign input_83 = ~keyinput_83 ^ SI_28_;
  assign AND_83 = input_83 & OR_82;
  assign input_84 = keyinput_84 ^ SI_27_;
  assign OR_84 = input_84 | AND_83;
  assign input_85 = keyinput_85 ^ SI_26_;
  assign AND_85 = input_85 & OR_84;
  assign input_86 = keyinput_86 ^ SI_25_;
  assign AND_86 = input_86 & AND_85;
  assign input_87 = keyinput_87 ^ SI_24_;
  assign OR_87 = input_87 | AND_86;
  assign input_88 = keyinput_88 ^ SI_23_;
  assign AND_88 = input_88 & OR_87;
  assign input_89 = keyinput_89 ^ SI_22_;
  assign OR_89 = input_89 | AND_88;
  assign input_90 = keyinput_90 ^ SI_21_;
  assign AND_90 = input_90 & OR_89;
  assign input_91 = ~keyinput_91 ^ SI_20_;
  assign OR_91 = input_91 | AND_90;
  assign input_92 = keyinput_92 ^ SI_19_;
  assign AND_92 = input_92 & OR_91;
  assign input_93 = keyinput_93 ^ SI_18_;
  assign OR_93 = input_93 | AND_92;
  assign input_94 = keyinput_94 ^ SI_17_;
  assign AND_94 = input_94 & OR_93;
  assign input_95 = ~keyinput_95 ^ SI_16_;
  assign OR_95 = input_95 | AND_94;
  assign input_96 = keyinput_96 ^ SI_15_;
  assign OR_96 = input_96 | OR_95;
  assign input_97 = ~keyinput_97 ^ SI_14_;
  assign OR_97 = input_97 | OR_96;
  assign input_98 = keyinput_98 ^ SI_13_;
  assign AND_98 = input_98 & OR_97;
  assign input_99 = ~keyinput_99 ^ SI_12_;
  assign OR_99 = input_99 | AND_98;
  assign input_100 = keyinput_100 ^ SI_11_;
  assign OR_100 = input_100 | OR_99;
  assign input_101 = keyinput_101 ^ SI_10_;
  assign OR_101 = input_101 | OR_100;
  assign input_102 = keyinput_102 ^ SI_9_;
  assign AND_102 = input_102 & OR_101;
  assign input_103 = ~keyinput_103 ^ SI_8_;
  assign OR_103 = input_103 | AND_102;
  assign input_104 = keyinput_104 ^ SI_7_;
  assign OR_104 = input_104 | OR_103;
  assign input_105 = keyinput_105 ^ SI_6_;
  assign AND_105 = input_105 & OR_104;
  assign input_106 = keyinput_106 ^ SI_5_;
  assign AND_106 = input_106 & AND_105;
  assign input_107 = keyinput_107 ^ SI_4_;
  assign OR_107 = input_107 | AND_106;
  assign input_108 = ~keyinput_108 ^ SI_3_;
  assign OR_108 = input_108 | OR_107;
  assign input_109 = keyinput_109 ^ SI_2_;
  assign AND_109 = input_109 & OR_108;
  assign input_110 = ~keyinput_110 ^ SI_1_;
  assign AND_110 = input_110 & AND_109;
  assign input_111 = keyinput_111 ^ SI_0_;
  assign AND_111 = input_111 & AND_110;
  assign input_112 = ~keyinput_112 ^ P2_RD_REG_SCAN_IN;
  assign OR_112 = input_112 | AND_111;
  assign input_113 = keyinput_113 ^ P2_DATAO_REG_31__SCAN_IN;
  assign AND_113 = input_113 & OR_112;
  assign input_114 = keyinput_114 ^ P2_DATAO_REG_30__SCAN_IN;
  assign AND_114 = input_114 & AND_113;
  assign input_115 = ~keyinput_115 ^ P2_DATAO_REG_29__SCAN_IN;
  assign OR_115 = input_115 | AND_114;
  assign input_116 = keyinput_116 ^ P2_DATAO_REG_28__SCAN_IN;
  assign AND_116 = input_116 & OR_115;
  assign input_117 = keyinput_117 ^ P2_DATAO_REG_27__SCAN_IN;
  assign OR_117 = input_117 | AND_116;
  assign input_118 = ~keyinput_118 ^ P2_DATAO_REG_26__SCAN_IN;
  assign OR_118 = input_118 | OR_117;
  assign input_119 = ~keyinput_119 ^ P2_DATAO_REG_25__SCAN_IN;
  assign AND_119 = input_119 & OR_118;
  assign input_120 = keyinput_120 ^ P2_DATAO_REG_24__SCAN_IN;
  assign AND_120 = input_120 & AND_119;
  assign input_121 = keyinput_121 ^ P2_DATAO_REG_23__SCAN_IN;
  assign AND_121 = input_121 & AND_120;
  assign input_122 = keyinput_122 ^ P2_DATAO_REG_22__SCAN_IN;
  assign OR_122 = input_122 | AND_121;
  assign input_123 = ~keyinput_123 ^ P2_DATAO_REG_21__SCAN_IN;
  assign OR_123 = input_123 | OR_122;
  assign input_124 = ~keyinput_124 ^ P2_DATAO_REG_20__SCAN_IN;
  assign AND_124 = input_124 & OR_123;
  assign input_125 = ~keyinput_125 ^ P2_DATAO_REG_19__SCAN_IN;
  assign OR_125 = input_125 | AND_124;
  assign input_126 = keyinput_126 ^ P2_DATAO_REG_18__SCAN_IN;
  assign OR_126 = input_126 | OR_125;
  assign input_127 = keyinput_127 ^ P2_DATAO_REG_17__SCAN_IN;
  assign OR_127 = input_127 | OR_126;
  assign input_128 = ~keyinput_128 ^ P2_DATAO_REG_16__SCAN_IN;
  assign OR_128 = input_128 | OR_127;
  assign input_129 = ~keyinput_129 ^ P2_DATAO_REG_15__SCAN_IN;
  assign AND_129 = input_129 & OR_128;
  assign input_130 = keyinput_130 ^ P2_DATAO_REG_14__SCAN_IN;
  assign AND_130 = input_130 & AND_129;
  assign input_131 = ~keyinput_131 ^ P2_DATAO_REG_13__SCAN_IN;
  assign OR_131 = input_131 | AND_130;
  assign input_132 = keyinput_132 ^ P2_DATAO_REG_12__SCAN_IN;
  assign OR_132 = input_132 | OR_131;
  assign input_133 = keyinput_133 ^ P2_DATAO_REG_11__SCAN_IN;
  assign AND_133 = input_133 & OR_132;
  assign input_134 = keyinput_134 ^ P2_DATAO_REG_10__SCAN_IN;
  assign OR_134 = input_134 | AND_133;
  assign input_135 = ~keyinput_135 ^ P2_DATAO_REG_9__SCAN_IN;
  assign OR_135 = input_135 | OR_134;
  assign input_136 = ~keyinput_136 ^ P2_DATAO_REG_8__SCAN_IN;
  assign AND_136 = input_136 & OR_135;
  assign input_137 = keyinput_137 ^ P2_DATAO_REG_7__SCAN_IN;
  assign OR_137 = input_137 | AND_136;
  assign input_138 = keyinput_138 ^ P2_DATAO_REG_6__SCAN_IN;
  assign AND_138 = input_138 & OR_137;
  assign input_139 = keyinput_139 ^ P1_IR_REG_0__SCAN_IN;
  assign OR_139 = input_139 | AND_138;
  assign input_140 = ~keyinput_140 ^ P1_IR_REG_1__SCAN_IN;
  assign OR_140 = input_140 | OR_139;
  assign input_141 = ~keyinput_141 ^ P1_IR_REG_2__SCAN_IN;
  assign AND_141 = input_141 & OR_140;
  assign input_142 = ~keyinput_142 ^ P1_IR_REG_3__SCAN_IN;
  assign OR_142 = input_142 | AND_141;
  assign input_143 = keyinput_143 ^ P1_IR_REG_4__SCAN_IN;
  assign AND_143 = input_143 & OR_142;
  assign input_144 = keyinput_144 ^ P1_IR_REG_5__SCAN_IN;
  assign AND_144 = input_144 & AND_143;
  assign input_145 = ~keyinput_145 ^ P1_IR_REG_6__SCAN_IN;
  assign AND_145 = input_145 & AND_144;
  assign input_146 = ~keyinput_146 ^ P1_IR_REG_7__SCAN_IN;
  assign OR_146 = input_146 | AND_145;
  assign input_147 = keyinput_147 ^ P1_IR_REG_8__SCAN_IN;
  assign AND_147 = input_147 & OR_146;
  assign input_148 = ~keyinput_148 ^ P1_IR_REG_9__SCAN_IN;
  assign AND_148 = input_148 & AND_147;
  assign input_149 = keyinput_149 ^ P1_IR_REG_10__SCAN_IN;
  assign OR_149 = input_149 | AND_148;
  assign input_150 = keyinput_150 ^ P1_IR_REG_11__SCAN_IN;
  assign OR_150 = input_150 | OR_149;
  assign input_151 = keyinput_151 ^ P1_IR_REG_12__SCAN_IN;
  assign AND_151 = input_151 & OR_150;
  assign input_152 = ~keyinput_152 ^ P1_IR_REG_13__SCAN_IN;
  assign AND_152 = input_152 & AND_151;
  assign input_153 = keyinput_153 ^ P1_IR_REG_14__SCAN_IN;
  assign AND_153 = input_153 & AND_152;
  assign input_154 = ~keyinput_154 ^ P1_IR_REG_15__SCAN_IN;
  assign OR_154 = input_154 | AND_153;
  assign input_155 = ~keyinput_155 ^ P1_IR_REG_16__SCAN_IN;
  assign AND_155 = input_155 & OR_154;
  assign input_156 = keyinput_156 ^ P1_IR_REG_17__SCAN_IN;
  assign AND_156 = input_156 & AND_155;
  assign input_157 = keyinput_157 ^ P1_IR_REG_18__SCAN_IN;
  assign OR_157 = input_157 | AND_156;
  assign input_158 = ~keyinput_158 ^ P1_IR_REG_19__SCAN_IN;
  assign AND_158 = input_158 & OR_157;
  assign input_159 = ~keyinput_159 ^ P1_IR_REG_20__SCAN_IN;
  assign AND_159 = input_159 & AND_158;
  assign AND_159_INV = ~AND_159;
  assign CASOP = AND_79 & AND_159_INV;
  assign P1_U3240 = P1_U3240_Lock ^ CASOP;
endmodule


