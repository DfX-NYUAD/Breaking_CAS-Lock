// Benchmark "b20_C_lock" written by ABC on Thu May 13 23:38:50 2021

module b20_C_lock ( 
    keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
    keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
    keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
    keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
    keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
    keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
    keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
    keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
    keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
    keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
    keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
    keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
    keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
    keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
    keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
    keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
    keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
    keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
    keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
    keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
    keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
    keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
    keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
    keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
    keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
    keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
    keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
    keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
    keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
    keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
    keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
    keyinput_156, keyinput_157, keyinput_158, keyinput_159, SI_31_, SI_30_,
    SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
    SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_,
    SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_,
    SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN,
    P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
    P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
    P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
    P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
    P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
    P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
    P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
    P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
    P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
    P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
    P1_IR_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
    P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
    P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
    P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    P1_U3242  );
  input  keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4,
    keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9,
    keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14,
    keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19,
    keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24,
    keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29,
    keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34,
    keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39,
    keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44,
    keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49,
    keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54,
    keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59,
    keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64,
    keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69,
    keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74,
    keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79,
    keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84,
    keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89,
    keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94,
    keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99,
    keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104,
    keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109,
    keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114,
    keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119,
    keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124,
    keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129,
    keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134,
    keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139,
    keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144,
    keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149,
    keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154,
    keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159,
    SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_,
    SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_,
    SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_,
    SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN,
    P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
    P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
    P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
    P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
    P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
    P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
    P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
    P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
    P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
    P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
    P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
    P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
    P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
    P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
    P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
    P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
    P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
    P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
    P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
    P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
    P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
    P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
    P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
    P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
    P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
    P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
    P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
    P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
    P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
    P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
    P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
    P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
    P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
    P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
    P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
    P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
    P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
    P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
    P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
    P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
    P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
    P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
    P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
    P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
    P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
    P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
    P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
    P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
    P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
    P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
    P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
    P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
    P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
    P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
    P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
    P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
    P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
    P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
    P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
    P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
    P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
    P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
    P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
    P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
    P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
    P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
    P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
    P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
    P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output P1_U3242;
  wire n9606, n8288, n7876, n9378, n15134, n13837, n14126, n13335, n14227,
    n14013, n14073, n14060, n11915, n9049, n7327, n9078, n9071, n7328,
    n13951, n13207, n9225, n7918, n7765, n9151, n9515, n7329, n7817, n7959,
    n7755, n7560, n7583, n7811, n10549, n10738, n7816, n8952, n7489, n7738,
    n7741, n10480, n8479, n7747, n7746, n10632, n7493, n7491, n7492, n7501,
    n7730, n7731, n7506, n7508, n7943, n7941, n10937, n10696, n10774,
    n7559, n7803, n7533, n7925, n7923, n7813, n7814, n7960, n8141, n8121,
    n8082, n9307, n8038, n7549, n8128, n15119, n14758, n7754, n13674,
    n8996, n8991, n7889, n7739, n7740, n7884, n7687, n8378, n7570, n7568,
    n8310, n7561, n8931, n7760, n7967, n7762, n9624, n7724, n7725, n7726,
    n10552, n10503, n9593, n14543, n14723, n14610, n14162, n9377, n8994,
    n8555, n8518, n8447, n9266, n8414, n9356, n7502, n7496, n10671, n7490,
    n7500, n7735, n7732, n7736, n7574, n10734, n7504, n10646, n7955, n7953,
    n8165, n7949, n7947, n10446, n10903, n7751, n7743, n7764, n7763, n8925,
    n8119, n7954, n8058, n7758, n8311, n8108, n8087, n7550, n8100, n7948,
    n10887, n13775, n13876, n7749, n7748, n7557, n7554, n7555, n7890,
    n7569, n7562, n7759, n8251, n8175, n8171, n7815, n7767, n7454, n15031,
    n13320, n11007, n7572, n13128, n14752, n12921, n13502, n13767, n12340,
    n14676, n14898, n15090, n14867, n14397, n13592, n13250, n13004, n12942,
    n12460, n11935, n7498, n9277, n11214, n7693, n8535, n11248, n8501,
    n8956, n7456, n8961, n9269, n8398, n9818, n8271, n11374, n7600, n7601,
    n7602, n9534, n7727, n7728, n7729, n10583, n7566, n11476, n13231,
    n12957, n13186, n12956, n12808, n10511, n10507, n14250, n8951, n13457,
    n7516, n7821, n8464, n8431, n7330, n9285, n7337, n7340, n7343, n7344,
    n7345, n7348, n7349, n7351, n9026, n8569, n9384, n7355, n7362, n7365,
    n7373, n12650, n10451, n7376, n7378, n7380, n11857, n13555, n7384,
    n7385, n7398, n10618, n7400, n14429, n7410, n7411, n7414, n7416,
    n10925, n7423, n7424, n7433, n7437, n12531, n7695, n7757, n7440, n8928,
    n7442, n7443, n7444, n7445, n7446, n7449, n7450, n7696, n7451, n12567,
    n10744, n7486, n7487, n7488, n7582, n10644, n7494, n7495, n7497,
    n10591, n10729, n7499, n10636, n7503, n7505, n7507, n7509, n7756,
    n7510, n7511, n7512, n7514, n7515, n8947, n8945, n7532, n7534, n7935,
    n11301, n7951, n11321, n7552, n8235, n7553, n7558, n7556, n7809, n7812,
    n8143, n7571, n8537, n7573, n7737, n7575, n9789, n7891, n7581, n7938,
    n9343, n7688, n8988, n12470, n8937, n7734, n7733, n7742, n7744, n7745,
    n7750, n7752, n7753, n10597, n10806, P1_U3242_Lock, n7761, n8212,
    n7766, n9514, n7961, n9327, n9345, n9519, n9535, n9553, n9572, n9597,
    n9628, n9655, n9686, n9715, n9744, n9767, n9794, n9819, n9846, n9869,
    n9275, n9308, n9288, n9287, n9742, n7885, n7900, n9721, n8929, n9076,
    n13237, n8169, n14856, n8953, n12357, n8503, n11612, n12815, n13561,
    n13957, n7905, n7904, n7970, n7971, n7907, n8497, n7906, n7969, n7909,
    n7908, n7966, n7968, n7911, n7910, n7964, n7965, n7913, n7912, n7914,
    n8213, n7916, n7915, n7917, n7963, n8195, n7920, n7919, n7921, n8176,
    n7922, n7962, n7924, n8047, n7927, n7926, n7929, n7928, n7933, n7930,
    n8026, n7931, n7932, n7934, n8059, n7936, n7937, n7939, n7940, n7942,
    n8080, n7945, n7944, n7946, n7950, n7952, n7956, n7957, n7958, n8234,
    n8250, n8270, n8287, n7973, n7972, n8308, n8309, n11905, n9763, n8039,
    n8060, n11289, n8081, n11316, n8101, n8120, n11025, n8142, n11274,
    n8170, n11306, n11347, n9567, n9594, n11415, n9622, n11512, n9651,
    n11672, n9678, n11743, n9711, n11828, n9738, n8312, n8314, n8313,
    n8333, n8332, n8331, n8356, n8357, n8334, n12119, n9816, n8355, n8354,
    n8377, n8379, n8358, n12295, n9840, n8376, n8375, n8397, n8399, n8380,
    n12426, n9867, n8401, n8400, n8413, n8415, n12727, n8416, n8418, n8417,
    n8430, n8432, n12849, n8433, n8435, n8434, n8446, n8448, n13040, n8449,
    n8451, n8450, n8463, n8465, n13171, n8467, n8466, n8478, n8480, n8482,
    n8481, n8484, n8483, n8500, n8502, n8499, n8498, n8517, n8519, n8504,
    n13464, n8520, n8522, n8521, n8534, n8536, n13658, n8538, n8540, n8539,
    n8554, n8556, n8553, n8552, n8572, n8574, n8558, n8557, n8573, n13943,
    n8571, n8570, n8577, n8594, n8576, n8575, n8593, n8579, n8578, n8584,
    n8581, n8580, n8582, n8583, n9376, n8926, n8927, n8930, n9680, n8932,
    n8933, n9842, n9268, n8934, n8958, n8935, n8944, n8936, n8938, n8940,
    n8949, n8939, n8941, n13338, n8943, n8942, n8946, n10960, P1_U3086,
    n8948, n8950, n8993, n8989, n8954, n8955, n12950, n8957, n8960, n8959,
    n8962, n12800, n11253, n8990, n8992, n11189, n11187, n9056, n9059,
    n11492, n9576, n12902, n8995, n8998, n9072, n8997, n9004, n9002, n8999,
    n9580, n9000, n9001, n9003, n9008, n9007, n9013, n9011, n9009, n9010,
    n9012, n12534, n9016, n9018, n9017, n9023, n9021, n9019, n9020, n9022,
    n9027, n9029, n9028, n9034, n9032, n9030, n9031, n9033, n12181, n9038,
    n9037, n9043, n9041, n9039, n9040, n9042, n10454, n9048, n9046, n9047,
    n9053, n9051, n9050, n9052, n9058, n9057, n9060, n12776, n9061, n9063,
    n9062, n9068, n9066, n9064, n9065, n9067, n9074, n9073, n9082, n9075,
    n9080, n9077, n9079, n9081, n11249, n9271, n9267, n9270, n14881, n9362,
    n9273, n9278, n9276, n9274, n11682, n11687, n12091, n9279, n9291,
    n9286, n11022, n12085, n10958, n9309, n9324, n11632, n11296, n9310,
    n9322, n9328, n9323, n9325, n9326, n11483, n11455, n9330, n9710, n9893,
    n9329, n12015, n9342, n9346, n9344, n11600, n11454, n9348, n9347,
    n12201, n10956, n10962, n9513, n9520, n9681, n9517, n9516, n9518,
    n11453, n9522, n9521, n9533, n9536, n9550, n11452, n11493, n9538,
    n9537, n9548, n9554, n9549, n9551, n9569, n9552, n11713, n11451, n9556,
    n9555, n12762, n9575, n9568, n9573, n9570, n9571, n11525, n9574, n9601,
    n12945, n9577, n9579, n9578, n9585, n9583, n9581, n9582, n9584, n9600,
    n9595, n9598, n9596, n11552, n11449, n9599, n11524, n9632, n12979,
    n9602, n9604, n9603, n9610, n9608, n9605, n9607, n9609, n9631, n9623,
    n9629, n9625, n9683, n9626, n9653, n9627, n11731, n11551, n9630, n9659,
    n13326, n9633, n9635, n9634, n9640, n9638, n9636, n9637, n9639, n9658,
    n9652, n9656, n9654, n11730, n9657, n9690, n13510, n9660, n9662, n9661,
    n9667, n9665, n9663, n9664, n9666, n9689, n9679, n9687, n9682, n9684,
    n9713, n9685, n12275, n11816, n9688, n9719, n13124, n9691, n9693,
    n9692, n9698, n9696, n9694, n9695, n9697, n9718, n9712, n9716, n9714,
    n12274, n9717, n9748, n13518, n9720, n9723, n9722, n9728, n9726, n9724,
    n9725, n9727, n9747, n9739, n9745, n9740, n9765, n9741, n9743, n13490,
    n12641, n9746, n9776, n13543, n9749, n9751, n9750, n9756, n9754, n9752,
    n9753, n9755, n9770, n9764, n9768, n9766, n13495, n9769, n9773, n9771,
    n9772, n9775, n9774, n9779, n9803, n14053, n9777, n9778, n13680, n9797,
    n9790, n9795, n9791, n9792, n9793, n14335, n13793, n9796, n9800, n9798,
    n9799, n9802, n9801, n9806, n9828, n14068, n9804, n9805, n13879, n9822,
    n9817, n9820, n9843, n14628, n14334, n9821, n9825, n9823, n9824, n9827,
    n9826, n9831, n9850, n14007, n9829, n9830, n13679, n9849, n9841, n9847,
    n9844, n9845, n14627, n9848, n9873, n13763, n9851, n9858, n9854, n9852,
    n9853, n9856, n9855, n9857, n14120, n9872, n9868, n9870, n9871, n9896,
    n14312, n9874, n9881, n9877, n9875, n9876, n9879, n9878, n9880, n14106,
    n9895, n12568, n9894, n9912, n14475, n9897, n9904, n9900, n9898, n9899,
    n9902, n9901, n9903, n14141, n9911, n12801, n9910, n9934, n14600,
    n9913, n9920, n9916, n9914, n9915, n9918, n9917, n9919, n14105, n9933,
    n12951, n9932, n9952, n14285, n9949, n9941, n9937, n9935, n9936, n9939,
    n9938, n9940, n14139, n10551, n10017, n14421, n10159, n9959, n9955,
    n9953, n9954, n9957, n9956, n9958, n11756, n10006, n13168, n10005,
    n10016, n13208, n10015, n10037, n14721, n10047, n10024, n10020, n10018,
    n10019, n10022, n10021, n10023, n11926, n10468, n10219, n14748, n10229,
    n10044, n10040, n10038, n10039, n10042, n10041, n10043, n12065, n10204,
    n10202, n10203, n10325, n14842, n10336, n10226, n10222, n10220, n10221,
    n10224, n10223, n10225, n12211, n10312, n13461, n10311, n10441, n10324,
    n10428, n15026, n10326, n10333, n10329, n10327, n10328, n10331, n10330,
    n10332, n12332, n13834, n10427, n10475, n15104, n10429, n10436, n10432,
    n10430, n10431, n10434, n10433, n10435, n12423, n10437, n10997, n10945,
    n10440, n10438, n10439, n10737, n10967, n10736, n10793, n10884, n10735,
    n14847, n10442, n10817, n10816, n10814, n10722, n10810, n10443, n10723,
    n14485, n10703, n10444, n10702, n10885, n10783, n10605, n10464, n10926,
    n10857, n10462, n10609, n10460, n10608, n10445, n10848, n13134, n10844,
    n10664, n10828, n10662, n10514, n10827, n12349, n10832, n10833, n10835,
    n10892, n10633, n11883, n11869, n12081, n12103, n10886, n10623, n10630,
    n11881, n10452, n11989, n10635, n10634, n11991, n11988, n10453, n12344,
    n12345, n10455, n10839, n12908, n10650, n12656, n10906, n12476, n10515,
    n10651, n10658, n10518, n10831, n12966, n10458, n10614, n13200, n10915,
    n10461, n10681, n10607, n10611, n13535, n10683, n10690, n10923, n10693,
    n10709, n10547, n10716, n14109, n10807, n10467, n10469, n10805, n10604,
    n10474, n13952, n10473, n15149, n15153, n10476, n10484, n10479, n10477,
    n10478, n10482, n10481, n10483, n12287, n10485, n10741, n10949, n10796,
    n10491, n10490, n10494, n10492, n10493, n11365, n12089, n12343, n13559,
    n13676, n10585, n10584, n14782, n14793, n10587, n10586, n10590, n10588,
    n10589, n11352, n14738, n10745, n10871, n10593, n11185, n10592, n14837,
    n10954, n10742, n10947, n10739, n10867, n10594, n10754, n10595, n10596,
    n10600, n10598, n10862, n10753, n10599, n10732, n10602, n10601, n10603,
    n10727, n10855, n10606, n10931, n10676, n10921, n10674, n10825, n10613,
    n10610, n10612, n10673, n10615, n10826, n10616, n10620, n10617, n10914,
    n10619, n10670, n10621, n10622, n10625, n10624, n10627, n10626, n10629,
    n10628, n10640, n10761, n10631, n10895, n10898, n10638, n10637, n10639,
    n10645, n10642, n10641, n10643, n10656, n10647, n10649, n10648, n10652,
    n10840, n10654, n10653, n10655, n10657, n10665, n10659, n10661, n10660,
    n10669, n10663, n10841, n10666, n10667, n10668, n10672, n10682, n10675,
    n10677, n10688, n10678, n10679, n10680, n10700, n10685, n10684, n10687,
    n10686, n10689, n10692, n10691, n10694, n10695, n10697, n10698, n10699,
    n10701, n10708, n10824, n10706, n10704, n10811, n10705, n10707, n10720,
    n10710, n10711, n10822, n10712, n10714, n10713, n10715, n10717, n10719,
    n10718, n10721, n10812, n10724, n10725, n10726, n10728, n10730, n10731,
    n10866, n10733, n10746, n10740, n10941, n10942, n10760, n10874, n10743,
    n10752, n10748, n10875, n10747, n10750, n10749, n10751, n10802, n10756,
    n10755, n10757, n10758, n10759, n10883, n10786, n10888, n11863, n10762,
    n10763, n12449, n10764, n10771, n10765, n10768, n10766, n10767, n10769,
    n10770, n10772, n10773, n10776, n10775, n10777, n10778, n10780, n10779,
    n10781, n10782, n10784, n10785, n10787, n10788, n10789, n10790, n10791,
    n10792, n10794, n10795, n10797, n10798, n10799, n10948, n10800, n10801,
    n10804, n10803, n10882, n10809, n10808, n10821, n10813, n10815, n10819,
    n10818, n10820, n10934, n10864, n10823, n10932, n10919, n10912, n10829,
    n10830, n10911, n10834, n10836, n10901, n10837, n10838, n10843, n10909,
    n10842, n10845, n10846, n10847, n10850, n10849, n10851, n10852, n10853,
    n10854, n10856, n10858, n10859, n10860, n10861, n10863, n10865, n10868,
    n10869, n10870, n10872, n10873, n10876, n10879, n10877, n10878, n10880,
    n10881, n10953, n10939, n10929, n10890, n10889, n10891, n10894, n10893,
    n10897, n10896, n10900, n10899, n10902, n10905, n10904, n10907, n10908,
    n10910, n10913, n10917, n10916, n10918, n10920, n10922, n10924, n10927,
    n10928, n10930, n10933, n10935, n10936, n10938, n10940, n10943, n10944,
    n10946, n10951, n10950, n10952, n10955, n10959, n10957, n10961, n13170,
    n11864, n10963, n11619, n10966, n10964, n10965, input_0, input_1,
    AND_1, input_2, AND_2, input_3, AND_3, input_4, OR_4, input_5, OR_5,
    input_6, OR_6, input_7, OR_7, input_8, OR_8, input_9, OR_9, input_10,
    AND_10, input_11, AND_11, input_12, OR_12, input_13, AND_13, input_14,
    OR_14, input_15, AND_15, input_16, AND_16, input_17, OR_17, input_18,
    OR_18, input_19, AND_19, input_20, AND_20, input_21, AND_21, input_22,
    AND_22, input_23, OR_23, input_24, OR_24, input_25, AND_25, input_26,
    AND_26, input_27, OR_27, input_28, OR_28, input_29, OR_29, input_30,
    AND_30, input_31, AND_31, input_32, OR_32, input_33, AND_33, input_34,
    AND_34, input_35, OR_35, input_36, OR_36, input_37, OR_37, input_38,
    AND_38, input_39, OR_39, input_40, OR_40, input_41, AND_41, input_42,
    OR_42, input_43, OR_43, input_44, OR_44, input_45, OR_45, input_46,
    OR_46, input_47, OR_47, input_48, AND_48, input_49, OR_49, input_50,
    OR_50, input_51, AND_51, input_52, AND_52, input_53, AND_53, input_54,
    AND_54, input_55, AND_55, input_56, OR_56, input_57, OR_57, input_58,
    AND_58, input_59, OR_59, input_60, OR_60, input_61, AND_61, input_62,
    OR_62, input_63, OR_63, input_64, AND_64, input_65, AND_65, input_66,
    AND_66, input_67, AND_67, input_68, AND_68, input_69, AND_69, input_70,
    AND_70, input_71, AND_71, input_72, OR_72, input_73, OR_73, input_74,
    AND_74, input_75, OR_75, input_76, AND_76, input_77, OR_77, input_78,
    AND_78, input_79, AND_79, input_80, input_81, AND_81, input_82, AND_82,
    input_83, AND_83, input_84, OR_84, input_85, OR_85, input_86, OR_86,
    input_87, OR_87, input_88, OR_88, input_89, OR_89, input_90, AND_90,
    input_91, AND_91, input_92, OR_92, input_93, AND_93, input_94, OR_94,
    input_95, AND_95, input_96, AND_96, input_97, OR_97, input_98, OR_98,
    input_99, AND_99, input_100, AND_100, input_101, AND_101, input_102,
    AND_102, input_103, OR_103, input_104, OR_104, input_105, AND_105,
    input_106, AND_106, input_107, OR_107, input_108, OR_108, input_109,
    OR_109, input_110, AND_110, input_111, AND_111, input_112, OR_112,
    input_113, AND_113, input_114, AND_114, input_115, OR_115, input_116,
    OR_116, input_117, OR_117, input_118, AND_118, input_119, OR_119,
    input_120, OR_120, input_121, AND_121, input_122, OR_122, input_123,
    OR_123, input_124, OR_124, input_125, OR_125, input_126, OR_126,
    input_127, OR_127, input_128, AND_128, input_129, OR_129, input_130,
    OR_130, input_131, AND_131, input_132, AND_132, input_133, AND_133,
    input_134, AND_134, input_135, AND_135, input_136, OR_136, input_137,
    OR_137, input_138, AND_138, input_139, OR_139, input_140, OR_140,
    input_141, AND_141, input_142, OR_142, input_143, OR_143, input_144,
    AND_144, input_145, AND_145, input_146, AND_146, input_147, AND_147,
    input_148, AND_148, input_149, AND_149, input_150, AND_150, input_151,
    AND_151, input_152, OR_152, input_153, OR_153, input_154, AND_154,
    input_155, OR_155, input_156, AND_156, input_157, OR_157, input_158,
    AND_158, input_159, AND_159, AND_159_INV, CASOP;
  assign n9606 = ~n9580;
  assign n8288 = n7562 & n7442;
  assign n7876 = ~n7328 | ~n11612;
  assign n9378 = ~n7918;
  assign n15134 = ~n11007;
  assign n13837 = n8555 ^ n8556;
  assign n14126 = ~n10783;
  assign n13335 = ~n8479 ^ n7821;
  assign n14227 = ~n9895 | ~n9894;
  assign n14013 = n9822 & n9821;
  assign n14073 = ~n9797 | ~n9796;
  assign n14060 = n9770 & n9769;
  assign n11915 = n9013 | n9012;
  assign n9049 = ~n9076;
  assign n7327 = ~n9026;
  assign n9078 = ~n8999 | ~n13951;
  assign n9071 = ~n13951 & ~n9377;
  assign n7328 = ~n7329;
  assign n13951 = ~n8996;
  assign n13207 = ~n7516 ^ n8936;
  assign n9225 = ~n8951 ^ n8989;
  assign n7918 = ~n9285;
  assign n7765 = n9307 & n7454;
  assign n9151 = ~P2_ADDR_REG_19__SCAN_IN ^ P1_ADDR_REG_19__SCAN_IN;
  assign n9515 = ~P1_IR_REG_5__SCAN_IN;
  assign n7329 = ~n9225;
  assign n7817 = ~n7960;
  assign n7959 = ~n7957 | ~n7755;
  assign n7755 = ~n7918 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n7560 = ~n8121 | ~n8119;
  assign n7583 = ~n7811 | ~n7936;
  assign n7811 = ~n8497 | ~P1_DATAO_REG_2__SCAN_IN;
  assign n10549 = ~n14610;
  assign n10738 = ~n11007 | ~n12423;
  assign n7816 = n8141 | n7817;
  assign n8952 = ~n7581 | ~P1_IR_REG_31__SCAN_IN;
  assign n7489 = n7884 & n8950;
  assign n7738 = ~n8378 | ~n7741;
  assign n7741 = ~n7743;
  assign n10480 = ~n9721;
  assign n8479 = ~n7746 | ~n7747;
  assign n7747 = ~n7748 & ~n7444;
  assign n7746 = ~n8447 | ~n7749;
  assign n10632 = ~n10622 | ~n7503;
  assign n7493 = ~n10668 | ~n10669;
  assign n7491 = ~n13134 & ~n7492;
  assign n7492 = ~n13200;
  assign n7501 = ~n7343 | ~n7423;
  assign n7730 = ~n7732 | ~n7731;
  assign n7731 = ~n10732;
  assign n7506 = ~n10867;
  assign n7508 = ~n10866;
  assign n7943 = ~n7941 | ~n7940;
  assign n7941 = n9285 | n8087;
  assign n10937 = ~n14752 & ~n12065;
  assign n10696 = n13767 | n14120;
  assign n10774 = n10461 | n10608;
  assign n7559 = ~n8416;
  assign n7803 = ~n7534 & ~n7532;
  assign n7533 = n9842 & n8933;
  assign n7925 = ~n7923 | ~n7922;
  assign n7923 = n8569 | n8165;
  assign n7813 = ~n7817 & ~n7814;
  assign n7814 = ~n7956;
  assign n7960 = ~n7959 | ~SI_6_;
  assign n8141 = ~n7959 ^ n7958;
  assign n8121 = ~n7951 | ~n7950;
  assign n8082 = ~n7939 | ~n7938;
  assign n9307 = ~P1_IR_REG_0__SCAN_IN & ~P1_IR_REG_1__SCAN_IN;
  assign n8038 = ~n7927 | ~n7926;
  assign n7549 = ~n7932 | ~n8026;
  assign n8128 = ~P1_DATAO_REG_5__SCAN_IN;
  assign n15119 = ~n10437 & ~n10945;
  assign n14758 = ~n7754 & ~n10937;
  assign n7754 = ~n10806;
  assign n13674 = n14060 & n13680;
  assign n8996 = ~n8991 ^ P1_IR_REG_29__SCAN_IN;
  assign n8991 = ~n8990 | ~P1_IR_REG_31__SCAN_IN;
  assign n7889 = n7890 & n8935;
  assign n7739 = ~n7740 & ~n7443;
  assign n7740 = ~n7743 & ~n8380;
  assign n7884 = n7688 & n7687;
  assign n7687 = n9680 & n8932;
  assign n8378 = ~n7570 | ~n8358;
  assign n7570 = ~n7569 | ~n7568;
  assign n7568 = ~n7571 & ~n8334;
  assign n8310 = ~n7561 & ~n7971;
  assign n7561 = ~n8288 & ~n8287;
  assign n8931 = ~n9624;
  assign n7760 = n7967 | n7968;
  assign n7967 = ~n8251 & ~n8250;
  assign n7762 = n7763 & n7963;
  assign n9624 = n9534 | n8927;
  assign n7724 = ~P2_ADDR_REG_19__SCAN_IN;
  assign n7725 = ~P1_RD_REG_SCAN_IN;
  assign n7726 = ~P2_RD_REG_SCAN_IN;
  assign n10552 = ~n14397;
  assign n10503 = ~n9034 & ~n9033;
  assign n9593 = n7876 & n9285;
  assign n14543 = n10006 & n10005;
  assign n14723 = ~n10016 | ~n10015;
  assign n14610 = n9911 & n9910;
  assign n14162 = ~n9872 | ~n9871;
  assign n9377 = ~n8994 ^ n11187;
  assign n8994 = ~n11189 | ~P1_IR_REG_31__SCAN_IN;
  assign n8555 = ~n8538 | ~n8537;
  assign n8518 = ~n8503 | ~n8504;
  assign n8447 = ~n7809 | ~n8433;
  assign n9266 = ~P1_IR_REG_20__SCAN_IN;
  assign n8414 = ~n7738 | ~n7739;
  assign n9356 = ~n8943 | ~n11248;
  assign n7502 = ~n10632 | ~n10631;
  assign n7496 = ~n10643 | ~n7337;
  assign n10671 = n7490 & n10670;
  assign n7490 = ~n7493 | ~n7491;
  assign n7500 = ~n7501 | ~n10724;
  assign n7735 = ~n10941 & ~n10731;
  assign n7732 = ~n10941;
  assign n7736 = ~n7737 | ~n7380;
  assign n7574 = ~n10740 & ~n10945;
  assign n10734 = n7505 & n7504;
  assign n7504 = ~n10947;
  assign n10646 = ~n10446;
  assign n7955 = ~n7953 | ~n7952;
  assign n7953 = n9378 | n8128;
  assign n8165 = ~P1_DATAO_REG_7__SCAN_IN;
  assign n7949 = ~n7947 | ~n7946;
  assign n7947 = n9384 | n8108;
  assign n10446 = ~n10903 | ~n12349;
  assign n10903 = ~n7696 | ~n7695;
  assign n7751 = ~n7752 | ~n8465;
  assign n7743 = ~n7744 | ~n8399;
  assign n7764 = n8195 & n7351;
  assign n7763 = ~n7764 | ~n8176;
  assign n8925 = ~P1_IR_REG_8__SCAN_IN;
  assign n8119 = ~n7955 ^ n7954;
  assign n7954 = ~SI_5_;
  assign n8058 = ~n7583 ^ n7937;
  assign n7758 = n8311 | n8312;
  assign n8311 = ~n8310 & ~n8309;
  assign n8108 = ~P1_DATAO_REG_4__SCAN_IN;
  assign n8087 = ~P1_DATAO_REG_3__SCAN_IN;
  assign n7550 = ~n7945 | ~n7944;
  assign n8100 = ~n7949 ^ n7948;
  assign n7948 = ~SI_4_;
  assign n10887 = ~n12800;
  assign n13775 = n10696 & n10605;
  assign n13876 = n10693 & n10464;
  assign n7749 = ~n7751;
  assign n7748 = ~n7751 & ~n8449;
  assign n7557 = n8415 | n7559;
  assign n7554 = ~n7555 & ~n7559;
  assign n7555 = ~n7739;
  assign n7890 = ~n8934 & ~P1_IR_REG_21__SCAN_IN;
  assign n7569 = ~n7758 | ~n7440;
  assign n7562 = ~n7760 | ~n7759;
  assign n7759 = ~n8270;
  assign n8251 = ~n7552 & ~n7965;
  assign n8175 = ~n7962 | ~n7961;
  assign n8171 = ~n7815 | ~n7960;
  assign n7815 = ~n8143 | ~n8141;
  assign n7767 = ~P1_IR_REG_4__SCAN_IN;
  assign n7454 = ~P1_IR_REG_2__SCAN_IN & ~P1_IR_REG_3__SCAN_IN;
  assign n15031 = n10440 & n10439;
  assign n13320 = n9631 & n9630;
  assign n11007 = n7572 & n10427;
  assign n7572 = ~n13837 | ~n9893;
  assign n13128 = n9689 & n9688;
  assign n14752 = n10204 & n10203;
  assign n12921 = n9600 & n9599;
  assign n13502 = n9658 & n9657;
  assign n13767 = n9849 & n9848;
  assign n12340 = ~n9068 & ~n9067;
  assign n14676 = ~n10604;
  assign n14898 = ~n14881;
  assign n15090 = ~n15031;
  assign n14867 = ~n10312 | ~n10311;
  assign n14397 = ~n9933 | ~n9932;
  assign n13592 = n9747 & n9746;
  assign n13250 = ~n9718 | ~n9717;
  assign n13004 = ~n13320;
  assign n12942 = ~n9575 | ~n9574;
  assign n12460 = n9522 & n9521;
  assign n11935 = ~n7373 | ~n7498;
  assign n7498 = n10591 | n9310;
  assign n9277 = n9276 & n9275;
  assign n11214 = n9356 & n11249;
  assign n7693 = n7891 & n7385;
  assign n8535 = ~n7573 & ~n8520;
  assign n11248 = ~n8942 ^ P1_IR_REG_26__SCAN_IN;
  assign n8501 = ~n8482 | ~n8481;
  assign n8956 = n7891 & n7456;
  assign n7456 = ~n8934;
  assign n8961 = ~n7891 | ~n7890;
  assign n9269 = n7891 | n9681;
  assign n8398 = ~n7742 | ~n8380;
  assign n9818 = ~n7884 | ~n8931;
  assign n8271 = ~n7760;
  assign n11374 = ~n7601 ^ n7600;
  assign n7600 = ~n8195;
  assign n7601 = ~n7602 | ~n7351;
  assign n7602 = n8175 | n8176;
  assign n9534 = ~n7765 | ~n7355;
  assign n7727 = ~n7729 | ~n7728;
  assign n7728 = ~n7726 | ~P1_ADDR_REG_19__SCAN_IN;
  assign n7729 = ~n7725 | ~n7724;
  assign n10583 = ~n9376;
  assign n7566 = ~n7330 & ~n7362;
  assign n11476 = n9728 | n9727;
  assign n13231 = n9698 | n9697;
  assign n12957 = n9667 | n9666;
  assign n13186 = n9640 | n9639;
  assign n12956 = n9610 | n9609;
  assign n12808 = n9585 | n9584;
  assign n10511 = n9004 | n9003;
  assign n10507 = ~n12340;
  assign n14250 = ~n8584 ^ n8583;
  assign n8951 = ~n8953 | ~P1_IR_REG_31__SCAN_IN;
  assign n13457 = n8501 ^ n8502;
  assign n7516 = ~n7514 | ~P1_IR_REG_31__SCAN_IN;
  assign n7821 = ~n8480;
  assign n8464 = ~n7750 | ~n8449;
  assign n8431 = ~n7556 | ~n8416;
  assign n7330 = n7344 & n12567;
  assign n9285 = n9151 & n7727;
  assign n7337 = n7497 & n10651;
  assign n7340 = n10633 & n10753;
  assign n7343 = n10715 & n10722;
  assign n7344 = n10957 | n10956;
  assign n7345 = n10759 | n12800;
  assign n7348 = n9680 & n8929;
  assign n7349 = n7348 & n7446;
  assign n7351 = SI_8_ | n7921;
  assign n9026 = ~n9071;
  assign n8569 = ~n8497;
  assign n9384 = ~n8497;
  assign n7355 = n7767 & n9515;
  assign n7362 = ~n10961 | ~n13170;
  assign n7365 = n8944 & n8936;
  assign n7373 = n9309 & n9308;
  assign n12650 = n10651 & n10827;
  assign n10451 = ~n9053 & ~n9052;
  assign n7376 = n7569 & n7757;
  assign n7378 = n7889 & n7365;
  assign n7380 = n10741 & n10754;
  assign n11857 = ~n9082 & ~n9081;
  assign n13555 = n13674 | n10683;
  assign n7384 = n7378 & n8949;
  assign n7385 = n8948 & n8989;
  assign n7398 = n7693 & n7384;
  assign n10618 = n13128 & n13231;
  assign n7400 = ~n7891 | ~n7378;
  assign n14429 = n10467 | n10816;
  assign n7410 = SI_10_ | n7914;
  assign n7411 = n10801 | n10887;
  assign n7414 = n7816 & n8169;
  assign n7416 = n7494 & n10827;
  assign n10925 = n14073 & n10462;
  assign n7423 = ~n10721 | ~n10720;
  assign n7424 = n7511 & n7344;
  assign n7433 = ~n10650 | ~n10903;
  assign n7437 = n7885 & n8929;
  assign n12531 = ~n9538 | ~n9537;
  assign n7695 = ~n12531;
  assign n7757 = ~n8334;
  assign n7440 = SI_16_ ^ n8333;
  assign n8928 = ~n8927;
  assign n7442 = SI_13_ | n7969;
  assign n7443 = SI_19_ & n8397;
  assign n7444 = SI_23_ & n8463;
  assign n7445 = n8931 & n7349;
  assign n7446 = n8930 & n7885;
  assign n7449 = n7557 & n8432;
  assign n7450 = n7348 & n8930;
  assign n7696 = n9022 | n9023;
  assign n7451 = n10966 | n10965;
  assign n12567 = ~n9267 ^ n9266;
  assign n10744 = ~n7486 | ~n10742;
  assign n7486 = ~n7487 | ~n10874;
  assign n7487 = ~n7488 | ~n7736;
  assign n7488 = ~n10746;
  assign n7582 = n7489 & n7803;
  assign n10644 = ~n7496 | ~n7416;
  assign n7494 = ~n7337 | ~n7495;
  assign n7495 = ~n10906;
  assign n7497 = ~n7433 | ~n10906;
  assign n10591 = ~n7876 | ~n7918;
  assign n10729 = ~n7499 | ~n10727;
  assign n7499 = ~n7500 | ~n10726;
  assign n10636 = ~n7502 | ~n10895;
  assign n7503 = ~n7340 | ~n10630;
  assign n7505 = ~n7507 | ~n7506;
  assign n7507 = ~n7509 | ~n7508;
  assign n7509 = ~n10731 | ~n10732;
  assign n7756 = ~n7510 | ~n7566;
  assign n7510 = ~n7512 | ~n7424;
  assign n7511 = ~n10882 | ~n10881;
  assign n7512 = ~n7345 | ~n7411;
  assign n7514 = ~n7515 | ~n8944;
  assign n7515 = ~n8937;
  assign n8947 = ~n8945 | ~n8944;
  assign n8945 = ~n8937 | ~P1_IR_REG_31__SCAN_IN;
  assign n7532 = ~n7533 | ~n7355;
  assign n7534 = ~n8928 | ~n7765;
  assign n7935 = ~n7933 | ~n7549;
  assign n11301 = ~n8039 ^ n7549;
  assign n7951 = ~n7550 | ~n8100;
  assign n11321 = ~n7550 ^ n8101;
  assign n7552 = ~n8235 & ~n8234;
  assign n8235 = n7553 & n7410;
  assign n7553 = n8212 | n8213;
  assign n7558 = ~n7738 | ~n7554;
  assign n7556 = ~n8414 | ~n8415;
  assign n7809 = ~n7558 | ~n7449;
  assign n7812 = ~n7560 | ~n7813;
  assign n8143 = ~n7560 | ~n7956;
  assign n7571 = ~n8357;
  assign n8537 = ~n8535 | ~n8536;
  assign n7573 = ~n8519 & ~n8518;
  assign n7737 = ~n7575 | ~n7574;
  assign n7575 = ~n7733 | ~n7730;
  assign n9789 = ~n7758 ^ n7440;
  assign n7891 = n7803 & n7884;
  assign n7581 = ~n7582 | ~n7378;
  assign n7938 = ~n7583 | ~SI_2_;
  assign n9343 = ~n7765;
  assign n7688 = n7437 & n8930;
  assign n8988 = ~n7384 | ~n7891;
  assign n12470 = ~n7696;
  assign n8937 = ~n7891 | ~n7889;
  assign n7734 = ~n10738 | ~n10737;
  assign n7733 = ~n7735 & ~n7734;
  assign n7742 = ~n8378 | ~n8379;
  assign n7744 = n8379 | n7745;
  assign n7745 = ~n8380;
  assign n7750 = ~n8447 | ~n8448;
  assign n7752 = n8448 | n7753;
  assign n7753 = ~n8449;
  assign n10597 = ~n14758 | ~n10594;
  assign n10806 = ~n14752 | ~n12065;
  assign P1_U3242_Lock = ~n7756 | ~n7451;
  assign n7761 = ~n8175 | ~n7764;
  assign n8212 = ~n7761 | ~n7762;
  assign n7766 = ~n7765 | ~n7767;
  assign n9514 = ~n7766 | ~P1_IR_REG_31__SCAN_IN;
  assign n7961 = ~n7812 | ~n7414;
  assign n9327 = n7876 | n11455;
  assign n9345 = n7876 | n11454;
  assign n9519 = n7876 | n11453;
  assign n9535 = n7876 | n11493;
  assign n9553 = n7876 | n11451;
  assign n9572 = n7876 | n11525;
  assign n9597 = n7876 | n11449;
  assign n9628 = n7876 | n11551;
  assign n9655 = n7876 | n11730;
  assign n9686 = n7876 | n11816;
  assign n9715 = n7876 | n12274;
  assign n9744 = n7876 | n12641;
  assign n9767 = n7876 | n13495;
  assign n9794 = n7876 | n13793;
  assign n9819 = n7876 | n14334;
  assign n9846 = n7876 | n14627;
  assign n9869 = n7876 | n14881;
  assign n9275 = n7876 | n11687;
  assign n9308 = n7876 | n11296;
  assign n9288 = n7876 | n9291;
  assign n9287 = ~n7876 | ~n11022;
  assign n9742 = ~n8931 | ~n7450;
  assign n7885 = ~P1_IR_REG_14__SCAN_IN;
  assign n7900 = n8993 & n8992;
  assign n9721 = ~n9072;
  assign n8929 = ~P1_IR_REG_13__SCAN_IN;
  assign n9076 = ~n13951 | ~n9377;
  assign n13237 = ~n10774;
  assign n8169 = ~n7925 ^ n7924;
  assign n14856 = ~n14867;
  assign n8953 = ~n8952 | ~n8993;
  assign n12357 = n10903 & n10835;
  assign n8503 = ~n8502 | ~n8501;
  assign n11612 = ~n8954 | ~n8953;
  assign n12815 = n10828 & n10662;
  assign n13561 = n9756 | n9755;
  assign n13957 = ~n13943;
  assign n7905 = ~n7918 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n7904 = ~n9378 | ~P2_DATAO_REG_14__SCAN_IN;
  assign n7970 = ~n7905 | ~n7904;
  assign n7971 = ~SI_14_ & ~n7970;
  assign n7907 = ~n7918 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n8497 = ~n9285;
  assign n7906 = ~n8569 | ~P2_DATAO_REG_13__SCAN_IN;
  assign n7969 = ~n7907 | ~n7906;
  assign n7909 = ~n7918 | ~P1_DATAO_REG_12__SCAN_IN;
  assign n7908 = ~n8569 | ~P2_DATAO_REG_12__SCAN_IN;
  assign n7966 = ~n7909 | ~n7908;
  assign n7968 = ~SI_12_ & ~n7966;
  assign n7911 = ~n7918 | ~P1_DATAO_REG_11__SCAN_IN;
  assign n7910 = ~n8569 | ~P2_DATAO_REG_11__SCAN_IN;
  assign n7964 = ~n7911 | ~n7910;
  assign n7965 = ~SI_11_ & ~n7964;
  assign n7913 = ~n7918 | ~P1_DATAO_REG_10__SCAN_IN;
  assign n7912 = ~n8569 | ~P2_DATAO_REG_10__SCAN_IN;
  assign n7914 = ~n7913 | ~n7912;
  assign n8213 = ~SI_10_ ^ n7914;
  assign n7916 = ~n7918 | ~P1_DATAO_REG_9__SCAN_IN;
  assign n7915 = ~n9378 | ~P2_DATAO_REG_9__SCAN_IN;
  assign n7917 = ~n7916 | ~n7915;
  assign n7963 = ~SI_9_ | ~n7917;
  assign n8195 = SI_9_ ^ n7917;
  assign n7920 = ~n7918 | ~P1_DATAO_REG_8__SCAN_IN;
  assign n7919 = ~n9378 | ~P2_DATAO_REG_8__SCAN_IN;
  assign n7921 = ~n7920 | ~n7919;
  assign n8176 = ~SI_8_ ^ n7921;
  assign n7922 = ~n9378 | ~P2_DATAO_REG_7__SCAN_IN;
  assign n7962 = ~SI_7_ | ~n7925;
  assign n7924 = ~SI_7_;
  assign n8047 = ~P1_DATAO_REG_1__SCAN_IN;
  assign n7927 = n9285 | n8047;
  assign n7926 = ~n9285 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n7929 = ~n8038;
  assign n7928 = ~SI_1_;
  assign n7933 = ~n7929 | ~n7928;
  assign n7930 = ~SI_0_ | ~P1_DATAO_REG_0__SCAN_IN;
  assign n8026 = n9285 | n7930;
  assign n7931 = SI_0_ & P2_DATAO_REG_0__SCAN_IN;
  assign n7932 = ~n9285 | ~n7931;
  assign n7934 = ~n8038 | ~SI_1_;
  assign n8059 = ~n7935 | ~n7934;
  assign n7936 = ~n9285 | ~P2_DATAO_REG_2__SCAN_IN;
  assign n7937 = ~SI_2_;
  assign n7939 = ~n8059 | ~n8058;
  assign n7940 = ~n9285 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n7942 = ~SI_3_;
  assign n8080 = ~n7943 ^ n7942;
  assign n7945 = ~n8082 | ~n8080;
  assign n7944 = ~n7943 | ~SI_3_;
  assign n7946 = ~n9378 | ~P2_DATAO_REG_4__SCAN_IN;
  assign n7950 = ~n7949 | ~SI_4_;
  assign n7952 = ~n8569 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n7956 = ~n7955 | ~SI_5_;
  assign n7957 = ~n9378 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n7958 = ~SI_6_;
  assign n8234 = ~SI_11_ ^ n7964;
  assign n8250 = ~SI_12_ ^ n7966;
  assign n8270 = ~SI_13_ ^ n7969;
  assign n8287 = ~SI_14_ ^ n7970;
  assign n7973 = ~n7918 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n7972 = ~n9384 | ~P2_DATAO_REG_15__SCAN_IN;
  assign n8308 = ~n7973 | ~n7972;
  assign n8309 = ~SI_15_ ^ n8308;
  assign n11905 = n8310 ^ n8309;
  assign n9763 = ~n11905;
  assign n8039 = ~n8038 ^ SI_1_;
  assign n8060 = ~n8058;
  assign n11289 = ~n8060 ^ n8059;
  assign n8081 = ~n8080;
  assign n11316 = ~n8082 ^ n8081;
  assign n8101 = ~n8100;
  assign n8120 = ~n8119;
  assign n11025 = ~n8121 ^ n8120;
  assign n8142 = ~n8141;
  assign n11274 = ~n8143 ^ n8142;
  assign n8170 = ~n8169;
  assign n11306 = ~n8171 ^ n8170;
  assign n11347 = n8176 ^ n8175;
  assign n9567 = ~n11347;
  assign n9594 = ~n11374;
  assign n11415 = n8213 ^ n8212;
  assign n9622 = ~n11415;
  assign n11512 = n8235 ^ n8234;
  assign n9651 = ~n11512;
  assign n11672 = n8251 ^ n8250;
  assign n9678 = ~n11672;
  assign n11743 = n8271 ^ n8270;
  assign n9711 = ~n11743;
  assign n11828 = n8288 ^ n8287;
  assign n9738 = ~n11828;
  assign n8312 = ~SI_15_ & ~n8308;
  assign n8314 = ~n7918 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n8313 = ~n9378 | ~P2_DATAO_REG_16__SCAN_IN;
  assign n8333 = ~n8314 | ~n8313;
  assign n8332 = ~n7918 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n8331 = ~n9384 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n8356 = ~n8332 | ~n8331;
  assign n8357 = SI_17_ ^ n8356;
  assign n8334 = ~SI_16_ & ~n8333;
  assign n12119 = ~n8357 ^ n7376;
  assign n9816 = ~n12119;
  assign n8355 = ~n7918 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n8354 = ~n9378 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n8377 = ~n8355 | ~n8354;
  assign n8379 = SI_18_ ^ n8377;
  assign n8358 = ~SI_17_ | ~n8356;
  assign n12295 = ~n8379 ^ n8378;
  assign n9840 = ~n12295;
  assign n8376 = ~n7918 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n8375 = ~n8569 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n8397 = ~n8376 | ~n8375;
  assign n8399 = SI_19_ ^ n8397;
  assign n8380 = ~SI_18_ | ~n8377;
  assign n12426 = ~n8399 ^ n8398;
  assign n9867 = ~n12426;
  assign n8401 = ~n7918 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n8400 = ~n8569 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n8413 = ~n8401 | ~n8400;
  assign n8415 = SI_20_ ^ n8413;
  assign n12727 = n8414 ^ n8415;
  assign n8416 = ~SI_20_ | ~n8413;
  assign n8418 = ~n7918 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n8417 = ~n8569 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n8430 = ~n8418 | ~n8417;
  assign n8432 = SI_21_ ^ n8430;
  assign n12849 = n8431 ^ n8432;
  assign n8433 = ~SI_21_ | ~n8430;
  assign n8435 = ~n7918 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n8434 = ~n9384 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n8446 = ~n8435 | ~n8434;
  assign n8448 = SI_22_ ^ n8446;
  assign n13040 = n8447 ^ n8448;
  assign n8449 = ~SI_22_ | ~n8446;
  assign n8451 = ~n7918 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n8450 = ~n9378 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n8463 = ~n8451 | ~n8450;
  assign n8465 = SI_23_ ^ n8463;
  assign n13171 = n8464 ^ n8465;
  assign n8467 = ~n7918 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n8466 = ~n9384 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n8478 = ~n8467 | ~n8466;
  assign n8480 = SI_24_ ^ n8478;
  assign n8482 = ~SI_24_ | ~n8478;
  assign n8481 = ~n8480 | ~n8479;
  assign n8484 = ~n8497 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n8483 = ~n9384 | ~P2_DATAO_REG_25__SCAN_IN;
  assign n8500 = ~n8484 | ~n8483;
  assign n8502 = SI_25_ ^ n8500;
  assign n8499 = ~n8497 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n8498 = ~n9384 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n8517 = ~n8499 | ~n8498;
  assign n8519 = ~SI_26_ ^ n8517;
  assign n8504 = ~SI_25_ | ~n8500;
  assign n13464 = ~n8519 ^ n8518;
  assign n8520 = ~SI_26_ & ~n8517;
  assign n8522 = ~n7918 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n8521 = ~n9378 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n8534 = ~n8522 | ~n8521;
  assign n8536 = SI_27_ ^ n8534;
  assign n13658 = n8535 ^ n8536;
  assign n8538 = ~SI_27_ | ~n8534;
  assign n8540 = ~n8497 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n8539 = ~n8569 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n8554 = ~n8540 | ~n8539;
  assign n8556 = SI_28_ ^ n8554;
  assign n8553 = ~n8497 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n8552 = ~n8569 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n8572 = ~n8553 | ~n8552;
  assign n8574 = SI_29_ ^ n8572;
  assign n8558 = ~SI_28_ | ~n8554;
  assign n8557 = ~n8556 | ~n8555;
  assign n8573 = ~n8558 | ~n8557;
  assign n13943 = ~n8574 ^ n8573;
  assign n8571 = ~n7918 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n8570 = ~n8569 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n8577 = ~n8571 | ~n8570;
  assign n8594 = SI_30_ ^ n8577;
  assign n8576 = ~SI_29_ | ~n8572;
  assign n8575 = ~n8574 | ~n8573;
  assign n8593 = ~n8576 | ~n8575;
  assign n8579 = ~n8594 | ~n8593;
  assign n8578 = ~SI_30_ | ~n8577;
  assign n8584 = ~n8579 | ~n8578;
  assign n8581 = ~n7918 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n8580 = ~n9384 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n8582 = ~n8581 | ~n8580;
  assign n8583 = ~n8582 ^ SI_31_;
  assign n9376 = ~n8594 ^ n8593;
  assign n8926 = ~P1_IR_REG_6__SCAN_IN & ~P1_IR_REG_7__SCAN_IN;
  assign n8927 = ~n8926 | ~n8925;
  assign n8930 = ~P1_IR_REG_9__SCAN_IN & ~P1_IR_REG_12__SCAN_IN;
  assign n9680 = ~P1_IR_REG_10__SCAN_IN & ~P1_IR_REG_11__SCAN_IN;
  assign n8932 = ~P1_IR_REG_15__SCAN_IN & ~P1_IR_REG_16__SCAN_IN;
  assign n8933 = ~P1_IR_REG_18__SCAN_IN;
  assign n9842 = ~P1_IR_REG_17__SCAN_IN;
  assign n9268 = ~P1_IR_REG_19__SCAN_IN;
  assign n8934 = ~n9268 | ~n9266;
  assign n8958 = ~P1_IR_REG_21__SCAN_IN;
  assign n8935 = ~P1_IR_REG_22__SCAN_IN;
  assign n8944 = ~P1_IR_REG_23__SCAN_IN;
  assign n8936 = ~P1_IR_REG_24__SCAN_IN;
  assign n8938 = ~n7400 | ~P1_IR_REG_31__SCAN_IN;
  assign n8940 = ~n8938 | ~P1_IR_REG_25__SCAN_IN;
  assign n8949 = ~P1_IR_REG_25__SCAN_IN;
  assign n8939 = ~n8949 | ~P1_IR_REG_31__SCAN_IN;
  assign n8941 = ~n8940 | ~n8939;
  assign n13338 = ~n8941 | ~n8988;
  assign n8943 = ~n13207 & ~n13338;
  assign n8942 = ~n8988 | ~P1_IR_REG_31__SCAN_IN;
  assign n8946 = n8945 | n8944;
  assign n10960 = ~n8947 | ~n8946;
  assign P1_U3086 = ~P1_STATE_REG_SCAN_IN;
  assign n8948 = ~P1_IR_REG_26__SCAN_IN;
  assign n8950 = n8949 & n8948;
  assign n8993 = ~P1_IR_REG_27__SCAN_IN;
  assign n8989 = ~P1_IR_REG_28__SCAN_IN;
  assign n8954 = n8952 | n8993;
  assign n8955 = ~n8961 | ~P1_IR_REG_31__SCAN_IN;
  assign n12950 = ~n8955 ^ n8935;
  assign n8957 = n8956 | n9681;
  assign n8960 = ~n8957 | ~P1_IR_REG_21__SCAN_IN;
  assign n8959 = ~n8958 | ~P1_IR_REG_31__SCAN_IN;
  assign n8962 = ~n8960 | ~n8959;
  assign n12800 = ~n8962 | ~n8961;
  assign n11253 = n12950 | n12800;
  assign n8990 = ~n7398 | ~n8993;
  assign n8992 = ~P1_IR_REG_29__SCAN_IN;
  assign n11189 = ~n7398 | ~n7900;
  assign n11187 = ~P1_IR_REG_30__SCAN_IN;
  assign n9056 = P1_REG3_REG_4__SCAN_IN & P1_REG3_REG_3__SCAN_IN;
  assign n9059 = ~n9056 | ~P1_REG3_REG_5__SCAN_IN;
  assign n11492 = ~P1_REG3_REG_6__SCAN_IN;
  assign n9576 = ~n9059 & ~n11492;
  assign n12902 = ~n9576 ^ P1_REG3_REG_7__SCAN_IN;
  assign n8995 = ~n12902;
  assign n8998 = ~n7327 | ~n8995;
  assign n9072 = n9377 & n8996;
  assign n8997 = ~n10480 | ~P1_REG1_REG_7__SCAN_IN;
  assign n9004 = ~n8998 | ~n8997;
  assign n9002 = ~n9049 | ~P1_REG0_REG_7__SCAN_IN;
  assign n8999 = ~n9377;
  assign n9580 = ~n9078;
  assign n9000 = ~P1_REG2_REG_7__SCAN_IN;
  assign n9001 = n9606 | n9000;
  assign n9003 = ~n9002 | ~n9001;
  assign n9008 = ~n9071 | ~P1_REG3_REG_0__SCAN_IN;
  assign n9007 = ~n9072 | ~P1_REG1_REG_0__SCAN_IN;
  assign n9013 = ~n9008 | ~n9007;
  assign n9011 = ~n9049 | ~P1_REG0_REG_0__SCAN_IN;
  assign n9009 = ~P1_REG2_REG_0__SCAN_IN;
  assign n9010 = n9078 | n9009;
  assign n9012 = ~n9011 | ~n9010;
  assign n12534 = ~n9059 ^ n11492;
  assign n9016 = ~n12534;
  assign n9018 = ~n7327 | ~n9016;
  assign n9017 = ~n10480 | ~P1_REG1_REG_6__SCAN_IN;
  assign n9023 = ~n9018 | ~n9017;
  assign n9021 = ~n9049 | ~P1_REG0_REG_6__SCAN_IN;
  assign n9019 = ~P1_REG2_REG_6__SCAN_IN;
  assign n9020 = n9606 | n9019;
  assign n9022 = ~n9021 | ~n9020;
  assign n9027 = ~P1_REG3_REG_3__SCAN_IN;
  assign n9029 = ~n7327 | ~n9027;
  assign n9028 = ~n10480 | ~P1_REG1_REG_3__SCAN_IN;
  assign n9034 = ~n9029 | ~n9028;
  assign n9032 = ~n9049 | ~P1_REG0_REG_3__SCAN_IN;
  assign n9030 = ~P1_REG2_REG_3__SCAN_IN;
  assign n9031 = n9078 | n9030;
  assign n9033 = ~n9032 | ~n9031;
  assign n12181 = P1_REG3_REG_4__SCAN_IN ^ P1_REG3_REG_3__SCAN_IN;
  assign n9038 = ~n7327 | ~n12181;
  assign n9037 = ~n10480 | ~P1_REG1_REG_4__SCAN_IN;
  assign n9043 = ~n9038 | ~n9037;
  assign n9041 = ~n9049 | ~P1_REG0_REG_4__SCAN_IN;
  assign n9039 = ~P1_REG2_REG_4__SCAN_IN;
  assign n9040 = n9606 | n9039;
  assign n9042 = ~n9041 | ~n9040;
  assign n10454 = ~n9043 & ~n9042;
  assign n9048 = ~n9071 | ~P1_REG3_REG_2__SCAN_IN;
  assign n9046 = ~P1_REG2_REG_2__SCAN_IN;
  assign n9047 = n9078 | n9046;
  assign n9053 = ~n9048 | ~n9047;
  assign n9051 = ~n9072 | ~P1_REG1_REG_2__SCAN_IN;
  assign n9050 = ~n9049 | ~P1_REG0_REG_2__SCAN_IN;
  assign n9052 = ~n9051 | ~n9050;
  assign n9058 = ~n9056;
  assign n9057 = ~P1_REG3_REG_5__SCAN_IN;
  assign n9060 = ~n9058 | ~n9057;
  assign n12776 = ~n9060 | ~n9059;
  assign n9061 = ~n12776;
  assign n9063 = ~n7327 | ~n9061;
  assign n9062 = ~n10480 | ~P1_REG1_REG_5__SCAN_IN;
  assign n9068 = ~n9063 | ~n9062;
  assign n9066 = ~n9049 | ~P1_REG0_REG_5__SCAN_IN;
  assign n9064 = ~P1_REG2_REG_5__SCAN_IN;
  assign n9065 = n9606 | n9064;
  assign n9067 = ~n9066 | ~n9065;
  assign n9074 = ~n9071 | ~P1_REG3_REG_1__SCAN_IN;
  assign n9073 = ~n9072 | ~P1_REG1_REG_1__SCAN_IN;
  assign n9082 = ~n9074 | ~n9073;
  assign n9075 = ~P1_REG0_REG_1__SCAN_IN;
  assign n9080 = n9076 | n9075;
  assign n9077 = ~P1_REG2_REG_1__SCAN_IN;
  assign n9079 = n9078 | n9077;
  assign n9081 = ~n9080 | ~n9079;
  assign n11249 = n10960 & P1_STATE_REG_SCAN_IN;
  assign n9271 = ~n9269 | ~n9268;
  assign n9267 = ~n9271 | ~P1_IR_REG_31__SCAN_IN;
  assign n9270 = n9269 | n9268;
  assign n14881 = ~n9271 | ~n9270;
  assign n9362 = ~n12567 | ~n14881;
  assign n9273 = ~n10591;
  assign n9278 = ~n9273 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n9276 = ~n9593 | ~n11301;
  assign n9274 = ~P1_IR_REG_31__SCAN_IN | ~P1_IR_REG_0__SCAN_IN;
  assign n11682 = ~n9274 ^ P1_IR_REG_1__SCAN_IN;
  assign n11687 = ~n11682;
  assign n12091 = ~n9278 | ~n9277;
  assign n9279 = ~n11857;
  assign n9291 = ~P1_IR_REG_0__SCAN_IN;
  assign n9286 = ~n9285 | ~SI_0_;
  assign n11022 = ~n9286 ^ P2_DATAO_REG_0__SCAN_IN;
  assign n12085 = ~n9288 | ~n9287;
  assign n10958 = ~n9362;
  assign n9309 = ~n9593 | ~n11289;
  assign n9324 = n9681 | n9307;
  assign n11632 = ~n9324 ^ P1_IR_REG_2__SCAN_IN;
  assign n11296 = ~n11632;
  assign n9310 = ~P2_DATAO_REG_2__SCAN_IN;
  assign n9322 = ~P2_DATAO_REG_3__SCAN_IN;
  assign n9328 = n10591 | n9322;
  assign n9323 = ~P1_IR_REG_2__SCAN_IN;
  assign n9325 = ~n9324 | ~n9323;
  assign n9326 = ~n9325 | ~P1_IR_REG_31__SCAN_IN;
  assign n11483 = ~n9326 ^ P1_IR_REG_3__SCAN_IN;
  assign n11455 = ~n11483;
  assign n9330 = n9328 & n9327;
  assign n9710 = ~n9593;
  assign n9893 = ~n9710;
  assign n9329 = ~n9893 | ~n11316;
  assign n12015 = ~n9330 | ~n9329;
  assign n9342 = ~P2_DATAO_REG_4__SCAN_IN;
  assign n9346 = n10591 | n9342;
  assign n9344 = ~n9343 | ~P1_IR_REG_31__SCAN_IN;
  assign n11600 = ~n9344 ^ P1_IR_REG_4__SCAN_IN;
  assign n11454 = ~n11600;
  assign n9348 = n9346 & n9345;
  assign n9347 = ~n9893 | ~n11321;
  assign n12201 = ~n9348 | ~n9347;
  assign n10956 = ~n12567;
  assign n10962 = n11253 | n9362;
  assign n9513 = ~P2_DATAO_REG_5__SCAN_IN;
  assign n9520 = n10591 | n9513;
  assign n9681 = ~P1_IR_REG_31__SCAN_IN;
  assign n9517 = ~n9514 | ~P1_IR_REG_5__SCAN_IN;
  assign n9516 = ~n9515 | ~P1_IR_REG_31__SCAN_IN;
  assign n9518 = ~n9517 | ~n9516;
  assign n11453 = ~n9518 | ~n9534;
  assign n9522 = n9520 & n9519;
  assign n9521 = ~n9893 | ~n11025;
  assign n9533 = ~P2_DATAO_REG_6__SCAN_IN;
  assign n9536 = n10591 | n9533;
  assign n9550 = ~n9534 | ~P1_IR_REG_31__SCAN_IN;
  assign n11452 = ~n9550 ^ P1_IR_REG_6__SCAN_IN;
  assign n11493 = ~n11452;
  assign n9538 = n9536 & n9535;
  assign n9537 = ~n9893 | ~n11274;
  assign n9548 = ~P2_DATAO_REG_7__SCAN_IN;
  assign n9554 = n10591 | n9548;
  assign n9549 = ~P1_IR_REG_6__SCAN_IN;
  assign n9551 = ~n9550 | ~n9549;
  assign n9569 = n9551 & P1_IR_REG_31__SCAN_IN;
  assign n9552 = ~P1_IR_REG_7__SCAN_IN;
  assign n11713 = ~n9569 ^ n9552;
  assign n11451 = ~n11713;
  assign n9556 = n9554 & n9553;
  assign n9555 = ~n9893 | ~n11306;
  assign n12762 = ~n9556 | ~n9555;
  assign n9575 = ~n9567 | ~n9893;
  assign n9568 = ~P2_DATAO_REG_8__SCAN_IN;
  assign n9573 = n10591 | n9568;
  assign n9570 = ~P1_IR_REG_7__SCAN_IN & ~n9569;
  assign n9571 = ~n9570 & ~n9681;
  assign n11525 = ~P1_IR_REG_8__SCAN_IN ^ n9571;
  assign n9574 = n9573 & n9572;
  assign n9601 = ~n9576 | ~P1_REG3_REG_7__SCAN_IN;
  assign n12945 = P1_REG3_REG_8__SCAN_IN ^ n9601;
  assign n9577 = ~n12945;
  assign n9579 = ~n7327 | ~n9577;
  assign n9578 = ~n10480 | ~P1_REG1_REG_8__SCAN_IN;
  assign n9585 = ~n9579 | ~n9578;
  assign n9583 = ~n9049 | ~P1_REG0_REG_8__SCAN_IN;
  assign n9581 = ~P1_REG2_REG_8__SCAN_IN;
  assign n9582 = n9606 | n9581;
  assign n9584 = ~n9583 | ~n9582;
  assign n9600 = ~n9594 | ~n9893;
  assign n9595 = ~P2_DATAO_REG_9__SCAN_IN;
  assign n9598 = n10591 | n9595;
  assign n9596 = ~n9624 | ~P1_IR_REG_31__SCAN_IN;
  assign n11552 = ~n9596 ^ P1_IR_REG_9__SCAN_IN;
  assign n11449 = ~n11552;
  assign n9599 = n9598 & n9597;
  assign n11524 = ~P1_REG3_REG_8__SCAN_IN;
  assign n9632 = ~n9601 & ~n11524;
  assign n12979 = ~P1_REG3_REG_9__SCAN_IN ^ n9632;
  assign n9602 = ~n12979;
  assign n9604 = ~n7327 | ~n9602;
  assign n9603 = ~n10480 | ~P1_REG1_REG_9__SCAN_IN;
  assign n9610 = ~n9604 | ~n9603;
  assign n9608 = ~n9049 | ~P1_REG0_REG_9__SCAN_IN;
  assign n9605 = ~P1_REG2_REG_9__SCAN_IN;
  assign n9607 = n9606 | n9605;
  assign n9609 = ~n9608 | ~n9607;
  assign n9631 = ~n9622 | ~n9893;
  assign n9623 = ~P2_DATAO_REG_10__SCAN_IN;
  assign n9629 = n10591 | n9623;
  assign n9625 = n9624 | P1_IR_REG_9__SCAN_IN;
  assign n9683 = ~n9625 | ~P1_IR_REG_31__SCAN_IN;
  assign n9626 = ~P1_IR_REG_10__SCAN_IN;
  assign n9653 = n9683 & n9626;
  assign n9627 = ~n9683 & ~n9626;
  assign n11731 = ~n9653 & ~n9627;
  assign n11551 = ~n11731;
  assign n9630 = n9629 & n9628;
  assign n9659 = n9632 & P1_REG3_REG_9__SCAN_IN;
  assign n13326 = ~P1_REG3_REG_10__SCAN_IN ^ n9659;
  assign n9633 = ~n13326;
  assign n9635 = ~n7327 | ~n9633;
  assign n9634 = ~n9072 | ~P1_REG1_REG_10__SCAN_IN;
  assign n9640 = ~n9635 | ~n9634;
  assign n9638 = ~n9049 | ~P1_REG0_REG_10__SCAN_IN;
  assign n9636 = ~P1_REG2_REG_10__SCAN_IN;
  assign n9637 = n9606 | n9636;
  assign n9639 = ~n9638 | ~n9637;
  assign n9658 = ~n9651 | ~n9893;
  assign n9652 = ~P2_DATAO_REG_11__SCAN_IN;
  assign n9656 = n10591 | n9652;
  assign n9654 = ~n9653 & ~n9681;
  assign n11730 = ~P1_IR_REG_11__SCAN_IN ^ n9654;
  assign n9657 = n9656 & n9655;
  assign n9690 = n9659 & P1_REG3_REG_10__SCAN_IN;
  assign n13510 = ~P1_REG3_REG_11__SCAN_IN ^ n9690;
  assign n9660 = ~n13510;
  assign n9662 = ~n7327 | ~n9660;
  assign n9661 = ~n9072 | ~P1_REG1_REG_11__SCAN_IN;
  assign n9667 = ~n9662 | ~n9661;
  assign n9665 = ~n9049 | ~P1_REG0_REG_11__SCAN_IN;
  assign n9663 = ~P1_REG2_REG_11__SCAN_IN;
  assign n9664 = n9606 | n9663;
  assign n9666 = ~n9665 | ~n9664;
  assign n9689 = ~n9678 | ~n9893;
  assign n9679 = ~P2_DATAO_REG_12__SCAN_IN;
  assign n9687 = n10591 | n9679;
  assign n9682 = n9681 | n9680;
  assign n9684 = ~n9683 | ~n9682;
  assign n9713 = ~n9684 & ~P1_IR_REG_12__SCAN_IN;
  assign n9685 = n9684 & P1_IR_REG_12__SCAN_IN;
  assign n12275 = ~n9713 & ~n9685;
  assign n11816 = ~n12275;
  assign n9688 = n9687 & n9686;
  assign n9719 = n9690 & P1_REG3_REG_11__SCAN_IN;
  assign n13124 = ~P1_REG3_REG_12__SCAN_IN ^ n9719;
  assign n9691 = ~n13124;
  assign n9693 = ~n7327 | ~n9691;
  assign n9692 = ~n9072 | ~P1_REG1_REG_12__SCAN_IN;
  assign n9698 = ~n9693 | ~n9692;
  assign n9696 = ~n9049 | ~P1_REG0_REG_12__SCAN_IN;
  assign n9694 = ~P1_REG2_REG_12__SCAN_IN;
  assign n9695 = n9606 | n9694;
  assign n9697 = ~n9696 | ~n9695;
  assign n9718 = ~n9711 | ~n9893;
  assign n9712 = ~P2_DATAO_REG_13__SCAN_IN;
  assign n9716 = n10591 | n9712;
  assign n9714 = ~n9713 & ~n9681;
  assign n12274 = ~P1_IR_REG_13__SCAN_IN ^ n9714;
  assign n9717 = n9716 & n9715;
  assign n9748 = n9719 & P1_REG3_REG_12__SCAN_IN;
  assign n13518 = ~P1_REG3_REG_13__SCAN_IN ^ n9748;
  assign n9720 = ~n13518;
  assign n9723 = ~n7327 | ~n9720;
  assign n9722 = ~n9072 | ~P1_REG1_REG_13__SCAN_IN;
  assign n9728 = ~n9723 | ~n9722;
  assign n9726 = ~n9049 | ~P1_REG0_REG_13__SCAN_IN;
  assign n9724 = ~P1_REG2_REG_13__SCAN_IN;
  assign n9725 = n9606 | n9724;
  assign n9727 = ~n9726 | ~n9725;
  assign n9747 = ~n9738 | ~n9893;
  assign n9739 = ~P2_DATAO_REG_14__SCAN_IN;
  assign n9745 = n10591 | n9739;
  assign n9740 = ~P1_IR_REG_31__SCAN_IN & ~P1_IR_REG_14__SCAN_IN;
  assign n9765 = n7445 | n9740;
  assign n9741 = P1_IR_REG_31__SCAN_IN & P1_IR_REG_14__SCAN_IN;
  assign n9743 = n9742 & n9741;
  assign n13490 = ~n9765 & ~n9743;
  assign n12641 = ~n13490;
  assign n9746 = n9745 & n9744;
  assign n9776 = n9748 & P1_REG3_REG_13__SCAN_IN;
  assign n13543 = ~P1_REG3_REG_14__SCAN_IN ^ n9776;
  assign n9749 = ~n13543;
  assign n9751 = ~n7327 | ~n9749;
  assign n9750 = ~n9072 | ~P1_REG1_REG_14__SCAN_IN;
  assign n9756 = ~n9751 | ~n9750;
  assign n9754 = ~n9049 | ~P1_REG0_REG_14__SCAN_IN;
  assign n9752 = ~P1_REG2_REG_14__SCAN_IN;
  assign n9753 = n9606 | n9752;
  assign n9755 = ~n9754 | ~n9753;
  assign n9770 = ~n9763 | ~n9893;
  assign n9764 = ~P2_DATAO_REG_15__SCAN_IN;
  assign n9768 = n10591 | n9764;
  assign n9766 = ~n9765 & ~n9681;
  assign n13495 = ~P1_IR_REG_15__SCAN_IN ^ n9766;
  assign n9769 = n9768 & n9767;
  assign n9773 = ~n9049 | ~P1_REG0_REG_15__SCAN_IN;
  assign n9771 = ~P1_REG2_REG_15__SCAN_IN;
  assign n9772 = n9606 | n9771;
  assign n9775 = ~n9773 | ~n9772;
  assign n9774 = n10480 & P1_REG1_REG_15__SCAN_IN;
  assign n9779 = ~n9775 & ~n9774;
  assign n9803 = n9776 & P1_REG3_REG_14__SCAN_IN;
  assign n14053 = ~P1_REG3_REG_15__SCAN_IN ^ n9803;
  assign n9777 = ~n14053;
  assign n9778 = ~n7327 | ~n9777;
  assign n13680 = ~n9779 | ~n9778;
  assign n9797 = ~n9789 | ~n9893;
  assign n9790 = ~P2_DATAO_REG_16__SCAN_IN;
  assign n9795 = n10591 | n9790;
  assign n9791 = ~P1_IR_REG_15__SCAN_IN;
  assign n9792 = ~n7445 | ~n9791;
  assign n9793 = ~n9792 | ~P1_IR_REG_31__SCAN_IN;
  assign n14335 = ~n9793 ^ P1_IR_REG_16__SCAN_IN;
  assign n13793 = ~n14335;
  assign n9796 = n9795 & n9794;
  assign n9800 = ~n9049 | ~P1_REG0_REG_16__SCAN_IN;
  assign n9798 = ~P1_REG2_REG_16__SCAN_IN;
  assign n9799 = n9606 | n9798;
  assign n9802 = ~n9800 | ~n9799;
  assign n9801 = n10480 & P1_REG1_REG_16__SCAN_IN;
  assign n9806 = ~n9802 & ~n9801;
  assign n9828 = n9803 & P1_REG3_REG_15__SCAN_IN;
  assign n14068 = ~P1_REG3_REG_16__SCAN_IN ^ n9828;
  assign n9804 = ~n14068;
  assign n9805 = ~n7327 | ~n9804;
  assign n13879 = ~n9806 | ~n9805;
  assign n9822 = ~n9816 | ~n9893;
  assign n9817 = ~P2_DATAO_REG_17__SCAN_IN;
  assign n9820 = n10591 | n9817;
  assign n9843 = ~n9818 | ~P1_IR_REG_31__SCAN_IN;
  assign n14628 = ~n9843 ^ P1_IR_REG_17__SCAN_IN;
  assign n14334 = ~n14628;
  assign n9821 = n9820 & n9819;
  assign n9825 = ~n9049 | ~P1_REG0_REG_17__SCAN_IN;
  assign n9823 = ~P1_REG2_REG_17__SCAN_IN;
  assign n9824 = n9606 | n9823;
  assign n9827 = ~n9825 | ~n9824;
  assign n9826 = n10480 & P1_REG1_REG_17__SCAN_IN;
  assign n9831 = ~n9827 & ~n9826;
  assign n9850 = n9828 & P1_REG3_REG_16__SCAN_IN;
  assign n14007 = ~P1_REG3_REG_17__SCAN_IN ^ n9850;
  assign n9829 = ~n14007;
  assign n9830 = ~n9829 | ~n7327;
  assign n13679 = ~n9831 | ~n9830;
  assign n9849 = ~n9840 | ~n9893;
  assign n9841 = ~P2_DATAO_REG_18__SCAN_IN;
  assign n9847 = n10591 | n9841;
  assign n9844 = n9843 & n9842;
  assign n9845 = ~n9844 & ~n9681;
  assign n14627 = ~P1_IR_REG_18__SCAN_IN ^ n9845;
  assign n9848 = n9847 & n9846;
  assign n9873 = n9850 & P1_REG3_REG_17__SCAN_IN;
  assign n13763 = ~P1_REG3_REG_18__SCAN_IN ^ n9873;
  assign n9851 = ~n13763;
  assign n9858 = ~n9851 | ~n7327;
  assign n9854 = ~n9049 | ~P1_REG0_REG_18__SCAN_IN;
  assign n9852 = ~P1_REG2_REG_18__SCAN_IN;
  assign n9853 = n9606 | n9852;
  assign n9856 = ~n9854 | ~n9853;
  assign n9855 = n9072 & P1_REG1_REG_18__SCAN_IN;
  assign n9857 = ~n9856 & ~n9855;
  assign n14120 = ~n9858 | ~n9857;
  assign n9872 = ~n9867 | ~n9893;
  assign n9868 = ~P2_DATAO_REG_19__SCAN_IN;
  assign n9870 = n10591 | n9868;
  assign n9871 = n9870 & n9869;
  assign n9896 = n9873 & P1_REG3_REG_18__SCAN_IN;
  assign n14312 = ~P1_REG3_REG_19__SCAN_IN ^ n9896;
  assign n9874 = ~n14312;
  assign n9881 = ~n9874 | ~n7327;
  assign n9877 = ~n9049 | ~P1_REG0_REG_19__SCAN_IN;
  assign n9875 = ~P1_REG2_REG_19__SCAN_IN;
  assign n9876 = n9606 | n9875;
  assign n9879 = ~n9877 | ~n9876;
  assign n9878 = n9072 & P1_REG1_REG_19__SCAN_IN;
  assign n9880 = ~n9879 & ~n9878;
  assign n14106 = ~n9881 | ~n9880;
  assign n9895 = ~n12727 | ~n9893;
  assign n12568 = ~P2_DATAO_REG_20__SCAN_IN;
  assign n9894 = n10591 | n12568;
  assign n9912 = n9896 & P1_REG3_REG_19__SCAN_IN;
  assign n14475 = ~P1_REG3_REG_20__SCAN_IN ^ n9912;
  assign n9897 = ~n14475;
  assign n9904 = ~n9897 | ~n7327;
  assign n9900 = ~n9049 | ~P1_REG0_REG_20__SCAN_IN;
  assign n9898 = ~P1_REG2_REG_20__SCAN_IN;
  assign n9899 = n9606 | n9898;
  assign n9902 = ~n9900 | ~n9899;
  assign n9901 = n9072 & P1_REG1_REG_20__SCAN_IN;
  assign n9903 = ~n9902 & ~n9901;
  assign n14141 = ~n9904 | ~n9903;
  assign n9911 = ~n12849 | ~n9893;
  assign n12801 = ~P2_DATAO_REG_21__SCAN_IN;
  assign n9910 = n10591 | n12801;
  assign n9934 = n9912 & P1_REG3_REG_20__SCAN_IN;
  assign n14600 = ~P1_REG3_REG_21__SCAN_IN ^ n9934;
  assign n9913 = ~n14600;
  assign n9920 = ~n9913 | ~n7327;
  assign n9916 = ~n9049 | ~P1_REG0_REG_21__SCAN_IN;
  assign n9914 = ~P1_REG2_REG_21__SCAN_IN;
  assign n9915 = n9606 | n9914;
  assign n9918 = ~n9916 | ~n9915;
  assign n9917 = n9072 & P1_REG1_REG_21__SCAN_IN;
  assign n9919 = ~n9918 & ~n9917;
  assign n14105 = ~n9920 | ~n9919;
  assign n9933 = ~n13040 | ~n9893;
  assign n12951 = ~P2_DATAO_REG_22__SCAN_IN;
  assign n9932 = n10591 | n12951;
  assign n9952 = n9934 & P1_REG3_REG_21__SCAN_IN;
  assign n14285 = ~P1_REG3_REG_22__SCAN_IN ^ n9952;
  assign n9949 = ~n14285;
  assign n9941 = ~n9949 | ~n7327;
  assign n9937 = ~n9049 | ~P1_REG0_REG_22__SCAN_IN;
  assign n9935 = ~P1_REG2_REG_22__SCAN_IN;
  assign n9936 = n9606 | n9935;
  assign n9939 = ~n9937 | ~n9936;
  assign n9938 = n9072 & P1_REG1_REG_22__SCAN_IN;
  assign n9940 = ~n9939 & ~n9938;
  assign n14139 = ~n9941 | ~n9940;
  assign n10551 = ~n14139;
  assign n10017 = n9952 & P1_REG3_REG_22__SCAN_IN;
  assign n14421 = ~P1_REG3_REG_23__SCAN_IN ^ n10017;
  assign n10159 = ~n14421;
  assign n9959 = ~n10159 | ~n7327;
  assign n9955 = ~n9049 | ~P1_REG0_REG_23__SCAN_IN;
  assign n9953 = ~P1_REG2_REG_23__SCAN_IN;
  assign n9954 = n9606 | n9953;
  assign n9957 = ~n9955 | ~n9954;
  assign n9956 = n9072 & P1_REG1_REG_23__SCAN_IN;
  assign n9958 = ~n9957 & ~n9956;
  assign n11756 = ~n9959 | ~n9958;
  assign n10006 = ~n13171 | ~n9893;
  assign n13168 = ~P2_DATAO_REG_23__SCAN_IN;
  assign n10005 = n10591 | n13168;
  assign n10016 = ~n13335 | ~n9893;
  assign n13208 = ~P2_DATAO_REG_24__SCAN_IN;
  assign n10015 = n10591 | n13208;
  assign n10037 = n10017 & P1_REG3_REG_23__SCAN_IN;
  assign n14721 = ~P1_REG3_REG_24__SCAN_IN ^ n10037;
  assign n10047 = ~n14721;
  assign n10024 = ~n10047 | ~n7327;
  assign n10020 = ~n9049 | ~P1_REG0_REG_24__SCAN_IN;
  assign n10018 = ~P1_REG2_REG_24__SCAN_IN;
  assign n10019 = n9606 | n10018;
  assign n10022 = ~n10020 | ~n10019;
  assign n10021 = n9072 & P1_REG1_REG_24__SCAN_IN;
  assign n10023 = ~n10022 & ~n10021;
  assign n11926 = ~n10024 | ~n10023;
  assign n10468 = ~n14723;
  assign n10219 = n10037 & P1_REG3_REG_24__SCAN_IN;
  assign n14748 = ~P1_REG3_REG_25__SCAN_IN ^ n10219;
  assign n10229 = ~n14748;
  assign n10044 = ~n10229 | ~n7327;
  assign n10040 = ~n9049 | ~P1_REG0_REG_25__SCAN_IN;
  assign n10038 = ~P1_REG2_REG_25__SCAN_IN;
  assign n10039 = n9606 | n10038;
  assign n10042 = ~n10040 | ~n10039;
  assign n10041 = n9072 & P1_REG1_REG_25__SCAN_IN;
  assign n10043 = ~n10042 & ~n10041;
  assign n12065 = ~n10044 | ~n10043;
  assign n10204 = ~n13457 | ~n9893;
  assign n10202 = ~P2_DATAO_REG_25__SCAN_IN;
  assign n10203 = n10591 | n10202;
  assign n10325 = ~n10219 | ~P1_REG3_REG_25__SCAN_IN;
  assign n14842 = P1_REG3_REG_26__SCAN_IN ^ n10325;
  assign n10336 = ~n14842;
  assign n10226 = ~n10336 | ~n7327;
  assign n10222 = ~n9049 | ~P1_REG0_REG_26__SCAN_IN;
  assign n10220 = ~P1_REG2_REG_26__SCAN_IN;
  assign n10221 = n9606 | n10220;
  assign n10224 = ~n10222 | ~n10221;
  assign n10223 = n9072 & P1_REG1_REG_26__SCAN_IN;
  assign n10225 = ~n10224 & ~n10223;
  assign n12211 = ~n10226 | ~n10225;
  assign n10312 = ~n13464 | ~n9893;
  assign n13461 = ~P2_DATAO_REG_26__SCAN_IN;
  assign n10311 = n10591 | n13461;
  assign n10441 = ~n12211;
  assign n10324 = ~P1_REG3_REG_26__SCAN_IN;
  assign n10428 = ~n10325 & ~n10324;
  assign n15026 = ~P1_REG3_REG_27__SCAN_IN ^ n10428;
  assign n10326 = ~n15026;
  assign n10333 = ~n10326 | ~n7327;
  assign n10329 = ~n9049 | ~P1_REG0_REG_27__SCAN_IN;
  assign n10327 = ~P1_REG2_REG_27__SCAN_IN;
  assign n10328 = n9606 | n10327;
  assign n10331 = ~n10329 | ~n10328;
  assign n10330 = n10480 & P1_REG1_REG_27__SCAN_IN;
  assign n10332 = ~n10331 & ~n10330;
  assign n12332 = ~n10333 | ~n10332;
  assign n13834 = ~P2_DATAO_REG_28__SCAN_IN;
  assign n10427 = n10591 | n13834;
  assign n10475 = n10428 & P1_REG3_REG_27__SCAN_IN;
  assign n15104 = ~P1_REG3_REG_28__SCAN_IN ^ n10475;
  assign n10429 = ~n15104;
  assign n10436 = ~n10429 | ~n7327;
  assign n10432 = ~n9049 | ~P1_REG0_REG_28__SCAN_IN;
  assign n10430 = ~P1_REG2_REG_28__SCAN_IN;
  assign n10431 = n9606 | n10430;
  assign n10434 = ~n10432 | ~n10431;
  assign n10433 = n10480 & P1_REG1_REG_28__SCAN_IN;
  assign n10435 = ~n10434 & ~n10433;
  assign n12423 = ~n10436 | ~n10435;
  assign n10437 = ~n10738;
  assign n10997 = ~n12423;
  assign n10945 = n15134 & n10997;
  assign n10440 = ~n13658 | ~n9593;
  assign n10438 = ~P2_DATAO_REG_27__SCAN_IN;
  assign n10439 = n10591 | n10438;
  assign n10737 = ~n15031 | ~n12332;
  assign n10967 = ~n12332;
  assign n10736 = ~n15090 | ~n10967;
  assign n10793 = ~n10736 | ~n10737;
  assign n10884 = ~n14856 | ~n12211;
  assign n10735 = ~n14867 | ~n10441;
  assign n14847 = ~n10884 | ~n10735;
  assign n10442 = ~n11926;
  assign n10817 = n14723 & n10442;
  assign n10816 = ~n14543 & ~n11756;
  assign n10814 = ~n10552 | ~n14139;
  assign n10722 = ~n14397 | ~n10551;
  assign n10810 = ~n14610 | ~n14105;
  assign n10443 = ~n14105;
  assign n10723 = ~n10549 | ~n10443;
  assign n14485 = ~n14227;
  assign n10703 = ~n14485 | ~n14141;
  assign n10444 = ~n14106;
  assign n10702 = n14162 | n10444;
  assign n10885 = ~n14162 | ~n10444;
  assign n10783 = ~n10702 | ~n10885;
  assign n10605 = ~n13767 | ~n14120;
  assign n10464 = ~n14013 | ~n13679;
  assign n10926 = ~n10605 | ~n10464;
  assign n10857 = ~n10926 | ~n10696;
  assign n10462 = ~n13879;
  assign n10609 = n13592 & n13561;
  assign n10460 = ~n11476;
  assign n10608 = ~n13250 & ~n10460;
  assign n10445 = ~n10618;
  assign n10848 = n13128 | n13231;
  assign n13134 = ~n10445 | ~n10848;
  assign n10844 = n13502 | n12957;
  assign n10664 = n13320 & n13186;
  assign n10828 = n12921 | n12956;
  assign n10662 = ~n12921 | ~n12956;
  assign n10514 = ~n12808;
  assign n10827 = ~n12942 | ~n10514;
  assign n12349 = ~n10507 | ~n12460;
  assign n10832 = ~n10454 | ~n12201;
  assign n10833 = n10507 | n12460;
  assign n10835 = ~n12470 | ~n12531;
  assign n10892 = n11935 | n10451;
  assign n10633 = ~n10451 | ~n11935;
  assign n11883 = n10892 & n10633;
  assign n11869 = ~n12085;
  assign n12081 = ~n11915 & ~n11869;
  assign n12103 = ~n12091;
  assign n10886 = ~n9279 | ~n12103;
  assign n10623 = ~n12081 | ~n10886;
  assign n10630 = ~n11857 | ~n12091;
  assign n11881 = ~n10623 | ~n10630;
  assign n10452 = ~n11883 | ~n11881;
  assign n11989 = ~n10452 | ~n10633;
  assign n10635 = n10503 | n12015;
  assign n10634 = ~n10503 | ~n12015;
  assign n11991 = ~n10635 | ~n10634;
  assign n11988 = ~n11991;
  assign n10453 = ~n11989 | ~n11988;
  assign n12344 = ~n10453 | ~n10634;
  assign n12345 = n10454 | n12201;
  assign n10455 = n10646 & n12345;
  assign n10839 = ~n12344 | ~n10455;
  assign n12908 = ~n12762;
  assign n10650 = ~n12908 | ~n10511;
  assign n12656 = ~n10511;
  assign n10906 = ~n12656 | ~n12762;
  assign n12476 = ~n10650 | ~n10906;
  assign n10515 = ~n12942;
  assign n10651 = ~n10515 | ~n12808;
  assign n10658 = ~n10664;
  assign n10518 = ~n13186;
  assign n10831 = ~n13004 | ~n10518;
  assign n12966 = ~n10658 | ~n10831;
  assign n10458 = ~n10844;
  assign n10614 = n13502 & n12957;
  assign n13200 = ~n10458 & ~n10614;
  assign n10915 = ~n13250 | ~n10460;
  assign n10461 = ~n10915;
  assign n10681 = ~n10609;
  assign n10607 = ~n13592 & ~n13561;
  assign n10611 = ~n10607;
  assign n13535 = ~n10681 | ~n10611;
  assign n10683 = ~n14060 & ~n13680;
  assign n10690 = ~n14073 & ~n10462;
  assign n10923 = n10690 | n13674;
  assign n10693 = n14013 | n13679;
  assign n10709 = ~n14141;
  assign n10547 = ~n14485 | ~n10709;
  assign n10716 = ~n14227 | ~n14141;
  assign n14109 = ~n10547 | ~n10716;
  assign n10807 = ~n14543 | ~n11756;
  assign n10467 = ~n10807;
  assign n10469 = ~n10817;
  assign n10805 = ~n10468 | ~n11926;
  assign n10604 = ~n10469 | ~n10805;
  assign n10474 = ~n13957 | ~n9893;
  assign n13952 = ~P2_DATAO_REG_29__SCAN_IN;
  assign n10473 = n10591 | n13952;
  assign n15149 = ~n10474 | ~n10473;
  assign n15153 = ~n10475 | ~P1_REG3_REG_28__SCAN_IN;
  assign n10476 = ~n15153;
  assign n10484 = ~n10476 | ~n7327;
  assign n10479 = ~n9049 | ~P1_REG0_REG_29__SCAN_IN;
  assign n10477 = ~P1_REG2_REG_29__SCAN_IN;
  assign n10478 = n9606 | n10477;
  assign n10482 = ~n10479 | ~n10478;
  assign n10481 = n10480 & P1_REG1_REG_29__SCAN_IN;
  assign n10483 = ~n10482 & ~n10481;
  assign n12287 = ~n10484 | ~n10483;
  assign n10485 = ~n12287;
  assign n10741 = n15149 | n10485;
  assign n10949 = ~n15149 | ~n10485;
  assign n10796 = ~n10741 | ~n10949;
  assign n10491 = ~n10480 | ~P1_REG1_REG_30__SCAN_IN;
  assign n10490 = ~n9049 | ~P1_REG0_REG_30__SCAN_IN;
  assign n10494 = ~n10491 | ~n10490;
  assign n10492 = ~P1_REG2_REG_30__SCAN_IN;
  assign n10493 = ~n9606 & ~n10492;
  assign n11365 = ~n10494 & ~n10493;
  assign n12089 = ~n10886 | ~n10630;
  assign n12343 = ~n12345 | ~n10832;
  assign n13559 = ~n13555;
  assign n13676 = ~n10925 & ~n10690;
  assign n10585 = ~n10583 | ~n9593;
  assign n10584 = ~n9273 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n14782 = ~n10585 | ~n10584;
  assign n14793 = ~n14782;
  assign n10587 = ~n9072 | ~P1_REG1_REG_31__SCAN_IN;
  assign n10586 = ~n9049 | ~P1_REG0_REG_31__SCAN_IN;
  assign n10590 = ~n10587 | ~n10586;
  assign n10588 = ~P1_REG2_REG_31__SCAN_IN;
  assign n10589 = ~n9606 & ~n10588;
  assign n11352 = n10590 | n10589;
  assign n14738 = ~n11352;
  assign n10745 = ~n14738 & ~n11365;
  assign n10871 = ~n14793 & ~n10745;
  assign n10593 = ~n14250 | ~n9593;
  assign n11185 = ~P2_DATAO_REG_31__SCAN_IN;
  assign n10592 = n10591 | n11185;
  assign n14837 = ~n10593 | ~n10592;
  assign n10954 = ~n14837 & ~n14738;
  assign n10742 = ~n10871 & ~n10954;
  assign n10947 = ~n10741 | ~n10738;
  assign n10739 = ~n10945;
  assign n10867 = ~n10739 | ~n10736;
  assign n10594 = ~n10805;
  assign n10754 = ~n12950 | ~n14898;
  assign n10595 = n10806 & n10754;
  assign n10596 = n10884 & n10595;
  assign n10600 = ~n10597 | ~n10596;
  assign n10598 = ~n10735;
  assign n10862 = ~n10598 & ~n10937;
  assign n10753 = ~n10754;
  assign n10599 = ~n10862 | ~n10753;
  assign n10732 = ~n10600 | ~n10599;
  assign n10602 = n10816 | n10753;
  assign n10601 = ~n10807 | ~n10753;
  assign n10603 = n10602 & n10601;
  assign n10727 = ~n10604 & ~n10603;
  assign n10855 = n10696 & n10693;
  assign n10606 = ~n10855;
  assign n10931 = ~n10606 | ~n10605;
  assign n10676 = ~n10923;
  assign n10921 = n10683 | n10607;
  assign n10674 = ~n10921;
  assign n10825 = ~n10609 & ~n10608;
  assign n10613 = ~n10825 | ~n10754;
  assign n10610 = n10915 & n10753;
  assign n10612 = ~n10611 | ~n10610;
  assign n10673 = ~n10613 | ~n10612;
  assign n10615 = ~n10848;
  assign n10826 = ~n10618 & ~n10614;
  assign n10616 = n10615 | n10826;
  assign n10620 = ~n10616 | ~n10753;
  assign n10617 = n10848 & n10844;
  assign n10914 = n10618 | n10617;
  assign n10619 = ~n10914 | ~n10754;
  assign n10670 = ~n10620 | ~n10619;
  assign n10621 = n10892 & n10754;
  assign n10622 = ~n10621 | ~n10886;
  assign n10625 = ~n10632 | ~n10623;
  assign n10624 = n10892 & n10635;
  assign n10627 = ~n10625 | ~n10624;
  assign n10626 = n10832 & n10634;
  assign n10629 = ~n10627 | ~n10626;
  assign n10628 = n12345 & n10753;
  assign n10640 = ~n10629 | ~n10628;
  assign n10761 = ~n12081;
  assign n10631 = ~n10761 | ~n10630;
  assign n10895 = n10634 & n10633;
  assign n10898 = n12345 & n10635;
  assign n10638 = ~n10636 | ~n10898;
  assign n10637 = n10832 & n10754;
  assign n10639 = ~n10638 | ~n10637;
  assign n10645 = ~n10640 | ~n10639;
  assign n10642 = ~n10645 | ~n12349;
  assign n10641 = n10833 & n10835;
  assign n10643 = ~n10642 | ~n10641;
  assign n10656 = ~n10644 | ~n10753;
  assign n10647 = ~n10645 | ~n10833;
  assign n10649 = ~n10647 | ~n10646;
  assign n10648 = n10906 & n10835;
  assign n10652 = ~n10649 | ~n10648;
  assign n10840 = n10651 & n10650;
  assign n10654 = ~n10652 | ~n10840;
  assign n10653 = n10827 & n10754;
  assign n10655 = ~n10654 | ~n10653;
  assign n10657 = ~n10656 | ~n10655;
  assign n10665 = ~n10657 | ~n12815;
  assign n10659 = ~n10665 | ~n10828;
  assign n10661 = ~n10659 | ~n10658;
  assign n10660 = n10831 & n10753;
  assign n10669 = ~n10661 | ~n10660;
  assign n10663 = ~n10662;
  assign n10841 = ~n10664 & ~n10663;
  assign n10666 = ~n10665 | ~n10841;
  assign n10667 = ~n10666 | ~n10831;
  assign n10668 = ~n10667 | ~n10754;
  assign n10672 = ~n10671 | ~n13237;
  assign n10682 = ~n10673 | ~n10672;
  assign n10675 = ~n10674 | ~n10682;
  assign n10677 = ~n10676 | ~n10675;
  assign n10688 = ~n10925;
  assign n10678 = n10677 & n10688;
  assign n10679 = n10926 | n10678;
  assign n10680 = n10679 & n10754;
  assign n10700 = ~n10931 | ~n10680;
  assign n10685 = ~n10682 | ~n10681;
  assign n10684 = ~n10683;
  assign n10687 = ~n10685 | ~n10684;
  assign n10686 = ~n13674;
  assign n10689 = ~n10687 | ~n10686;
  assign n10692 = ~n10689 | ~n10688;
  assign n10691 = ~n10690;
  assign n10694 = ~n10692 | ~n10691;
  assign n10695 = n10694 & n10693;
  assign n10697 = n10695 | n10926;
  assign n10698 = ~n10697 | ~n10696;
  assign n10699 = ~n10698 | ~n10753;
  assign n10701 = ~n10700 | ~n10699;
  assign n10708 = ~n10701 | ~n14126;
  assign n10824 = ~n10703 | ~n10702;
  assign n10706 = ~n10824 & ~n10753;
  assign n10704 = ~n10885 | ~n10753;
  assign n10811 = n14227 & n10709;
  assign n10705 = ~n10704 & ~n10811;
  assign n10707 = n10706 | n10705;
  assign n10720 = ~n10708 | ~n10707;
  assign n10710 = ~n10720 | ~n10709;
  assign n10711 = ~n10710 | ~n10723;
  assign n10822 = n10814 & n10810;
  assign n10712 = ~n10711 | ~n10822;
  assign n10714 = ~n10712 | ~n10753;
  assign n10713 = ~n10810 | ~n10754;
  assign n10715 = ~n10714 | ~n10713;
  assign n10717 = ~n10716;
  assign n10719 = ~n10822 | ~n10717;
  assign n10718 = ~n14485 | ~n10754;
  assign n10721 = ~n10719 | ~n10718;
  assign n10812 = n10723 & n10722;
  assign n10724 = n10812 | n10753;
  assign n10725 = ~n10814 & ~n10753;
  assign n10726 = ~n14429 & ~n10725;
  assign n10728 = ~n10817 | ~n10753;
  assign n10730 = ~n10729 | ~n10728;
  assign n10731 = ~n14758 | ~n10730;
  assign n10866 = ~n10737 | ~n10884;
  assign n10733 = ~n10949 | ~n10753;
  assign n10746 = ~n10734 & ~n10733;
  assign n10740 = ~n10949;
  assign n10941 = ~n10736 | ~n10735;
  assign n10942 = ~n10737;
  assign n10760 = ~n14782 & ~n11365;
  assign n10874 = ~n10760 | ~n11352;
  assign n10743 = ~n14782 | ~n10753;
  assign n10752 = ~n10744 | ~n10743;
  assign n10748 = ~n10746 | ~n10745;
  assign n10875 = n14837 & n14738;
  assign n10747 = ~n10875;
  assign n10750 = ~n10748 | ~n10747;
  assign n10749 = ~n10874 & ~n10754;
  assign n10751 = ~n10750 & ~n10749;
  assign n10802 = n10752 & n10751;
  assign n10756 = n10875 | n10753;
  assign n10755 = n10954 | n10754;
  assign n10757 = ~n10756 | ~n10755;
  assign n10758 = ~n10757 | ~n12950;
  assign n10759 = ~n10802 & ~n10758;
  assign n10883 = ~n10760 & ~n10875;
  assign n10786 = ~n10822;
  assign n10888 = ~n11915 | ~n11869;
  assign n11863 = n10761 & n10888;
  assign n10762 = ~n11863 | ~n11883;
  assign n10763 = ~n10762 & ~n12089;
  assign n12449 = ~n12460 ^ n12340;
  assign n10764 = n10763 & n12449;
  assign n10771 = ~n12650 | ~n10764;
  assign n10765 = ~n12476;
  assign n10768 = ~n10765 | ~n12357;
  assign n10766 = ~n12343;
  assign n10767 = ~n10766 | ~n11988;
  assign n10769 = ~n10768 & ~n10767;
  assign n10770 = ~n12815 | ~n10769;
  assign n10772 = ~n10771 & ~n10770;
  assign n10773 = ~n13200 | ~n10772;
  assign n10776 = ~n12966 & ~n10773;
  assign n10775 = ~n13535 & ~n10774;
  assign n10777 = ~n10776 | ~n10775;
  assign n10778 = ~n13134 & ~n10777;
  assign n10780 = ~n13676 | ~n10778;
  assign n10779 = ~n13559 | ~n13876;
  assign n10781 = ~n10780 & ~n10779;
  assign n10782 = ~n10781 | ~n14109;
  assign n10784 = ~n10783 & ~n10782;
  assign n10785 = ~n13775 | ~n10784;
  assign n10787 = ~n10786 & ~n10785;
  assign n10788 = ~n10812 | ~n10787;
  assign n10789 = ~n14429 & ~n10788;
  assign n10790 = ~n14758 | ~n10789;
  assign n10791 = ~n14847 & ~n10790;
  assign n10792 = ~n14676 | ~n10791;
  assign n10794 = ~n10793 & ~n10792;
  assign n10795 = ~n15119 | ~n10794;
  assign n10797 = ~n10796 & ~n10795;
  assign n10798 = ~n10883 | ~n10797;
  assign n10799 = ~n10954 & ~n10798;
  assign n10948 = ~n11365 | ~n14782;
  assign n10800 = ~n10799 | ~n10948;
  assign n10801 = ~n10800 ^ n14898;
  assign n10804 = ~n10802;
  assign n10803 = ~n10875 & ~n14881;
  assign n10882 = ~n10804 | ~n10803;
  assign n10809 = ~n10806 | ~n10805;
  assign n10808 = ~n10817 & ~n10807;
  assign n10821 = ~n10809 & ~n10808;
  assign n10813 = ~n10811 | ~n10810;
  assign n10815 = ~n10813 | ~n10812;
  assign n10819 = ~n10815 | ~n10814;
  assign n10818 = ~n10817 & ~n10816;
  assign n10820 = ~n10819 | ~n10818;
  assign n10934 = ~n10821 | ~n10820;
  assign n10864 = ~n10934;
  assign n10823 = ~n10822 | ~n10821;
  assign n10932 = ~n10824 & ~n10823;
  assign n10919 = ~n10825;
  assign n10912 = ~n10826;
  assign n10829 = ~n10828 | ~n10827;
  assign n10830 = ~n10841 | ~n10829;
  assign n10911 = ~n10831 | ~n10830;
  assign n10834 = ~n10833 | ~n10832;
  assign n10836 = ~n10834 | ~n12349;
  assign n10901 = ~n10836 | ~n10835;
  assign n10837 = ~n10901 | ~n10903;
  assign n10838 = n10837 & n10906;
  assign n10843 = ~n10839 | ~n10838;
  assign n10909 = ~n10841 | ~n10840;
  assign n10842 = ~n10909;
  assign n10845 = ~n10843 | ~n10842;
  assign n10846 = ~n10845 | ~n10844;
  assign n10847 = ~n10911 & ~n10846;
  assign n10850 = ~n10912 & ~n10847;
  assign n10849 = ~n10848 | ~n10915;
  assign n10851 = ~n10850 & ~n10849;
  assign n10852 = ~n10919 & ~n10851;
  assign n10853 = ~n10921 & ~n10852;
  assign n10854 = ~n10923 & ~n10853;
  assign n10856 = ~n10925 & ~n10854;
  assign n10858 = ~n10856 | ~n10855;
  assign n10859 = ~n10858 | ~n10857;
  assign n10860 = ~n10859 | ~n10885;
  assign n10861 = ~n10932 | ~n10860;
  assign n10863 = ~n10862 | ~n10861;
  assign n10865 = ~n10864 & ~n10863;
  assign n10868 = ~n10866 & ~n10865;
  assign n10869 = ~n10868 & ~n10867;
  assign n10870 = ~n10947 & ~n10869;
  assign n10872 = ~n10871 & ~n10870;
  assign n10873 = ~n10872 | ~n10949;
  assign n10876 = ~n10874 | ~n10873;
  assign n10879 = ~n10876 & ~n10875;
  assign n10877 = ~n10954;
  assign n10878 = ~n10877 | ~n14881;
  assign n10880 = ~n10879 & ~n10878;
  assign n10881 = ~n10880 & ~n11253;
  assign n10953 = ~n10883;
  assign n10939 = ~n10884;
  assign n10929 = ~n10885;
  assign n10890 = ~n10886;
  assign n10889 = ~n10888 | ~n10887;
  assign n10891 = ~n10890 & ~n10889;
  assign n10894 = ~n10891 & ~n11881;
  assign n10893 = ~n10892;
  assign n10897 = ~n10894 & ~n10893;
  assign n10896 = ~n10895;
  assign n10900 = ~n10897 & ~n10896;
  assign n10899 = ~n10898 | ~n12349;
  assign n10902 = ~n10900 & ~n10899;
  assign n10905 = ~n10902 & ~n10901;
  assign n10904 = ~n10903;
  assign n10907 = ~n10905 & ~n10904;
  assign n10908 = ~n10907 & ~n7495;
  assign n10910 = ~n10909 & ~n10908;
  assign n10913 = ~n10911 & ~n10910;
  assign n10917 = ~n10913 & ~n10912;
  assign n10916 = ~n10915 | ~n10914;
  assign n10918 = ~n10917 & ~n10916;
  assign n10920 = ~n10919 & ~n10918;
  assign n10922 = ~n10921 & ~n10920;
  assign n10924 = ~n10923 & ~n10922;
  assign n10927 = ~n10925 & ~n10924;
  assign n10928 = ~n10927 & ~n10926;
  assign n10930 = ~n10929 & ~n10928;
  assign n10933 = ~n10931 | ~n10930;
  assign n10935 = ~n10933 | ~n10932;
  assign n10936 = ~n10935 | ~n10934;
  assign n10938 = ~n10937 & ~n10936;
  assign n10940 = ~n10939 & ~n10938;
  assign n10943 = ~n10941 & ~n10940;
  assign n10944 = ~n10943 & ~n10942;
  assign n10946 = ~n10945 & ~n10944;
  assign n10951 = ~n10947 & ~n10946;
  assign n10950 = ~n10949 | ~n10948;
  assign n10952 = ~n10951 & ~n10950;
  assign n10955 = ~n10953 & ~n10952;
  assign n10959 = ~n10955 & ~n10954;
  assign n10957 = ~n10959 & ~n14881;
  assign n10961 = ~n10959 | ~n10958;
  assign n13170 = ~n10960 & ~P1_U3086;
  assign n11864 = ~n10962;
  assign n10963 = ~n11214 | ~n11864;
  assign n11619 = n7328 | n11612;
  assign n10966 = ~n10963 & ~n11619;
  assign n10964 = ~n13170 | ~n12950;
  assign n10965 = ~n10964 | ~P1_B_REG_SCAN_IN;
  assign input_0 = keyinput_0 ^ SI_31_;
  assign input_1 = keyinput_1 ^ SI_30_;
  assign AND_1 = input_0 & input_1;
  assign input_2 = ~keyinput_2 ^ SI_29_;
  assign AND_2 = input_2 & AND_1;
  assign input_3 = ~keyinput_3 ^ SI_28_;
  assign AND_3 = input_3 & AND_2;
  assign input_4 = ~keyinput_4 ^ SI_27_;
  assign OR_4 = input_4 | AND_3;
  assign input_5 = keyinput_5 ^ SI_26_;
  assign OR_5 = input_5 | OR_4;
  assign input_6 = ~keyinput_6 ^ SI_25_;
  assign OR_6 = input_6 | OR_5;
  assign input_7 = keyinput_7 ^ SI_24_;
  assign OR_7 = input_7 | OR_6;
  assign input_8 = ~keyinput_8 ^ SI_23_;
  assign OR_8 = input_8 | OR_7;
  assign input_9 = ~keyinput_9 ^ SI_22_;
  assign OR_9 = input_9 | OR_8;
  assign input_10 = keyinput_10 ^ SI_21_;
  assign AND_10 = input_10 & OR_9;
  assign input_11 = keyinput_11 ^ SI_20_;
  assign AND_11 = input_11 & AND_10;
  assign input_12 = keyinput_12 ^ SI_19_;
  assign OR_12 = input_12 | AND_11;
  assign input_13 = ~keyinput_13 ^ SI_18_;
  assign AND_13 = input_13 & OR_12;
  assign input_14 = keyinput_14 ^ SI_17_;
  assign OR_14 = input_14 | AND_13;
  assign input_15 = keyinput_15 ^ SI_16_;
  assign AND_15 = input_15 & OR_14;
  assign input_16 = ~keyinput_16 ^ SI_15_;
  assign AND_16 = input_16 & AND_15;
  assign input_17 = ~keyinput_17 ^ SI_14_;
  assign OR_17 = input_17 | AND_16;
  assign input_18 = keyinput_18 ^ SI_13_;
  assign OR_18 = input_18 | OR_17;
  assign input_19 = ~keyinput_19 ^ SI_12_;
  assign AND_19 = input_19 & OR_18;
  assign input_20 = keyinput_20 ^ SI_11_;
  assign AND_20 = input_20 & AND_19;
  assign input_21 = ~keyinput_21 ^ SI_10_;
  assign AND_21 = input_21 & AND_20;
  assign input_22 = keyinput_22 ^ SI_9_;
  assign AND_22 = input_22 & AND_21;
  assign input_23 = ~keyinput_23 ^ SI_8_;
  assign OR_23 = input_23 | AND_22;
  assign input_24 = ~keyinput_24 ^ SI_7_;
  assign OR_24 = input_24 | OR_23;
  assign input_25 = keyinput_25 ^ SI_6_;
  assign AND_25 = input_25 & OR_24;
  assign input_26 = ~keyinput_26 ^ SI_5_;
  assign AND_26 = input_26 & AND_25;
  assign input_27 = ~keyinput_27 ^ SI_4_;
  assign OR_27 = input_27 | AND_26;
  assign input_28 = keyinput_28 ^ SI_3_;
  assign OR_28 = input_28 | OR_27;
  assign input_29 = keyinput_29 ^ SI_2_;
  assign OR_29 = input_29 | OR_28;
  assign input_30 = ~keyinput_30 ^ SI_1_;
  assign AND_30 = input_30 & OR_29;
  assign input_31 = keyinput_31 ^ SI_0_;
  assign AND_31 = input_31 & AND_30;
  assign input_32 = ~keyinput_32 ^ P2_RD_REG_SCAN_IN;
  assign OR_32 = input_32 | AND_31;
  assign input_33 = keyinput_33 ^ P2_DATAO_REG_31__SCAN_IN;
  assign AND_33 = input_33 & OR_32;
  assign input_34 = ~keyinput_34 ^ P2_DATAO_REG_30__SCAN_IN;
  assign AND_34 = input_34 & AND_33;
  assign input_35 = ~keyinput_35 ^ P2_DATAO_REG_29__SCAN_IN;
  assign OR_35 = input_35 | AND_34;
  assign input_36 = ~keyinput_36 ^ P2_DATAO_REG_28__SCAN_IN;
  assign OR_36 = input_36 | OR_35;
  assign input_37 = ~keyinput_37 ^ P2_DATAO_REG_27__SCAN_IN;
  assign OR_37 = input_37 | OR_36;
  assign input_38 = ~keyinput_38 ^ P2_DATAO_REG_26__SCAN_IN;
  assign AND_38 = input_38 & OR_37;
  assign input_39 = keyinput_39 ^ P2_DATAO_REG_25__SCAN_IN;
  assign OR_39 = input_39 | AND_38;
  assign input_40 = ~keyinput_40 ^ P2_DATAO_REG_24__SCAN_IN;
  assign OR_40 = input_40 | OR_39;
  assign input_41 = keyinput_41 ^ P2_DATAO_REG_23__SCAN_IN;
  assign AND_41 = input_41 & OR_40;
  assign input_42 = keyinput_42 ^ P2_DATAO_REG_22__SCAN_IN;
  assign OR_42 = input_42 | AND_41;
  assign input_43 = ~keyinput_43 ^ P2_DATAO_REG_21__SCAN_IN;
  assign OR_43 = input_43 | OR_42;
  assign input_44 = ~keyinput_44 ^ P2_DATAO_REG_20__SCAN_IN;
  assign OR_44 = input_44 | OR_43;
  assign input_45 = keyinput_45 ^ P2_DATAO_REG_19__SCAN_IN;
  assign OR_45 = input_45 | OR_44;
  assign input_46 = ~keyinput_46 ^ P2_DATAO_REG_18__SCAN_IN;
  assign OR_46 = input_46 | OR_45;
  assign input_47 = ~keyinput_47 ^ P2_DATAO_REG_17__SCAN_IN;
  assign OR_47 = input_47 | OR_46;
  assign input_48 = ~keyinput_48 ^ P2_DATAO_REG_16__SCAN_IN;
  assign AND_48 = input_48 & OR_47;
  assign input_49 = ~keyinput_49 ^ P2_DATAO_REG_15__SCAN_IN;
  assign OR_49 = input_49 | AND_48;
  assign input_50 = keyinput_50 ^ P2_DATAO_REG_14__SCAN_IN;
  assign OR_50 = input_50 | OR_49;
  assign input_51 = keyinput_51 ^ P2_DATAO_REG_13__SCAN_IN;
  assign AND_51 = input_51 & OR_50;
  assign input_52 = keyinput_52 ^ P2_DATAO_REG_12__SCAN_IN;
  assign AND_52 = input_52 & AND_51;
  assign input_53 = ~keyinput_53 ^ P2_DATAO_REG_11__SCAN_IN;
  assign AND_53 = input_53 & AND_52;
  assign input_54 = keyinput_54 ^ P2_DATAO_REG_10__SCAN_IN;
  assign AND_54 = input_54 & AND_53;
  assign input_55 = ~keyinput_55 ^ P2_DATAO_REG_9__SCAN_IN;
  assign AND_55 = input_55 & AND_54;
  assign input_56 = keyinput_56 ^ P2_DATAO_REG_8__SCAN_IN;
  assign OR_56 = input_56 | AND_55;
  assign input_57 = keyinput_57 ^ P2_DATAO_REG_7__SCAN_IN;
  assign OR_57 = input_57 | OR_56;
  assign input_58 = keyinput_58 ^ P1_IR_REG_0__SCAN_IN;
  assign AND_58 = input_58 & OR_57;
  assign input_59 = ~keyinput_59 ^ P1_IR_REG_1__SCAN_IN;
  assign OR_59 = input_59 | AND_58;
  assign input_60 = keyinput_60 ^ P1_IR_REG_2__SCAN_IN;
  assign OR_60 = input_60 | OR_59;
  assign input_61 = keyinput_61 ^ P1_IR_REG_3__SCAN_IN;
  assign AND_61 = input_61 & OR_60;
  assign input_62 = ~keyinput_62 ^ P1_IR_REG_4__SCAN_IN;
  assign OR_62 = input_62 | AND_61;
  assign input_63 = ~keyinput_63 ^ P1_IR_REG_5__SCAN_IN;
  assign OR_63 = input_63 | OR_62;
  assign input_64 = ~keyinput_64 ^ P1_IR_REG_6__SCAN_IN;
  assign AND_64 = input_64 & OR_63;
  assign input_65 = keyinput_65 ^ P1_IR_REG_7__SCAN_IN;
  assign AND_65 = input_65 & AND_64;
  assign input_66 = keyinput_66 ^ P1_IR_REG_8__SCAN_IN;
  assign AND_66 = input_66 & AND_65;
  assign input_67 = ~keyinput_67 ^ P1_IR_REG_9__SCAN_IN;
  assign AND_67 = input_67 & AND_66;
  assign input_68 = keyinput_68 ^ P1_IR_REG_10__SCAN_IN;
  assign AND_68 = input_68 & AND_67;
  assign input_69 = keyinput_69 ^ P1_IR_REG_11__SCAN_IN;
  assign AND_69 = input_69 & AND_68;
  assign input_70 = ~keyinput_70 ^ P1_IR_REG_12__SCAN_IN;
  assign AND_70 = input_70 & AND_69;
  assign input_71 = ~keyinput_71 ^ P1_IR_REG_13__SCAN_IN;
  assign AND_71 = input_71 & AND_70;
  assign input_72 = keyinput_72 ^ P1_IR_REG_14__SCAN_IN;
  assign OR_72 = input_72 | AND_71;
  assign input_73 = ~keyinput_73 ^ P1_IR_REG_15__SCAN_IN;
  assign OR_73 = input_73 | OR_72;
  assign input_74 = keyinput_74 ^ P1_IR_REG_16__SCAN_IN;
  assign AND_74 = input_74 & OR_73;
  assign input_75 = keyinput_75 ^ P1_IR_REG_17__SCAN_IN;
  assign OR_75 = input_75 | AND_74;
  assign input_76 = ~keyinput_76 ^ P1_IR_REG_18__SCAN_IN;
  assign AND_76 = input_76 & OR_75;
  assign input_77 = ~keyinput_77 ^ P1_IR_REG_19__SCAN_IN;
  assign OR_77 = input_77 | AND_76;
  assign input_78 = ~keyinput_78 ^ P1_IR_REG_20__SCAN_IN;
  assign AND_78 = input_78 & OR_77;
  assign input_79 = ~keyinput_79 ^ P1_IR_REG_21__SCAN_IN;
  assign AND_79 = input_79 & AND_78;
  assign input_80 = keyinput_80 ^ SI_31_;
  assign input_81 = keyinput_81 ^ SI_30_;
  assign AND_81 = input_80 & input_81;
  assign input_82 = keyinput_82 ^ SI_29_;
  assign AND_82 = input_82 & AND_81;
  assign input_83 = ~keyinput_83 ^ SI_28_;
  assign AND_83 = input_83 & AND_82;
  assign input_84 = ~keyinput_84 ^ SI_27_;
  assign OR_84 = input_84 | AND_83;
  assign input_85 = keyinput_85 ^ SI_26_;
  assign OR_85 = input_85 | OR_84;
  assign input_86 = keyinput_86 ^ SI_25_;
  assign OR_86 = input_86 | OR_85;
  assign input_87 = ~keyinput_87 ^ SI_24_;
  assign OR_87 = input_87 | OR_86;
  assign input_88 = ~keyinput_88 ^ SI_23_;
  assign OR_88 = input_88 | OR_87;
  assign input_89 = keyinput_89 ^ SI_22_;
  assign OR_89 = input_89 | OR_88;
  assign input_90 = ~keyinput_90 ^ SI_21_;
  assign AND_90 = input_90 & OR_89;
  assign input_91 = keyinput_91 ^ SI_20_;
  assign AND_91 = input_91 & AND_90;
  assign input_92 = ~keyinput_92 ^ SI_19_;
  assign OR_92 = input_92 | AND_91;
  assign input_93 = keyinput_93 ^ SI_18_;
  assign AND_93 = input_93 & OR_92;
  assign input_94 = ~keyinput_94 ^ SI_17_;
  assign OR_94 = input_94 | AND_93;
  assign input_95 = keyinput_95 ^ SI_16_;
  assign AND_95 = input_95 & OR_94;
  assign input_96 = ~keyinput_96 ^ SI_15_;
  assign AND_96 = input_96 & AND_95;
  assign input_97 = ~keyinput_97 ^ SI_14_;
  assign OR_97 = input_97 | AND_96;
  assign input_98 = ~keyinput_98 ^ SI_13_;
  assign OR_98 = input_98 | OR_97;
  assign input_99 = ~keyinput_99 ^ SI_12_;
  assign AND_99 = input_99 & OR_98;
  assign input_100 = ~keyinput_100 ^ SI_11_;
  assign AND_100 = input_100 & AND_99;
  assign input_101 = ~keyinput_101 ^ SI_10_;
  assign AND_101 = input_101 & AND_100;
  assign input_102 = keyinput_102 ^ SI_9_;
  assign AND_102 = input_102 & AND_101;
  assign input_103 = ~keyinput_103 ^ SI_8_;
  assign OR_103 = input_103 | AND_102;
  assign input_104 = ~keyinput_104 ^ SI_7_;
  assign OR_104 = input_104 | OR_103;
  assign input_105 = ~keyinput_105 ^ SI_6_;
  assign AND_105 = input_105 & OR_104;
  assign input_106 = ~keyinput_106 ^ SI_5_;
  assign AND_106 = input_106 & AND_105;
  assign input_107 = ~keyinput_107 ^ SI_4_;
  assign OR_107 = input_107 | AND_106;
  assign input_108 = keyinput_108 ^ SI_3_;
  assign OR_108 = input_108 | OR_107;
  assign input_109 = ~keyinput_109 ^ SI_2_;
  assign OR_109 = input_109 | OR_108;
  assign input_110 = ~keyinput_110 ^ SI_1_;
  assign AND_110 = input_110 & OR_109;
  assign input_111 = ~keyinput_111 ^ SI_0_;
  assign AND_111 = input_111 & AND_110;
  assign input_112 = keyinput_112 ^ P2_RD_REG_SCAN_IN;
  assign OR_112 = input_112 | AND_111;
  assign input_113 = ~keyinput_113 ^ P2_DATAO_REG_31__SCAN_IN;
  assign AND_113 = input_113 & OR_112;
  assign input_114 = keyinput_114 ^ P2_DATAO_REG_30__SCAN_IN;
  assign AND_114 = input_114 & AND_113;
  assign input_115 = keyinput_115 ^ P2_DATAO_REG_29__SCAN_IN;
  assign OR_115 = input_115 | AND_114;
  assign input_116 = ~keyinput_116 ^ P2_DATAO_REG_28__SCAN_IN;
  assign OR_116 = input_116 | OR_115;
  assign input_117 = keyinput_117 ^ P2_DATAO_REG_27__SCAN_IN;
  assign OR_117 = input_117 | OR_116;
  assign input_118 = ~keyinput_118 ^ P2_DATAO_REG_26__SCAN_IN;
  assign AND_118 = input_118 & OR_117;
  assign input_119 = ~keyinput_119 ^ P2_DATAO_REG_25__SCAN_IN;
  assign OR_119 = input_119 | AND_118;
  assign input_120 = keyinput_120 ^ P2_DATAO_REG_24__SCAN_IN;
  assign OR_120 = input_120 | OR_119;
  assign input_121 = keyinput_121 ^ P2_DATAO_REG_23__SCAN_IN;
  assign AND_121 = input_121 & OR_120;
  assign input_122 = keyinput_122 ^ P2_DATAO_REG_22__SCAN_IN;
  assign OR_122 = input_122 | AND_121;
  assign input_123 = keyinput_123 ^ P2_DATAO_REG_21__SCAN_IN;
  assign OR_123 = input_123 | OR_122;
  assign input_124 = keyinput_124 ^ P2_DATAO_REG_20__SCAN_IN;
  assign OR_124 = input_124 | OR_123;
  assign input_125 = keyinput_125 ^ P2_DATAO_REG_19__SCAN_IN;
  assign OR_125 = input_125 | OR_124;
  assign input_126 = ~keyinput_126 ^ P2_DATAO_REG_18__SCAN_IN;
  assign OR_126 = input_126 | OR_125;
  assign input_127 = ~keyinput_127 ^ P2_DATAO_REG_17__SCAN_IN;
  assign OR_127 = input_127 | OR_126;
  assign input_128 = ~keyinput_128 ^ P2_DATAO_REG_16__SCAN_IN;
  assign AND_128 = input_128 & OR_127;
  assign input_129 = ~keyinput_129 ^ P2_DATAO_REG_15__SCAN_IN;
  assign OR_129 = input_129 | AND_128;
  assign input_130 = ~keyinput_130 ^ P2_DATAO_REG_14__SCAN_IN;
  assign OR_130 = input_130 | OR_129;
  assign input_131 = keyinput_131 ^ P2_DATAO_REG_13__SCAN_IN;
  assign AND_131 = input_131 & OR_130;
  assign input_132 = keyinput_132 ^ P2_DATAO_REG_12__SCAN_IN;
  assign AND_132 = input_132 & AND_131;
  assign input_133 = keyinput_133 ^ P2_DATAO_REG_11__SCAN_IN;
  assign AND_133 = input_133 & AND_132;
  assign input_134 = ~keyinput_134 ^ P2_DATAO_REG_10__SCAN_IN;
  assign AND_134 = input_134 & AND_133;
  assign input_135 = keyinput_135 ^ P2_DATAO_REG_9__SCAN_IN;
  assign AND_135 = input_135 & AND_134;
  assign input_136 = ~keyinput_136 ^ P2_DATAO_REG_8__SCAN_IN;
  assign OR_136 = input_136 | AND_135;
  assign input_137 = ~keyinput_137 ^ P2_DATAO_REG_7__SCAN_IN;
  assign OR_137 = input_137 | OR_136;
  assign input_138 = keyinput_138 ^ P1_IR_REG_0__SCAN_IN;
  assign AND_138 = input_138 & OR_137;
  assign input_139 = keyinput_139 ^ P1_IR_REG_1__SCAN_IN;
  assign OR_139 = input_139 | AND_138;
  assign input_140 = ~keyinput_140 ^ P1_IR_REG_2__SCAN_IN;
  assign OR_140 = input_140 | OR_139;
  assign input_141 = ~keyinput_141 ^ P1_IR_REG_3__SCAN_IN;
  assign AND_141 = input_141 & OR_140;
  assign input_142 = ~keyinput_142 ^ P1_IR_REG_4__SCAN_IN;
  assign OR_142 = input_142 | AND_141;
  assign input_143 = ~keyinput_143 ^ P1_IR_REG_5__SCAN_IN;
  assign OR_143 = input_143 | OR_142;
  assign input_144 = keyinput_144 ^ P1_IR_REG_6__SCAN_IN;
  assign AND_144 = input_144 & OR_143;
  assign input_145 = ~keyinput_145 ^ P1_IR_REG_7__SCAN_IN;
  assign AND_145 = input_145 & AND_144;
  assign input_146 = ~keyinput_146 ^ P1_IR_REG_8__SCAN_IN;
  assign AND_146 = input_146 & AND_145;
  assign input_147 = ~keyinput_147 ^ P1_IR_REG_9__SCAN_IN;
  assign AND_147 = input_147 & AND_146;
  assign input_148 = ~keyinput_148 ^ P1_IR_REG_10__SCAN_IN;
  assign AND_148 = input_148 & AND_147;
  assign input_149 = ~keyinput_149 ^ P1_IR_REG_11__SCAN_IN;
  assign AND_149 = input_149 & AND_148;
  assign input_150 = keyinput_150 ^ P1_IR_REG_12__SCAN_IN;
  assign AND_150 = input_150 & AND_149;
  assign input_151 = keyinput_151 ^ P1_IR_REG_13__SCAN_IN;
  assign AND_151 = input_151 & AND_150;
  assign input_152 = keyinput_152 ^ P1_IR_REG_14__SCAN_IN;
  assign OR_152 = input_152 | AND_151;
  assign input_153 = ~keyinput_153 ^ P1_IR_REG_15__SCAN_IN;
  assign OR_153 = input_153 | OR_152;
  assign input_154 = keyinput_154 ^ P1_IR_REG_16__SCAN_IN;
  assign AND_154 = input_154 & OR_153;
  assign input_155 = keyinput_155 ^ P1_IR_REG_17__SCAN_IN;
  assign OR_155 = input_155 | AND_154;
  assign input_156 = keyinput_156 ^ P1_IR_REG_18__SCAN_IN;
  assign AND_156 = input_156 & OR_155;
  assign input_157 = ~keyinput_157 ^ P1_IR_REG_19__SCAN_IN;
  assign OR_157 = input_157 | AND_156;
  assign input_158 = keyinput_158 ^ P1_IR_REG_20__SCAN_IN;
  assign AND_158 = input_158 & OR_157;
  assign input_159 = ~keyinput_159 ^ P1_IR_REG_21__SCAN_IN;
  assign AND_159 = input_159 & AND_158;
  assign AND_159_INV = ~AND_159;
  assign CASOP = AND_79 & AND_159_INV;
  assign P1_U3242 = P1_U3242_Lock ^ CASOP;
endmodule


