// Benchmark "b17_C_lock" written by ABC on Thu May 13 23:44:09 2021

module b17_C_lock ( 
    keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
    keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
    keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
    keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
    keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
    keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
    keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
    keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
    keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
    keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
    keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
    keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
    keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
    keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
    keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
    keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
    keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
    keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
    keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
    keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
    keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
    keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
    keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
    keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
    keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
    keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
    keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
    keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
    keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
    keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
    keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
    keyinput_156, keyinput_157, keyinput_158, keyinput_159,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, P2_STATE_REG_2__SCAN_IN,
    P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
    P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
    P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
    P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
    P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
    P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
    P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
    P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
    P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
    P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
    P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
    P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
    P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
    P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
    P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
    P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
    P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
    P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
    P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
    P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
    P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
    P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
    P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
    P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
    P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
    P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
    P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
    P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
    P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
    P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
    P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
    P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
    P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
    P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
    P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
    P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
    P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
    P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
    P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
    P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
    P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
    P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
    P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
    P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
    P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
    P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
    P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
    P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
    P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
    P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
    P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
    P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
    P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
    P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
    P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
    P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
    P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
    P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
    P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
    P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
    P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
    P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
    P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
    P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
    P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
    P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
    P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN,
    P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_INSTADDRPOINTER_REG_3__SCAN_IN,
    P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_INSTADDRPOINTER_REG_5__SCAN_IN,
    P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_INSTADDRPOINTER_REG_7__SCAN_IN,
    P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_INSTADDRPOINTER_REG_9__SCAN_IN,
    P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_INSTADDRPOINTER_REG_11__SCAN_IN,
    P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_INSTADDRPOINTER_REG_13__SCAN_IN,
    P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_INSTADDRPOINTER_REG_15__SCAN_IN,
    P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_INSTADDRPOINTER_REG_17__SCAN_IN,
    P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_INSTADDRPOINTER_REG_19__SCAN_IN,
    P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_INSTADDRPOINTER_REG_21__SCAN_IN,
    P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_INSTADDRPOINTER_REG_23__SCAN_IN,
    P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_INSTADDRPOINTER_REG_25__SCAN_IN,
    P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_INSTADDRPOINTER_REG_27__SCAN_IN,
    P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_INSTADDRPOINTER_REG_29__SCAN_IN,
    P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_INSTADDRPOINTER_REG_31__SCAN_IN,
    P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_PHYADDRPOINTER_REG_1__SCAN_IN,
    P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_PHYADDRPOINTER_REG_3__SCAN_IN,
    P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_PHYADDRPOINTER_REG_5__SCAN_IN,
    P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_PHYADDRPOINTER_REG_7__SCAN_IN,
    P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_PHYADDRPOINTER_REG_9__SCAN_IN,
    P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_PHYADDRPOINTER_REG_11__SCAN_IN,
    P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_PHYADDRPOINTER_REG_13__SCAN_IN,
    P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_PHYADDRPOINTER_REG_15__SCAN_IN,
    P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_PHYADDRPOINTER_REG_17__SCAN_IN,
    P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_PHYADDRPOINTER_REG_19__SCAN_IN,
    P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_PHYADDRPOINTER_REG_21__SCAN_IN,
    P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_PHYADDRPOINTER_REG_23__SCAN_IN,
    P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_PHYADDRPOINTER_REG_25__SCAN_IN,
    P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_PHYADDRPOINTER_REG_27__SCAN_IN,
    P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_PHYADDRPOINTER_REG_29__SCAN_IN,
    P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_PHYADDRPOINTER_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, P2_FLUSH_REG_SCAN_IN,
    P2_U3015  );
  input  keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4,
    keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9,
    keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14,
    keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19,
    keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24,
    keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29,
    keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34,
    keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39,
    keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44,
    keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49,
    keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54,
    keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59,
    keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64,
    keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69,
    keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74,
    keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79,
    keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84,
    keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89,
    keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94,
    keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99,
    keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104,
    keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109,
    keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114,
    keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119,
    keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124,
    keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129,
    keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134,
    keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139,
    keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144,
    keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149,
    keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154,
    keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, P2_STATE_REG_2__SCAN_IN,
    P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
    P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
    P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
    P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
    P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
    P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
    P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
    P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
    P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
    P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
    P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
    P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
    P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
    P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
    P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
    P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
    P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
    P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
    P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
    P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
    P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
    P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
    P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
    P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
    P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
    P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
    P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
    P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
    P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
    P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
    P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
    P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
    P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
    P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
    P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
    P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
    P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
    P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
    P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
    P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
    P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
    P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
    P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
    P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
    P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
    P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
    P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
    P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
    P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
    P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
    P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
    P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
    P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
    P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
    P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
    P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
    P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
    P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
    P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
    P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
    P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
    P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
    P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
    P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
    P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
    P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
    P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_1__SCAN_IN,
    P2_INSTADDRPOINTER_REG_2__SCAN_IN, P2_INSTADDRPOINTER_REG_3__SCAN_IN,
    P2_INSTADDRPOINTER_REG_4__SCAN_IN, P2_INSTADDRPOINTER_REG_5__SCAN_IN,
    P2_INSTADDRPOINTER_REG_6__SCAN_IN, P2_INSTADDRPOINTER_REG_7__SCAN_IN,
    P2_INSTADDRPOINTER_REG_8__SCAN_IN, P2_INSTADDRPOINTER_REG_9__SCAN_IN,
    P2_INSTADDRPOINTER_REG_10__SCAN_IN, P2_INSTADDRPOINTER_REG_11__SCAN_IN,
    P2_INSTADDRPOINTER_REG_12__SCAN_IN, P2_INSTADDRPOINTER_REG_13__SCAN_IN,
    P2_INSTADDRPOINTER_REG_14__SCAN_IN, P2_INSTADDRPOINTER_REG_15__SCAN_IN,
    P2_INSTADDRPOINTER_REG_16__SCAN_IN, P2_INSTADDRPOINTER_REG_17__SCAN_IN,
    P2_INSTADDRPOINTER_REG_18__SCAN_IN, P2_INSTADDRPOINTER_REG_19__SCAN_IN,
    P2_INSTADDRPOINTER_REG_20__SCAN_IN, P2_INSTADDRPOINTER_REG_21__SCAN_IN,
    P2_INSTADDRPOINTER_REG_22__SCAN_IN, P2_INSTADDRPOINTER_REG_23__SCAN_IN,
    P2_INSTADDRPOINTER_REG_24__SCAN_IN, P2_INSTADDRPOINTER_REG_25__SCAN_IN,
    P2_INSTADDRPOINTER_REG_26__SCAN_IN, P2_INSTADDRPOINTER_REG_27__SCAN_IN,
    P2_INSTADDRPOINTER_REG_28__SCAN_IN, P2_INSTADDRPOINTER_REG_29__SCAN_IN,
    P2_INSTADDRPOINTER_REG_30__SCAN_IN, P2_INSTADDRPOINTER_REG_31__SCAN_IN,
    P2_PHYADDRPOINTER_REG_0__SCAN_IN, P2_PHYADDRPOINTER_REG_1__SCAN_IN,
    P2_PHYADDRPOINTER_REG_2__SCAN_IN, P2_PHYADDRPOINTER_REG_3__SCAN_IN,
    P2_PHYADDRPOINTER_REG_4__SCAN_IN, P2_PHYADDRPOINTER_REG_5__SCAN_IN,
    P2_PHYADDRPOINTER_REG_6__SCAN_IN, P2_PHYADDRPOINTER_REG_7__SCAN_IN,
    P2_PHYADDRPOINTER_REG_8__SCAN_IN, P2_PHYADDRPOINTER_REG_9__SCAN_IN,
    P2_PHYADDRPOINTER_REG_10__SCAN_IN, P2_PHYADDRPOINTER_REG_11__SCAN_IN,
    P2_PHYADDRPOINTER_REG_12__SCAN_IN, P2_PHYADDRPOINTER_REG_13__SCAN_IN,
    P2_PHYADDRPOINTER_REG_14__SCAN_IN, P2_PHYADDRPOINTER_REG_15__SCAN_IN,
    P2_PHYADDRPOINTER_REG_16__SCAN_IN, P2_PHYADDRPOINTER_REG_17__SCAN_IN,
    P2_PHYADDRPOINTER_REG_18__SCAN_IN, P2_PHYADDRPOINTER_REG_19__SCAN_IN,
    P2_PHYADDRPOINTER_REG_20__SCAN_IN, P2_PHYADDRPOINTER_REG_21__SCAN_IN,
    P2_PHYADDRPOINTER_REG_22__SCAN_IN, P2_PHYADDRPOINTER_REG_23__SCAN_IN,
    P2_PHYADDRPOINTER_REG_24__SCAN_IN, P2_PHYADDRPOINTER_REG_25__SCAN_IN,
    P2_PHYADDRPOINTER_REG_26__SCAN_IN, P2_PHYADDRPOINTER_REG_27__SCAN_IN,
    P2_PHYADDRPOINTER_REG_28__SCAN_IN, P2_PHYADDRPOINTER_REG_29__SCAN_IN,
    P2_PHYADDRPOINTER_REG_30__SCAN_IN, P2_PHYADDRPOINTER_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, P2_FLUSH_REG_SCAN_IN;
  output P2_U3015;
  wire n34982, n21475, n40626, n26095, n20338, n30005, n25608, n21353,
    n26187, n21498, n25836, n21791, n25810, n20333, n22568, n34908, n21369,
    n25478, n40860, n20337, n21268, n21253, n26070, n40817, n34001, n25616,
    n20332, n22371, n35516, n25531, n40702, n39539, n36597, n34713, n21505,
    n35866, n21480, n20827, n21476, n21519, n20618, n20623, n35527, n35075,
    n33203, n21471, n21464, n21458, n22379, n22155, n27051, n21373, n21415,
    n21361, n21330, n22389, n22360, n21354, n22153, n22088, n35031, n22370,
    n21362, n21265, n21327, n21320, n21170, n20339, n26132, n21212, n21313,
    n21549, n22222, n26137, n21312, n40788, n26169, n34008, n34021, n33988,
    n25782, n22328, n25822, n25513, n21779, n20353, n20354, n21404, n21666,
    n21851, n21377, n20656, n20657, n22181, n20512, n20507, n20508, n20509,
    n20708, n20710, n20785, n20786, n34467, n38064, n21197, n21754, n20782,
    n21753, n20783, n21496, n20824, n20823, n20712, n22323, n21384, n21407,
    n21399, n21300, n20997, n20585, n20791, n21762, n20825, n21860, n21755,
    n20501, n21836, n27052, n20800, n20795, n21225, n25218, n25206, n21927,
    n21872, n20511, n20967, n21444, n21965, n21438, n20648, n31666, n25485,
    n20787, n20554, n27013, n20688, n21520, n20624, n20799, n21459, n20801,
    n21164, n21194, n29331, n29333, n20660, n20703, n37916, n20555, n20556,
    n34233, n20550, n20694, n20639, n20640, n25379, n25334, n20638, n37331,
    n20692, n20691, n40719, n40931, n21695, n21623, n26175, n20634, n20635,
    n20636, n20637, n20933, n21497, n20923, n40469, n21176, n21391, n21352,
    n21333, n21198, n21210, n21204, n21224, n21889, n21885, n20951, n21840,
    n21833, n20504, n26066, n21395, n26147, n26100, n25182, n21913, n20713,
    n21857, n21856, n20584, n21751, n20876, n21450, n20877, n21456, n21457,
    n21501, n20689, n21512, n20705, n25332, n25240, n25215, n21921, n20714,
    n20715, n21896, n21894, n21888, n20707, n21845, n20704, n21443, n21425,
    n21423, n20882, n25364, n25312, n25854, n33607, n21376, n21303, n20872,
    n20873, n21014, n25441, n20869, n20870, n20697, n38068, n26215, n25280,
    n35684, n35691, n35501, n25167, n34622, n20878, n40137, n35671, n35358,
    n33140, n32109, n31875, n22176, n20655, n21858, n25968, n25974, n20662,
    n21756, n36596, n33541, n22420, n20647, n21245, n25475, n37920, n20510,
    n25222, n21879, n21878, n21880, n20981, n20701, n20702, n38250, n34624,
    n20552, n20553, n32963, n33551, n34510, n21461, n21441, n21442, n25693,
    n35494, n20794, n20695, n20696, n25238, n20643, n25237, n25209, n25174,
    n35952, n40118, n20690, n21247, n21544, n26048, n20952, n20359, n20360,
    n20361, n20363, n20364, n20788, n21257, n20377, n20378, n20379, n20381,
    n20383, n21148, n20386, n20387, n20389, n20706, n20394, n20396, n20398,
    n30599, n21004, n22341, n20402, n20406, n21842, n20413, n20414, n20415,
    n20416, n20418, n20423, n20424, n20426, n20427, n20428, n20430, n20432,
    n20438, n20442, n20443, n20444, n20447, n34004, n20450, n21925, n20455,
    n22361, n20505, n20456, n20460, n20467, n20468, n21972, n20617, n25440,
    n20709, n40929, n20471, n20483, n37335, n20485, n20831, n25219, n20506,
    n21919, n20513, n20551, n20578, n34716, n21737, n20582, n20579, n20580,
    n20581, n20644, n40212, n20590, n34839, n20619, n20620, n22027, n20798,
    n38451, n20646, n20826, n25257, n25383, n20632, n20641, n40161, n21914,
    n20645, n22380, n30480, n37914, n26982, n20649, n20650, n20658, n22422,
    n20659, n25415, n20687, n20693, n25501, n20700, n25496, n21773, n21853,
    n20711, n21823, n21832, n20784, n21750, n21761, n20790, n20822, n20796,
    n21509, n34064, n20797, n21241, n21207, n21141, n21278, n20993, n20962,
    n26167, n20875, n20879, n20881, n21446, n21418, n20883, n20884, n25443,
    n30816, n21226, n20890, n25486, n22194, n20896, n22571, n20898, n20900,
    n20901, n20903, n21759, n20904, n21147, n21256, n22285, n25753, n21206,
    n20984, n20985, n21357, n21234, n21231, n20910, n20960, n21454, n21274,
    n21057, n21871, n25488, n25565, n21365, n21439, n21263, n25389, n21906,
    n21766, n25514, n21859, n40439, n33655, n25970, n21460, n22122, n22143,
    n25472, n36439, n32242, n22174, n34075, n36540, n41068, n40868, n40691,
    n34028, n21056, n21018, n21017, n20909, n21053, n21051, n20913, n20911,
    n20912, n21123, n21122, n21125, n21447, n20914, n20916, n34046, n20915,
    n22120, n21019, n20918, n20917, n20922, n20920, n26069, n20919, n20921,
    n20949, n20953, n20928, n20924, n25799, n20926, n25794, n35840, n20925,
    n20927, n20930, n26127, n20929, n20947, n20932, n20931, n20937, n26146,
    n20935, n20934, n20936, n20945, n40820, n20939, n20938, n20943, n20941,
    n20940, n20942, n20944, n20946, n20948, n31893, n20950, n20958, n20955,
    n20954, n20956, n22324, n20957, n20961, n20959, n20965, n20963, n20964,
    n20966, n20969, n20968, n20973, n20971, n20970, n20972, n20979, n20975,
    n20974, n20977, n20976, n20978, n20980, n20983, n20982, n21474, n20990,
    n20988, n20986, n20987, n20989, n20998, n20992, n39604, n20991, n20996,
    n21469, n20994, n20995, n21000, n20999, n21003, n21001, n21002, n21012,
    n21006, n21005, n21010, n21008, n21007, n21009, n21011, n21013, n25564,
    n21016, n21943, n21015, n21827, n21942, n21949, n21055, n21021, n21020,
    n21025, n21023, n21022, n21024, n21033, n21027, n21026, n21031, n21029,
    n21028, n21030, n21032, n21050, n21035, n21034, n21039, n21037, n21036,
    n21038, n21048, n21041, n25744, n21040, n21046, n21044, n21042, n21535,
    n21043, n21045, n21047, n21049, n21745, n21054, n21052, n21951, n21936,
    n21128, n21091, n21059, n21058, n21063, n21061, n21060, n21062, n21069,
    n25783, n21065, n21648, n21064, n21067, n40482, n21066, n21068, n21089,
    n21071, n40468, n21070, n21077, n22211, n22246, n21075, n21073, n21072,
    n21074, n21076, n21087, n21079, n21152, n21078, n21085, n21080, n21083,
    n21081, n21082, n21084, n21086, n21088, n21736, n21090, n21780, n21093,
    n21092, n21097, n21095, n21094, n21096, n21105, n21099, n21098, n21103,
    n21101, n21100, n21102, n21104, n21121, n21107, n21106, n21111, n21109,
    n21108, n21110, n21119, n21113, n21112, n21117, n21115, n21114, n21116,
    n21118, n21120, n22396, n21127, n21124, n21332, n21126, n21776, n21939,
    n21129, n30072, n21331, n21131, n21130, n21133, n22247, n21132, n21137,
    n21135, n21134, n21136, n21146, n21140, n21138, n21139, n21144, n22250,
    n21142, n21143, n21145, n21151, n21149, n21321, n21150, n21154, n21153,
    n21162, n21156, n21155, n21160, n21158, n21157, n21159, n21161, n21163,
    n21166, n21165, n21168, n21674, n21167, n21169, n21173, n21171, n21172,
    n21181, n21175, n21792, n21174, n21179, n22207, n21177, n40787, n21178,
    n21180, n21183, n21182, n21185, n22208, n21184, n21193, n21187, n21186,
    n21191, n21189, n21188, n21190, n21192, n34924, n21227, n21196, n21195,
    n21611, n21202, n21200, n21199, n21201, n21211, n21205, n21203, n21209,
    n21615, n21208, n21214, n21213, n21218, n21216, n21215, n21217, n21220,
    n21219, n21222, n21221, n21223, n21229, n21228, n21232, n21230, n21237,
    n21233, n21235, n21236, n21246, n21239, n22288, n21238, n21244, n21240,
    n21242, n21243, n21249, n21248, n21252, n21250, n21251, n21255, n21254,
    n21261, n21259, n21258, n21260, n21262, n21264, n34783, n21267, n21266,
    n21270, n25821, n21269, n21271, n21272, n21273, n21283, n21277, n21275,
    n21276, n21281, n21580, n21279, n21280, n21282, n21298, n21285, n21284,
    n21288, n21286, n21287, n21296, n21290, n21289, n21294, n21292, n21291,
    n21293, n21295, n21297, n21301, n21299, n21302, n21304, n26136, n21311,
    n21306, n21305, n21309, n21307, n21308, n21310, n21329, n40816, n21315,
    n40839, n21314, n21319, n40838, n21317, n21316, n21318, n21323, n21322,
    n21325, n21324, n21326, n21328, n25855, n30492, n29786, n34035, n22114,
    n21959, n21335, n21334, n21338, n21337, n21336, n29821, n21339, n21343,
    n21340, n21341, n30489, n21342, n22100, n30086, n34609, n29819, n34083,
    n40434, n40368, n40109, n21390, n21351, n21374, n22175, n33974, n21355,
    n21356, n21359, n21358, n21360, n21934, n26203, n21363, n21364, n25610,
    n22132, n21366, n22139, n21367, n21368, n29336, n25448, n21370, n21403,
    n25847, n21371, n22103, n35016, n22110, n21372, n22147, n21375, n22135,
    n21405, n22136, n21383, n25690, n21378, n21381, n21431, n34078, n21379,
    n21380, n21382, n21386, n21385, n21401, n21387, n21389, n25691, n21388,
    n22142, n21393, n21392, n21394, n21397, n21396, n21398, n21400, n21402,
    n21406, n21412, n25583, n30495, n21410, n21408, n21409, n21411, n21463,
    n21413, n27016, n21414, n21416, n34005, n21417, n21426, n21420, n21419,
    n21427, n21421, n21422, n21424, n21429, n21428, n21430, n21434, n21432,
    n21433, n21435, n21440, n21436, n21437, n21445, n21449, n21448, n34831,
    n21455, n21451, n21453, n21452, n21462, n21466, n21465, n21467, n21468,
    n36849, n21470, n21472, n21473, n35590, n21478, n21477, n35376, n21479,
    n21481, n34862, n21482, n21486, n21483, n36500, n21484, n21485, n21494,
    n21487, n36170, n21488, n21492, n21489, n36075, n21490, n21491, n21493,
    n21495, n21508, n36457, n21500, n37332, n21499, n21506, n36552, n21504,
    n21502, n21503, n21507, n21526, n21510, n37718, n39591, n21511, n21516,
    n21513, n35265, n21514, n21515, n21518, n21517, n21524, n35843, n21522,
    n34805, n21521, n21523, n21525, n21562, n21528, n21527, n21532, n21530,
    n21529, n21531, n21541, n21534, n21533, n21539, n21537, n21536, n21538,
    n21540, n21559, n21543, n21542, n21548, n21546, n21545, n21547, n21557,
    n21551, n21550, n21555, n21553, n25827, n21552, n21554, n21556, n21558,
    n21560, n21743, n22382, n21561, n21564, n21563, n21567, n21566, n21565,
    n21588, n21570, n21568, n21569, n21575, n21571, n21573, n25818, n21572,
    n21574, n21586, n21576, n21579, n21577, n21578, n21584, n25817, n21582,
    n21581, n21583, n21585, n21587, n21596, n21590, n21589, n21594, n21592,
    n21591, n21593, n21595, n22359, n21667, n21598, n21597, n21602, n21600,
    n21599, n21601, n21603, n21605, n40631, n21604, n21610, n21606, n21608,
    n21651, n21607, n21609, n21621, n26065, n21613, n21612, n21619, n21614,
    n21617, n21616, n21618, n21620, n21622, n21631, n21625, n21624, n21629,
    n21627, n21626, n21628, n21630, n21665, n21633, n21632, n21637, n21635,
    n21634, n21636, n21645, n21639, n21638, n21643, n21641, n21640, n21642,
    n21644, n21663, n21647, n21646, n21650, n21649, n21655, n21653, n21652,
    n21654, n21661, n21657, n21656, n21659, n21658, n21660, n21662, n22408,
    n21664, n21669, n21668, n21673, n21671, n21670, n21672, n21676, n21675,
    n21682, n21677, n21680, n21678, n21679, n21681, n21693, n21683, n21686,
    n21684, n21685, n21691, n21687, n21689, n40773, n21688, n21690, n21692,
    n21694, n21703, n21697, n21696, n21701, n21699, n21698, n21700, n21702,
    n21758, n21704, n21706, n21705, n21710, n21708, n21707, n21709, n21718,
    n21712, n21711, n21716, n21714, n21713, n21715, n21717, n21735, n21719,
    n21723, n21721, n21720, n21722, n21727, n21725, n21724, n21726, n21733,
    n21731, n21729, n21728, n21730, n21732, n21734, n21765, n39141, n21738,
    n31887, n21741, n25658, n21739, n21740, n21742, n21747, n31245, n21744,
    n31244, n21746, n21748, n34717, n21749, n21752, n36591, n21757, n36592,
    n21760, n25965, n21763, n21764, n39136, n26977, n40398, n40318, n40409,
    n40103, n40107, n40384, n40360, n40153, n21767, n40328, n22167, n22169,
    n40573, n21768, n21772, n21775, n21774, n21778, n21777, n21822, n21782,
    n21781, n21838, n21784, n38471, n21783, n21844, n21786, n21785, n21790,
    n21788, n21787, n21789, n21816, n21796, n21794, n21793, n21795, n21798,
    n21797, n21814, n21800, n21799, n21804, n21802, n21801, n21803, n21812,
    n21806, n21805, n21810, n21808, n21807, n21809, n21811, n21813, n21815,
    n22358, n21817, n21819, n21818, n21852, n21821, n35557, n21820, n21866,
    n21893, n21863, n21901, n21907, n21911, n21918, n21916, n21926, n25205,
    n37860, n25227, n21824, n37025, n21825, n21826, n35534, n21831, n31882,
    n21829, n21828, n35510, n31881, n21830, n31242, n38436, n31243, n21835,
    n21834, n34712, n21837, n21839, n38663, n35084, n35090, n21841, n21843,
    n21847, n21846, n38476, n21848, n21850, n21849, n25973, n21854, n37882,
    n21855, n21861, n35556, n38853, n38688, n21862, n21870, n21864, n38705,
    n40020, n40290, n40012, n21865, n40123, n21867, n37662, n39536, n39714,
    n21868, n40025, n21869, n21877, n21874, n21873, n37679, n40000, n21876,
    n21875, n40027, n21882, n21881, n38765, n40125, n21884, n40021, n21883,
    n21890, n21887, n39139, n37145, n39140, n39143, n21886, n26958, n38415,
    n26960, n39996, n40022, n21892, n21891, n21899, n21895, n38740, n40165,
    n21898, n21897, n40119, n21900, n21902, n38723, n21905, n40221, n40222,
    n21908, n37427, n21909, n21910, n40546, n21912, n34615, n40160, n21915,
    n21917, n35489, n21920, n35946, n21922, n40209, n21923, n21924, n40210,
    n21929, n21928, n35678, n29793, n21938, n21937, n21941, n21940, n21956,
    n21948, n21946, n21944, n21945, n21947, n21950, n21953, n21952, n21954,
    n21955, n21958, n21957, n21961, n21960, n21963, n21962, n21967, n21966,
    n21971, n21969, n21968, n21970, n25175, n21974, n21973, n21978, n21976,
    n21975, n21977, n35495, n21980, n21979, n21984, n21982, n21981, n21983,
    n34625, n21986, n21985, n21990, n21988, n21987, n21989, n35581, n21992,
    n21991, n21996, n21994, n21993, n21995, n34468, n21998, n21997, n22002,
    n22000, n21999, n22001, n33877, n22004, n22003, n22008, n22006, n22005,
    n22007, n26965, n22010, n22009, n22014, n22012, n22011, n22013, n32243,
    n22016, n22015, n22020, n22018, n22017, n22019, n25969, n22022, n22021,
    n22026, n22024, n22023, n22025, n33542, n22028, n37823, n22032, n22030,
    n22029, n22031, n22034, n22033, n34509, n22038, n22036, n22035, n22037,
    n22040, n22039, n33550, n22046, n22044, n22042, n22041, n22043, n22045,
    n32962, n40334, n22052, n22050, n22048, n22047, n22049, n22051, n33703,
    n22056, n22054, n22053, n22055, n22058, n22057, n34232, n22064, n22062,
    n22060, n22059, n22061, n22063, n34777, n22068, n22066, n22065, n22067,
    n22070, n22069, n36043, n22077, n22071, n22075, n22073, n22072, n22074,
    n22076, n35951, n22084, n22078, n22082, n22080, n22079, n22081, n22083,
    n35683, n22089, n22118, n34073, n25567, n27360, n27446, n27361, n27839,
    n22090, n27785, n22091, n27436, n30125, n22092, n22093, n22096, n22094,
    n22095, n22097, n22102, n22098, n22099, n22101, n22116, n22104, n22108,
    n22123, n22105, n22106, n22107, n22113, n22109, n22111, n22112, n25574,
    n22115, n22117, n22125, n22119, n22121, n22124, n22126, n30818, n22131,
    n22133, n39129, n25959, n25963, n22134, n39715, n26975, n40331, n22165,
    n22159, n34726, n33171, n22156, n22137, n22138, n22140, n22141, n22149,
    n22144, n22145, n30003, n22146, n22148, n25609, n22150, n22151, n22152,
    n33170, n33176, n22158, n22154, n25617, n30075, n33158, n33156, n22157,
    n40332, n40152, n34065, n22161, n40148, n33157, n22163, n22162, n22164,
    n25962, n22166, n40173, n22180, n25568, n22178, n30078, n30073, n22177,
    n22179, n40710, n22185, n22183, n22182, n22184, n25281, n22187, n22186,
    n22189, n22188, n35502, n22191, n22190, n22193, n22192, n34623, n22196,
    n22195, n22198, n22197, n35359, n22200, n22199, n22239, n22237, n22202,
    n22201, n22206, n22204, n22203, n22205, n22234, n22210, n22209, n22215,
    n22213, n36001, n22212, n22214, n22232, n22217, n22216, n22221, n22219,
    n22218, n22220, n22230, n26139, n22523, n22224, n22223, n22228, n22226,
    n22225, n22227, n22229, n22231, n22233, n34463, n22235, n22236, n22238,
    n33656, n22274, n22241, n22240, n22245, n22243, n22242, n22244, n22272,
    n22249, n22248, n22254, n22252, n36056, n22251, n22253, n22270, n22256,
    n22255, n22260, n22258, n22257, n22259, n22268, n22262, n22261, n22266,
    n22264, n22263, n22265, n22267, n22269, n22271, n33874, n22273, n22278,
    n22276, n22275, n22277, n32110, n22312, n22280, n22279, n22284, n22282,
    n22281, n22283, n22310, n37448, n22287, n39645, n22286, n22292, n22290,
    n36226, n22289, n22291, n22308, n22294, n22293, n22298, n22296, n22295,
    n22297, n22306, n22300, n22299, n22304, n22302, n22301, n22303, n22305,
    n22307, n22309, n33214, n22311, n22316, n22314, n22313, n22315, n26983,
    n22353, n22318, n22317, n22322, n22320, n22319, n22321, n22351, n22326,
    n22325, n22332, n22330, n22327, n22329, n22331, n22349, n22334, n22333,
    n22338, n22336, n22335, n22337, n22347, n22340, n22339, n22345, n22343,
    n22342, n22344, n22346, n22348, n22350, n32237, n22352, n22357, n22355,
    n22354, n22356, n30575, n22415, n22403, n30543, n22363, n22362, n22365,
    n22364, n22378, n22367, n27841, n22366, n22381, n22369, n22368, n30490,
    n22383, n22372, n30532, n22374, n22373, n22377, n22375, n22376, n30531,
    n30481, n22387, n22384, n22386, n22385, n22388, n31195, n22391, n27840,
    n22390, n22393, n22392, n31194, n22395, n22394, n22400, n22398, n22397,
    n22399, n22402, n22401, n33202, n27493, n22405, n22404, n22407, n22406,
    n35074, n22410, n22409, n27503, n22412, n22411, n22414, n22413, n35071,
    n37878, n22417, n22416, n22419, n22418, n25956, n22421, n30652, n38844,
    n22424, n22423, n22426, n22425, n30651, n30574, n31116, n22428, n22427,
    n22460, n22430, n22429, n22434, n22432, n22431, n22433, n22442, n22436,
    n22435, n22440, n22438, n22437, n22439, n22441, n22458, n22444, n22443,
    n22448, n22446, n22445, n22447, n22456, n22450, n22449, n22454, n22452,
    n22451, n22453, n22455, n22457, n25737, n22459, n22462, n22461, n31115,
    n22464, n22463, n22496, n22466, n22465, n22470, n22468, n22467, n22469,
    n22478, n22472, n22471, n22476, n22474, n22473, n22475, n22477, n22494,
    n22480, n22479, n22484, n22482, n22481, n22483, n22492, n22486, n22485,
    n22490, n22488, n22487, n22489, n22491, n22493, n25739, n22495, n22498,
    n22497, n31874, n22500, n22499, n22533, n22502, n22501, n22506, n22504,
    n22503, n22505, n22514, n22508, n22507, n22512, n22510, n22509, n22511,
    n22513, n22531, n22516, n22515, n22520, n22518, n22517, n22519, n22529,
    n22522, n22521, n22527, n22525, n22524, n22526, n22528, n22530, n25740,
    n22532, n22535, n22534, n33139, n22537, n22536, n22570, n22539, n22538,
    n22543, n22541, n22540, n22542, n22551, n22545, n22544, n22549, n22547,
    n22546, n22548, n22550, n22567, n22553, n22552, n22557, n22555, n22554,
    n22556, n22565, n22559, n22558, n22563, n22561, n22560, n22562, n22564,
    n22566, n25741, n22569, n22573, n22572, n33606, n37425, n22575, n22574,
    n22577, n22576, n35670, n22579, n22578, n22581, n22580, n25853, n22583,
    n22582, n22585, n22584, n35690, n25277, n25272, n25287, n25301, n25169,
    n25168, n25173, n25171, n25170, n25172, n37917, n25282, n25179, n25177,
    n25176, n25178, n25181, n25180, n38249, n25186, n25184, n25183, n25185,
    n25188, n25187, n38063, n25195, n25193, n25189, n25191, n25190, n25192,
    n25194, n25256, n25220, n25217, n25213, n25207, n25208, n39014, n25211,
    n25210, n25214, n38069, n25216, n40877, n25228, n40879, n25223, n25221,
    n38251, n25229, n40580, n25224, n25225, n40878, n25226, n40578, n25231,
    n40882, n40697, n40581, n25230, n25232, n25245, n25239, n25241, n39272,
    n25242, n25243, n25244, n25376, n25255, n25253, n25249, n25251, n25250,
    n25252, n25254, n25346, n25269, n25298, n40713, n25318, n25420, n25271,
    n25270, n25274, n25273, n25313, n25276, n25275, n25279, n25278, n37915,
    n40567, n25284, n25283, n25286, n25285, n26214, n40869, n25289, n25288,
    n25291, n25290, n38067, n27810, n25293, n25292, n25295, n25294, n25363,
    n25422, n25299, n25300, n40715, n40923, n25302, n25426, n25329, n25331,
    n25385, n25333, n39749, n25338, n25345, n25343, n25339, n25341, n25340,
    n25342, n25344, n25400, n25360, n25359, n25362, n25361, n25414, n25413,
    n25421, n25424, n25381, n25382, n25390, n25388, n25384, n25386, n39935,
    n25387, n25442, n25523, n25399, n25393, n25395, n25394, n25397, n25396,
    n25398, n25456, n25512, n27816, n25417, n25416, n25419, n25418, n25511,
    n25522, n25423, n25425, n25556, n25439, n27060, n25444, n25468, n25553,
    n25455, n25453, n25449, n25451, n25450, n25452, n25454, n25495, n25471,
    n25469, n25470, n25481, n25474, n25473, n25477, n25476, n39888, n25479,
    n25480, n25506, n25657, n25484, n25494, n25492, n25487, n25490, n25489,
    n25491, n25493, n25499, n25497, n25498, n37757, n25528, n25526, n25532,
    n25508, n25507, n25510, n25509, n25552, n25551, n25521, n25516, n25515,
    n25519, n25517, n25518, n25520, n39881, n25530, n25524, n25554, n25525,
    n25527, n25529, P2_U3015_Lock, n35860, input_0, input_1, AND_1,
    input_2, OR_2, input_3, OR_3, input_4, AND_4, input_5, OR_5, input_6,
    OR_6, input_7, AND_7, input_8, OR_8, input_9, AND_9, input_10, OR_10,
    input_11, OR_11, input_12, AND_12, input_13, AND_13, input_14, AND_14,
    input_15, AND_15, input_16, AND_16, input_17, AND_17, input_18, OR_18,
    input_19, AND_19, input_20, AND_20, input_21, AND_21, input_22, AND_22,
    input_23, OR_23, input_24, AND_24, input_25, OR_25, input_26, OR_26,
    input_27, AND_27, input_28, OR_28, input_29, OR_29, input_30, OR_30,
    input_31, AND_31, input_32, OR_32, input_33, AND_33, input_34, AND_34,
    input_35, OR_35, input_36, AND_36, input_37, AND_37, input_38, OR_38,
    input_39, OR_39, input_40, OR_40, input_41, OR_41, input_42, OR_42,
    input_43, OR_43, input_44, OR_44, input_45, OR_45, input_46, OR_46,
    input_47, OR_47, input_48, OR_48, input_49, AND_49, input_50, AND_50,
    input_51, AND_51, input_52, OR_52, input_53, OR_53, input_54, AND_54,
    input_55, OR_55, input_56, AND_56, input_57, OR_57, input_58, AND_58,
    input_59, AND_59, input_60, AND_60, input_61, AND_61, input_62, OR_62,
    input_63, AND_63, input_64, AND_64, input_65, OR_65, input_66, AND_66,
    input_67, AND_67, input_68, AND_68, input_69, AND_69, input_70, AND_70,
    input_71, OR_71, input_72, AND_72, input_73, OR_73, input_74, OR_74,
    input_75, AND_75, input_76, OR_76, input_77, AND_77, input_78, AND_78,
    input_79, AND_79, input_80, input_81, AND_81, input_82, OR_82,
    input_83, OR_83, input_84, AND_84, input_85, OR_85, input_86, OR_86,
    input_87, AND_87, input_88, OR_88, input_89, AND_89, input_90, OR_90,
    input_91, OR_91, input_92, AND_92, input_93, AND_93, input_94, AND_94,
    input_95, AND_95, input_96, AND_96, input_97, AND_97, input_98, OR_98,
    input_99, AND_99, input_100, AND_100, input_101, AND_101, input_102,
    AND_102, input_103, OR_103, input_104, AND_104, input_105, OR_105,
    input_106, OR_106, input_107, AND_107, input_108, OR_108, input_109,
    OR_109, input_110, OR_110, input_111, AND_111, input_112, OR_112,
    input_113, AND_113, input_114, AND_114, input_115, OR_115, input_116,
    AND_116, input_117, AND_117, input_118, OR_118, input_119, OR_119,
    input_120, OR_120, input_121, OR_121, input_122, OR_122, input_123,
    OR_123, input_124, OR_124, input_125, OR_125, input_126, OR_126,
    input_127, OR_127, input_128, OR_128, input_129, AND_129, input_130,
    AND_130, input_131, AND_131, input_132, OR_132, input_133, OR_133,
    input_134, AND_134, input_135, OR_135, input_136, AND_136, input_137,
    OR_137, input_138, AND_138, input_139, AND_139, input_140, AND_140,
    input_141, AND_141, input_142, OR_142, input_143, AND_143, input_144,
    AND_144, input_145, OR_145, input_146, AND_146, input_147, AND_147,
    input_148, AND_148, input_149, AND_149, input_150, AND_150, input_151,
    OR_151, input_152, AND_152, input_153, OR_153, input_154, OR_154,
    input_155, AND_155, input_156, OR_156, input_157, AND_157, input_158,
    AND_158, input_159, AND_159, AND_159_INV, CASOP;
  assign n34982 = ~n20827 & ~n20646;
  assign n21475 = n35590 | n21474;
  assign n40626 = ~n25564;
  assign n26095 = ~n26137;
  assign n20338 = ~n21147;
  assign n30005 = ~n27016 | ~n21414;
  assign n25608 = ~n21353 | ~n21330;
  assign n21353 = ~n21227 & ~n21779;
  assign n26187 = ~n20824 | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n21498 = n38451 | n21470;
  assign n25836 = ~n22285;
  assign n21791 = ~n21648;
  assign n25810 = ~n21544;
  assign n20333 = ~n20332;
  assign n22568 = n22235 | n21779;
  assign n34908 = ~n20337;
  assign n21369 = n22139 | n34783;
  assign n25478 = ~n21735 | ~n21734;
  assign n40860 = ~n25855;
  assign n20337 = ~n21779;
  assign n21268 = ~n21019;
  assign n21253 = ~n26187 & ~n34021;
  assign n26070 = ~n20353 | ~n34021;
  assign n40817 = ~n34001 | ~n26167;
  assign n34001 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n25616 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n20332 = ~n20952;
  assign n22371 = ~n40860 & ~P2_STATE2_REG_3__SCAN_IN;
  assign n35516 = ~n20981 & ~n20980;
  assign n25531 = n25530 & n20690;
  assign n40702 = ~n39539 | ~n20485;
  assign n39539 = ~n20619 | ~n21766;
  assign n36597 = ~n20582 | ~n21841;
  assign n34713 = n21836 ^ ~n34831;
  assign n21505 = n21504 & n21503;
  assign n35866 = ~n20827 & ~n20826;
  assign n21480 = n21476 & n21475;
  assign n20827 = ~n21459 | ~n21502;
  assign n21476 = n36849 | n21469;
  assign n21519 = n34839 | n21497;
  assign n20618 = n20798 & n20424;
  assign n20623 = n21461 | n21460;
  assign n35527 = ~n34064;
  assign n35075 = ~n20649 | ~n22403;
  assign n33203 = n20650 & n20423;
  assign n21471 = ~n21464 | ~n21463;
  assign n21464 = ~n21403 | ~n21402;
  assign n21458 = ~n21457 | ~n21456;
  assign n22379 = n22366 | n20648;
  assign n22155 = n21361 & n21360;
  assign n27051 = ~n29786;
  assign n21373 = n22103 | n21372;
  assign n21415 = n22181 | n21363;
  assign n21361 = n21354 | n21353;
  assign n21330 = ~n22153 & ~n25855;
  assign n22389 = ~n40626 | ~n37335;
  assign n22360 = n22370 & n21362;
  assign n21354 = n21362 & n34783;
  assign n22153 = ~n34783 | ~n35031;
  assign n22088 = ~n21164 & ~n21163;
  assign n35031 = n21298 | n21297;
  assign n22370 = n21779 | n34924;
  assign n21362 = ~n25855;
  assign n21265 = ~n21246 | ~n21245;
  assign n21327 = n21320 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n21320 = n21319 | n21318;
  assign n21170 = n21168 & n21167;
  assign n20339 = ~n21042;
  assign n26132 = ~n21148;
  assign n21212 = ~n21549;
  assign n21313 = ~n21312;
  assign n21549 = n26175 | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n22222 = n40820 & n34021;
  assign n26137 = n40469 | P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n21312 = ~n34008 & ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n40788 = ~n20923 | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n26169 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n34008 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n34021 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n33988 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n25782 = ~n40817 & ~n34021;
  assign n22328 = ~n21312 | ~n34021;
  assign n25822 = ~n21312 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n25513 = ~n25415;
  assign n21779 = ~n21226 & ~n21225;
  assign n20353 = ~n20933 & ~n25616;
  assign n20354 = ~n40626 | ~n37335;
  assign n21404 = ~n21384;
  assign n21666 = ~n21753;
  assign n21851 = n20790 ^ ~n21758;
  assign n21377 = ~n25693 & ~n25690;
  assign n20656 = ~n20377 | ~n20657;
  assign n20657 = ~n35071;
  assign n22181 = ~n21362 | ~n26203;
  assign n20512 = ~n21859 & ~n21852;
  assign n20507 = ~n21927 & ~n20508;
  assign n20508 = ~n20708 | ~n20509;
  assign n20509 = ~n21926;
  assign n20708 = ~n25220 & ~n20709;
  assign n20710 = n20364 | P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n20785 = ~n20786 & ~n20456;
  assign n20786 = ~n20361 & ~n20413;
  assign n34467 = ~n34233 | ~n34232;
  assign n38064 = ~n37917 & ~n37916;
  assign n21197 = n21019 | n21611;
  assign n21754 = ~n20782 | ~n20783;
  assign n20782 = n21737 & n22359;
  assign n21753 = ~n21665 | ~n21664;
  assign n20783 = ~n20877;
  assign n21496 = n21480 & n21479;
  assign n20824 = ~n20823 & ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n20823 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n20712 = n21774 & n21833;
  assign n22323 = ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n21384 = n31666 | n30492;
  assign n21407 = ~n21399 & ~n21398;
  assign n21399 = ~n22142 & ~n34075;
  assign n21300 = n26137 | n21299;
  assign n20997 = ~n20996 & ~n20995;
  assign n20585 = ~n20645 | ~n20791;
  assign n20791 = n21858 & n20406;
  assign n21762 = ~n20825 | ~n20389;
  assign n20825 = n25970 | n25965;
  assign n21860 = ~n20707 | ~n20706;
  assign n21755 = ~n20501 | ~n21752;
  assign n20501 = n20875 | n35084;
  assign n21836 = ~n20578 | ~n37025;
  assign n27052 = ~n22176;
  assign n20800 = n22027 ^ ~n20795;
  assign n20795 = ~n21450;
  assign n21225 = ~n21224 | ~n21223;
  assign n25218 = ~n20507;
  assign n25206 = ~n21927 & ~n21926;
  assign n21927 = n21921 | n21916;
  assign n21872 = n21888 | n21889;
  assign n20511 = ~n21885;
  assign n20967 = ~n20958 & ~n20957;
  assign n21444 = ~n20822 | ~n21430;
  assign n21965 = ~n29333 & ~n21384;
  assign n21438 = n25488 | n21436;
  assign n20648 = n20386 | n22367;
  assign n31666 = ~n29331 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n25485 = n22132 | n29336;
  assign n20787 = ~n20788 & ~n20442;
  assign n20554 = n20555 | n35581;
  assign n27013 = ~n22122 | ~n22121;
  assign n20688 = n21762 ^ ~n21763;
  assign n21520 = ~n21478 | ~n21477;
  assign n20624 = ~n20800 | ~n20799;
  assign n20799 = ~n21458;
  assign n21459 = ~n20801 | ~n21458;
  assign n20801 = ~n20800;
  assign n21164 = ~n21146 | ~n21145;
  assign n21194 = n21181 & n21180;
  assign n29331 = ~n35516;
  assign n29333 = ~n22175;
  assign n20660 = ~n22409;
  assign n20703 = ~n20704 | ~n25400;
  assign n37916 = ~n38250 | ~n38249;
  assign n20555 = ~n20556 | ~n34777;
  assign n20556 = ~n34468;
  assign n34233 = n32963 & n20467;
  assign n20550 = ~n33877;
  assign n20694 = ~n20695 & ~n25553;
  assign n20639 = ~n20641 | ~n20640;
  assign n20640 = ~n20904;
  assign n25379 = n25334 ^ ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n25334 = n39749 | n25440;
  assign n20638 = ~n20710 | ~n20396;
  assign n37331 = ~P2_STATE2_REG_2__SCAN_IN;
  assign n20692 = n25528 & n40719;
  assign n20691 = ~n25527 | ~n20450;
  assign n40719 = n22174 & n34035;
  assign n40931 = n22174 & n30086;
  assign n21695 = n21673 | n21672;
  assign n21623 = n21602 | n21601;
  assign n26175 = ~n33988 | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n20634 = ~n20636 & ~n20635;
  assign n20635 = ~n25379;
  assign n20636 = ~n20639 & ~n20637;
  assign n20637 = ~n20638;
  assign n20933 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n21497 = ~n38451 | ~n30599;
  assign n20923 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n40469 = ~n34001 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n21176 = ~n22222 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n21391 = ~n22360 | ~n21352;
  assign n21352 = n21351 & n21374;
  assign n21333 = n21057 & n21056;
  assign n21198 = n21196 & n21195;
  assign n21210 = ~n21209 & ~n21208;
  assign n21204 = n22328 | n21203;
  assign n21224 = ~n21218 & ~n21217;
  assign n21889 = n34908 & P2_EBX_REG_10__SCAN_IN;
  assign n21885 = n34908 & P2_EBX_REG_8__SCAN_IN;
  assign n20951 = ~n25799 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n21840 = n21823 | n21822;
  assign n21833 = n20438 & n20504;
  assign n20504 = n20505 | n34908;
  assign n26066 = ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n21395 = n22136 & P2_STATE2_REG_0__SCAN_IN;
  assign n26147 = ~n25822;
  assign n26100 = ~n26132;
  assign n25182 = ~n25488;
  assign n21913 = ~n21880 & ~n20713;
  assign n20713 = n20714 | n21907;
  assign n21857 = ~n21856 | ~n21855;
  assign n21856 = n21851 | n25478;
  assign n20584 = ~n34712;
  assign n21751 = ~n20876 | ~n21749;
  assign n20876 = ~n34716 | ~n34717;
  assign n21450 = n21449 & n21448;
  assign n20877 = ~n21562 | ~n21561;
  assign n21456 = n21455 & n21454;
  assign n21457 = n25448 | n34831;
  assign n21501 = ~n20689 | ~n20617;
  assign n20689 = ~n21498;
  assign n21512 = ~n21470 | ~n20796;
  assign n20705 = ~n22176 | ~n21936;
  assign n25332 = ~n25240 & ~n25239;
  assign n25240 = n25215 | n25207;
  assign n25215 = ~n25219 | ~n25213;
  assign n21921 = n21919 | n21918;
  assign n20714 = n20715 | n21901;
  assign n20715 = n20471 | n21879;
  assign n21896 = ~n21894 | ~n21893;
  assign n21894 = ~n21872 & ~n21871;
  assign n21888 = ~n20707 | ~n20394;
  assign n20707 = ~n21853;
  assign n21845 = ~n21840 & ~n21838;
  assign n20704 = n25346 & n25256;
  assign n21443 = n21434 & n21433;
  assign n21425 = ~n21423 | ~n21422;
  assign n21423 = n25488 | n21421;
  assign n20882 = ~n21413 | ~n34004;
  assign n25364 = ~n25312 & ~n25313;
  assign n25312 = ~n38068 | ~n38067;
  assign n25854 = ~n34623 & ~n34622;
  assign n33607 = ~n33656 & ~n33655;
  assign n21376 = ~n35031;
  assign n21303 = n26070 | n26136;
  assign n20872 = ~n26977 & ~n20873;
  assign n20873 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN | ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n21014 = ~n20998 | ~n20997;
  assign n25441 = n27060 | n25440;
  assign n20869 = ~n21768 & ~n20870;
  assign n20870 = ~n20872;
  assign n20697 = n25301 & P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n38068 = ~n37914 & ~n37915;
  assign n26215 = ~n25281 & ~n25280;
  assign n25280 = ~n35691 | ~n35690;
  assign n35684 = ~n35495 & ~n35494;
  assign n35691 = ~n35502 & ~n35501;
  assign n35501 = ~n25854 | ~n25853;
  assign n25167 = ~n25448;
  assign n34622 = ~n35671 | ~n35670;
  assign n20878 = n20879 & n21910;
  assign n40137 = n21909 ^ ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n35671 = ~n35359 & ~n35358;
  assign n35358 = ~n33607 | ~n33606;
  assign n33140 = ~n32109 & ~n32110;
  assign n32109 = ~n31875 | ~n31874;
  assign n31875 = ~n26982 & ~n26983;
  assign n22176 = ~n29331 | ~n40626;
  assign n20655 = n20656 & n25956;
  assign n21858 = n21857 | n25965;
  assign n25968 = ~n34510 | ~n34509;
  assign n25974 = n21857 ^ ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n20662 = ~n21779 | ~n37335;
  assign n21756 = ~n21755;
  assign n36596 = n21848 ^ ~n37823;
  assign n33541 = ~n20624 | ~n22028;
  assign n22420 = ~n22568;
  assign n20647 = ~n38451;
  assign n21245 = ~n21244 & ~n21243;
  assign n25475 = ~n20707 | ~n20512;
  assign n37920 = n25219 | n20510;
  assign n20510 = ~n20507 & ~n20506;
  assign n25222 = ~n25206 | ~n25205;
  assign n21879 = n34908 & P2_EBX_REG_14__SCAN_IN;
  assign n21878 = ~n21880 & ~n21879;
  assign n21880 = n21896 | n21863;
  assign n20981 = ~n20967 | ~n20966;
  assign n20701 = ~n20703 & ~n20702;
  assign n20702 = ~n25456;
  assign n38250 = ~n25175 & ~n25174;
  assign n34624 = ~n20552 | ~n20455;
  assign n20552 = ~n34467;
  assign n20553 = ~n20554;
  assign n32963 = ~n32243 & ~n32242;
  assign n33551 = ~n25969 & ~n25968;
  assign n34510 = ~n33542 & ~n33541;
  assign n21461 = n21444 ^ ~n21443;
  assign n21441 = n21440 & n21439;
  assign n21442 = n25448 | n21435;
  assign n25693 = n21375 | n21374;
  assign n35494 = ~n35952 | ~n35951;
  assign n20794 = ~n25529 | ~n25526;
  assign n20695 = ~n20697 | ~n20696;
  assign n20696 = ~n25424;
  assign n25238 = ~n20643 | ~n20378;
  assign n20643 = ~n40212 | ~n20785;
  assign n25237 = n25209 ^ ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n25209 = n39014 | n25440;
  assign n25174 = ~n35684 | ~n35683;
  assign n35952 = ~n34624 & ~n34625;
  assign n40118 = n38688 & n25478;
  assign n20690 = ~n20692 & ~n20691;
  assign n21247 = ~n26187 & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n21544 = ~n25794;
  assign n26048 = ~n26069;
  assign n20952 = ~n40817 & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n20359 = n20623 | n20387;
  assign n20360 = n40137 & n20881;
  assign n20361 = n20884 & n21925;
  assign n20363 = n22222 & P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n20364 = ~n39272 & ~n25329;
  assign n20788 = ~n21925;
  assign n21257 = ~n40788 & ~n34021;
  assign n20377 = n20659 & n22415;
  assign n20378 = n20513 & n25232;
  assign n20379 = n21193 & n21192;
  assign n20381 = n20512 & n20511;
  assign n20383 = ~n21877 & ~n40027;
  assign n21148 = ~n26175 & ~n34021;
  assign n20386 = n22371 & P2_EAX_REG_1__SCAN_IN;
  assign n20387 = n21458 ^ n21450;
  assign n20389 = n21760 | n21759;
  assign n20706 = ~n21852;
  assign n20394 = n20381 & n21866;
  assign n20396 = n20364 | n20711;
  assign n20398 = n25211 & n25210;
  assign n30599 = ~n21471 | ~n21467;
  assign n21004 = ~n21253;
  assign n22341 = ~n21004;
  assign n20402 = n25441 ^ P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n20406 = n20383 & n20483;
  assign n21842 = n21754 ^ ~n21753;
  assign n20413 = n20884 & n40210;
  assign n20414 = n20884 & n20787;
  assign n20415 = n21900 & n20360;
  assign n20416 = n21406 & n21413;
  assign n20418 = n21270 & n21269;
  assign n20423 = n22387 | n22388;
  assign n20424 = n21445 | n20387;
  assign n20426 = n21019 | n22324;
  assign n20427 = n21880 | n20715;
  assign n20428 = n20579 & n35090;
  assign n20430 = n20687 & n39136;
  assign n20432 = n21445 & n20387;
  assign n20438 = ~n34908 | ~n21772;
  assign n20442 = n40209 & n21923;
  assign n20443 = n32962 & n20551;
  assign n20444 = n20443 & n33703;
  assign n20447 = n25524 & n25554;
  assign n34004 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n20450 = ~n20447 & ~n20794;
  assign n21925 = ~n35489 & ~n25440;
  assign n20455 = n20553 & n36043;
  assign n22361 = ~n20505;
  assign n20505 = n21558 | n21559;
  assign n20456 = n20442 & n20788;
  assign n20460 = n21880 | n20714;
  assign n20467 = n20444 & n20550;
  assign n20468 = n20707 & n20381;
  assign n21972 = ~n21965;
  assign n20617 = ~n34839;
  assign n25440 = ~n25478;
  assign n20709 = ~n25205;
  assign n40929 = n22174 & n22133;
  assign n20471 = n34908 & P2_EBX_REG_15__SCAN_IN;
  assign n20483 = n35556 | n38853;
  assign n37335 = ~P2_STATE2_REG_3__SCAN_IN;
  assign n20485 = n20869 & P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n20831 = ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n25219 = ~n25218 & ~n25217;
  assign n20506 = ~n25217;
  assign n21919 = ~n21913 | ~n21911;
  assign n20513 = ~n20785 | ~n20414;
  assign n20551 = ~n26965;
  assign n20578 = ~n34716 | ~n25440;
  assign n34716 = n20877 ^ ~n21737;
  assign n21737 = ~n21596 | ~n21595;
  assign n20582 = ~n20580 | ~n20428;
  assign n20579 = ~n21837 | ~n20584;
  assign n20580 = ~n20581 | ~n21837;
  assign n20581 = ~n34713;
  assign n20644 = ~n20585 | ~n20415;
  assign n40212 = ~n20590 | ~n21915;
  assign n20590 = ~n40161 | ~n40160;
  assign n34839 = ~n20359 | ~n20618;
  assign n20619 = ~n20430 | ~n20620;
  assign n20620 = ~n20688 | ~n21764;
  assign n22027 = ~n20623 | ~n21445;
  assign n20798 = ~n20623 | ~n20432;
  assign n38451 = n21462 & n20623;
  assign n20646 = ~n20624 | ~n20647;
  assign n20826 = ~n38451 | ~n20624;
  assign n25257 = ~n38064 | ~n38063;
  assign n25383 = ~n20632 | ~n20634;
  assign n20632 = ~n25245 | ~n20638;
  assign n20641 = ~n20710;
  assign n40161 = n21914 ^ ~n40546;
  assign n21914 = ~n20644 | ~n20878;
  assign n20645 = ~n25973 | ~n25974;
  assign n22380 = ~n30480 & ~n30481;
  assign n30480 = n22379 ^ ~n22378;
  assign n37914 = ~n26215 | ~n26214;
  assign n26982 = ~n31116 | ~n31115;
  assign n20649 = ~n33203 | ~n33202;
  assign n20650 = n31195 | n31194;
  assign n20658 = ~n22410 | ~n20377;
  assign n22422 = ~n20658 | ~n20655;
  assign n20659 = ~n35071 | ~n20660;
  assign n25415 = n22181 | n20662;
  assign n20687 = ~n21764 | ~n38853;
  assign n20693 = ~n40702;
  assign n25501 = ~n20693 | ~n20694;
  assign n20700 = ~n25257;
  assign n25496 = ~n20700 | ~n20701;
  assign n21773 = ~n21054 | ~n20705;
  assign n21853 = ~n21845 | ~n21844;
  assign n20711 = ~n25244;
  assign n21823 = ~n21775 | ~n20712;
  assign n21832 = ~n21775 | ~n21774;
  assign n20784 = ~n20783 | ~n21737;
  assign n21750 = n20784 ^ ~n22359;
  assign n21761 = ~n20790 & ~n21704;
  assign n20790 = ~n21667 | ~n21666;
  assign n20822 = ~n21471 | ~n20797;
  assign n20796 = ~n20797;
  assign n21509 = ~n21470 | ~n20797;
  assign n34064 = n21472 ^ ~n20797;
  assign n20797 = n21424 ^ ~n21426;
  assign n21241 = ~n22222 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n21207 = ~n22222 | ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n21141 = ~n22222 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n21278 = ~n22222 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n20993 = ~n22222 | ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n20962 = ~n22222 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n26167 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n20875 = n21750 ^ ~n21751;
  assign n20879 = ~n20360 | ~n40222;
  assign n20881 = ~n40221 | ~n21906;
  assign n21446 = ~n21407 | ~n21406;
  assign n21418 = ~n20883 | ~n20882;
  assign n20883 = ~n20416 | ~n21407;
  assign n20884 = n25224 & n20398;
  assign n25443 = ~n25388 | ~n25387;
  assign n30816 = ~n26169 & ~n34004;
  assign n21226 = ~n21211 | ~n21210;
  assign n20890 = P2_STATE2_REG_0__SCAN_IN & P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n25486 = ~n21972;
  assign n22194 = ~n22371;
  assign n20896 = n21323 & n21322;
  assign n22571 = ~n22389;
  assign n20898 = n21309 & n21308;
  assign n20900 = n21306 & n21305;
  assign n20901 = n21325 & n21324;
  assign n20903 = n21566 & n21565;
  assign n21759 = ~n21851;
  assign n20904 = n25242 & n25478;
  assign n21147 = ~n21247;
  assign n21256 = ~n40788 & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n22285 = ~n25782;
  assign n25753 = ~n25799;
  assign n21206 = n25822 | n21615;
  assign n20984 = n21019 | n21474;
  assign n20985 = n20983 & n20982;
  assign n21357 = n21355 | n21779;
  assign n21234 = ~n25782 | ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n21231 = n21019 | n21230;
  assign n20910 = n21018 | n21017;
  assign n20960 = n25822 | n20959;
  assign n21454 = n21453 & n21452;
  assign n21274 = ~n20418 | ~n21271;
  assign n21057 = n21125 & n20914;
  assign n21871 = n34908 & P2_EBX_REG_11__SCAN_IN;
  assign n25488 = ~n21377 | ~n21404;
  assign n25565 = ~n31666;
  assign n21365 = ~n21376 | ~n35516;
  assign n21439 = n21438 & n21437;
  assign n21263 = ~n21252 & ~n21251;
  assign n25389 = ~n39935 & ~n25440;
  assign n21906 = ~n40222;
  assign n21766 = n21765 | n39141;
  assign n25514 = ~n22194;
  assign n21859 = n21821 & n21820;
  assign n40439 = n35678 | n25440;
  assign n33655 = ~n33140 | ~n33139;
  assign n25970 = n21760 ^ ~n21759;
  assign n21460 = ~n21442 | ~n21441;
  assign n22122 = ~n21963 | ~n21962;
  assign n22143 = ~n21368 | ~n22088;
  assign n25472 = n25385 | n25384;
  assign n36439 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n32242 = ~n33551 | ~n33550;
  assign n22174 = n22126 & n34083;
  assign n34075 = ~P2_STATE2_REG_0__SCAN_IN;
  assign n36540 = ~P2_STATE2_REG_2__SCAN_IN & ~P2_STATE2_REG_3__SCAN_IN;
  assign n41068 = ~n36540 | ~n21431;
  assign n40868 = P2_STATE2_REG_0__SCAN_IN | n41068;
  assign n40691 = ~n40868;
  assign n34028 = ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n21056 = ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~n34028;
  assign n21018 = P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n21017 = ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~n36439;
  assign n20909 = ~n35860 | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n21053 = ~n20910 | ~n20909;
  assign n21051 = P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n20913 = ~n21053 | ~n21051;
  assign n20911 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n20912 = ~n20911 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n21123 = ~n20913 | ~n20912;
  assign n21122 = P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n21125 = ~n21123 | ~n21122;
  assign n21447 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n20914 = ~n21447 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n20916 = ~n21056 & ~n21057;
  assign n34046 = ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n20915 = ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & ~n34046;
  assign n22120 = ~n20916 & ~n20915;
  assign n21019 = ~n30816 | ~n20933;
  assign n20918 = ~n21268 | ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n20917 = ~n20333 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n20922 = ~n20918 | ~n20917;
  assign n20920 = ~n26095 | ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n26069 = ~n22341;
  assign n20919 = ~n26048 | ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n20921 = ~n20920 | ~n20919;
  assign n20949 = ~n20922 & ~n20921;
  assign n20953 = ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n20928 = ~n21648 & ~n20953;
  assign n20924 = ~n26169;
  assign n25799 = n20924 & n34001;
  assign n20926 = ~n25827 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n25794 = ~n26169 & ~n34008;
  assign n35840 = ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n20925 = ~n25810 | ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n20927 = ~n20926 | ~n20925;
  assign n20930 = ~n20928 & ~n20927;
  assign n26127 = ~n22328;
  assign n20929 = ~n26127 | ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n20947 = ~n20930 | ~n20929;
  assign n20932 = ~n25836 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n20931 = ~n25783 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n20937 = ~n20932 | ~n20931;
  assign n26146 = ~n26070;
  assign n20935 = ~n26146 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n20934 = ~n26100 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n20936 = ~n20935 | ~n20934;
  assign n20945 = ~n20937 & ~n20936;
  assign n40820 = ~n25616 & ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n20939 = ~n22222 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n20938 = ~n20338 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n20943 = ~n20939 | ~n20938;
  assign n20941 = ~n26147 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n20940 = ~n25744 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n20942 = ~n20941 | ~n20940;
  assign n20944 = ~n20943 & ~n20942;
  assign n20946 = ~n20945 | ~n20944;
  assign n20948 = ~n20947 & ~n20946;
  assign n31893 = ~n20949 | ~n20948;
  assign n20950 = ~n25794 | ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n20958 = ~n20951 | ~n20950;
  assign n20955 = ~n20332 & ~n35840;
  assign n20954 = ~n22328 & ~n20953;
  assign n20956 = ~n20955 & ~n20954;
  assign n22324 = ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n20957 = ~n20956 | ~n20426;
  assign n20961 = ~n25782 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n20959 = ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n20965 = ~n20961 | ~n20960;
  assign n20963 = ~n26146 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n20964 = ~n20963 | ~n20962;
  assign n20966 = ~n20965 & ~n20964;
  assign n20969 = ~n21247 | ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n20968 = ~n21256 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n20973 = ~n20969 | ~n20968;
  assign n20971 = ~n22341 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n20970 = ~n21212 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n20972 = ~n20971 | ~n20970;
  assign n20979 = ~n20973 & ~n20972;
  assign n20975 = ~n21148 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n20974 = ~n20339 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n20977 = ~n20975 | ~n20974;
  assign n20976 = ~n26137 & ~n22323;
  assign n20978 = ~n20977 & ~n20976;
  assign n20980 = ~n20979 | ~n20978;
  assign n20983 = ~n25799 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n20982 = ~n25794 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n21474 = ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n20990 = ~n20985 | ~n20984;
  assign n20988 = ~n25782 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n20986 = ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n20987 = n26070 | n20986;
  assign n20989 = ~n20988 | ~n20987;
  assign n20998 = ~n20990 & ~n20989;
  assign n20992 = ~n20952 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n39604 = ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n20991 = n22328 | n39604;
  assign n20996 = ~n20992 | ~n20991;
  assign n21469 = ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n20994 = n25822 | n21469;
  assign n20995 = ~n20994 | ~n20993;
  assign n21000 = ~n21247 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n20999 = ~n21321 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n21003 = ~n21000 | ~n20999;
  assign n21001 = ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n21002 = ~n26137 & ~n21001;
  assign n21012 = ~n21003 & ~n21002;
  assign n21006 = ~n22341 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n21005 = ~n21212 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n21010 = ~n21006 | ~n21005;
  assign n21008 = ~n21256 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n21007 = ~n20339 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n21009 = ~n21008 | ~n21007;
  assign n21011 = ~n21010 & ~n21009;
  assign n21013 = ~n21012 | ~n21011;
  assign n25564 = ~n21014 & ~n21013;
  assign n21016 = ~n31893 | ~n27052;
  assign n21943 = P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ^ ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n21015 = ~n22176 | ~n21943;
  assign n21827 = ~n21016 | ~n21015;
  assign n21942 = n21018 ^ ~n21017;
  assign n21949 = ~n22176 | ~n21942;
  assign n21055 = ~n21827 | ~n21949;
  assign n21021 = ~n21268 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n21020 = ~n21791 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n21025 = ~n21021 | ~n21020;
  assign n21023 = ~n26127 | ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n21022 = ~n20333 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n21024 = ~n21023 | ~n21022;
  assign n21033 = ~n21025 & ~n21024;
  assign n21027 = ~n25827 | ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n21026 = ~n25810 | ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n21031 = ~n21027 | ~n21026;
  assign n21029 = ~n26146 | ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n21028 = ~n26147 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n21030 = ~n21029 | ~n21028;
  assign n21032 = ~n21031 & ~n21030;
  assign n21050 = n21033 & n21032;
  assign n21035 = ~n26095 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n21034 = ~n22222 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n21039 = ~n21035 | ~n21034;
  assign n21037 = ~n20338 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n21036 = ~n25836 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n21038 = ~n21037 | ~n21036;
  assign n21048 = ~n21039 & ~n21038;
  assign n21041 = ~n26100 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n25744 = ~n21549;
  assign n21040 = ~n25744 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n21046 = ~n21041 | ~n21040;
  assign n21044 = ~n26048 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n21042 = ~n21257;
  assign n21535 = ~n20339;
  assign n21043 = ~n25783 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n21045 = ~n21044 | ~n21043;
  assign n21047 = ~n21046 & ~n21045;
  assign n21049 = n21048 & n21047;
  assign n21745 = ~n21050 | ~n21049;
  assign n21054 = n21745 | n22176;
  assign n21052 = ~n21051;
  assign n21951 = n21053 ^ ~n21052;
  assign n21936 = ~n21951;
  assign n21128 = ~n21055 | ~n21773;
  assign n21091 = ~n21333 | ~n22176;
  assign n21059 = ~n20338 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n21058 = ~n26048 | ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n21063 = ~n21059 | ~n21058;
  assign n21061 = ~n25744 | ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n21060 = ~n26100 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n21062 = ~n21061 | ~n21060;
  assign n21069 = ~n21063 & ~n21062;
  assign n25783 = ~n21535;
  assign n21065 = ~n25783 | ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n21648 = ~n21256;
  assign n21064 = ~n21791 | ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n21067 = ~n21065 | ~n21064;
  assign n40482 = ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n21066 = ~n26139 & ~n40482;
  assign n21068 = ~n21067 & ~n21066;
  assign n21089 = ~n21069 | ~n21068;
  assign n21071 = ~n20333 | ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n40468 = ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n21070 = n26070 | n40468;
  assign n21077 = n21071 & n21070;
  assign n22211 = ~n21268;
  assign n22246 = ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n21075 = ~n22211 & ~n22246;
  assign n21073 = ~n25799 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n21072 = ~n25794 | ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n21074 = ~n21073 | ~n21072;
  assign n21076 = ~n21075 & ~n21074;
  assign n21087 = ~n21077 | ~n21076;
  assign n21079 = ~n25782 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n21152 = ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n21078 = n22328 | n21152;
  assign n21085 = n21079 & n21078;
  assign n21080 = ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n21083 = ~n26137 & ~n21080;
  assign n21081 = ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n21082 = ~n25822 & ~n21081;
  assign n21084 = ~n21083 & ~n21082;
  assign n21086 = ~n21085 | ~n21084;
  assign n21088 = n21087 | n21086;
  assign n21736 = ~n21089 & ~n21088;
  assign n21090 = ~n27052 | ~n21736;
  assign n21780 = ~n21091 | ~n21090;
  assign n21093 = ~n26146 | ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n21092 = ~n26100 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n21097 = ~n21093 | ~n21092;
  assign n21095 = ~n26147 | ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n21094 = ~n25782 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n21096 = ~n21095 | ~n21094;
  assign n21105 = ~n21097 & ~n21096;
  assign n21099 = ~n22222 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n21098 = ~n20338 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n21103 = ~n21099 | ~n21098;
  assign n21101 = ~n26048 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n21100 = ~n25744 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n21102 = ~n21101 | ~n21100;
  assign n21104 = ~n21103 & ~n21102;
  assign n21121 = ~n21105 | ~n21104;
  assign n21107 = ~n26127 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n21106 = ~n25810 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n21111 = ~n21107 | ~n21106;
  assign n21109 = ~n21268 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n21108 = ~n21791 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n21110 = ~n21109 | ~n21108;
  assign n21119 = ~n21111 & ~n21110;
  assign n21113 = ~n20333 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n21112 = ~n25799 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n21117 = ~n21113 | ~n21112;
  assign n21115 = ~n26095 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n21114 = ~n25783 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n21116 = ~n21115 | ~n21114;
  assign n21118 = ~n21117 & ~n21116;
  assign n21120 = ~n21119 | ~n21118;
  assign n22396 = ~n21121 & ~n21120;
  assign n21127 = ~n22396 | ~n27052;
  assign n21124 = n21123 | n21122;
  assign n21332 = ~n21125 | ~n21124;
  assign n21126 = ~n22176 | ~n21332;
  assign n21776 = ~n21127 | ~n21126;
  assign n21939 = ~n21780 & ~n21776;
  assign n21129 = ~n21128 | ~n21939;
  assign n30072 = ~n22120 | ~n21129;
  assign n21331 = ~n30072;
  assign n21131 = ~n25799 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n21130 = ~n25794 | ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n21133 = n21131 & n21130;
  assign n22247 = ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n21132 = n21019 | n22247;
  assign n21137 = ~n21133 | ~n21132;
  assign n21135 = ~n21233 | ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n21134 = ~n25782 | ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n21136 = ~n21135 | ~n21134;
  assign n21146 = ~n21137 & ~n21136;
  assign n21140 = ~n20952 | ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n21138 = ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n21139 = n22328 | n21138;
  assign n21144 = ~n21140 | ~n21139;
  assign n22250 = ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n21142 = n25822 | n22250;
  assign n21143 = ~n21142 | ~n21141;
  assign n21145 = ~n21144 & ~n21143;
  assign n21151 = ~n21247 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n21149 = ~n21148;
  assign n21321 = ~n21149;
  assign n21150 = ~n21321 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n21154 = ~n21151 | ~n21150;
  assign n21153 = ~n26137 & ~n21152;
  assign n21162 = ~n21154 & ~n21153;
  assign n21156 = ~n22341 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n21155 = ~n21212 | ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n21160 = ~n21156 | ~n21155;
  assign n21158 = ~n21256 | ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n21157 = ~n20339 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n21159 = ~n21158 | ~n21157;
  assign n21161 = ~n21160 & ~n21159;
  assign n21163 = ~n21162 | ~n21161;
  assign n21166 = ~n25799 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n21165 = ~n25794 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n21168 = n21166 & n21165;
  assign n21674 = ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n21167 = n21019 | n21674;
  assign n21169 = ~n25782 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n21173 = ~n21170 | ~n21169;
  assign n21171 = ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n21172 = ~n26070 & ~n21171;
  assign n21181 = ~n21173 & ~n21172;
  assign n21175 = ~n20952 | ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n21792 = ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n21174 = n22328 | n21792;
  assign n21179 = ~n21175 | ~n21174;
  assign n22207 = ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n21177 = n25822 | n22207;
  assign n40787 = ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n21178 = ~n21177 | ~n21176;
  assign n21180 = ~n21179 & ~n21178;
  assign n21183 = ~n21247 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n21182 = ~n21321 | ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n21185 = ~n21183 | ~n21182;
  assign n22208 = ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n21184 = ~n26137 & ~n22208;
  assign n21193 = ~n21185 & ~n21184;
  assign n21187 = ~n21253 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n21186 = ~n21212 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n21191 = ~n21187 | ~n21186;
  assign n21189 = ~n21256 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n21188 = ~n20339 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n21190 = ~n21189 | ~n21188;
  assign n21192 = ~n21191 & ~n21190;
  assign n34924 = ~n21194 | ~n20379;
  assign n21227 = ~n22088 | ~n34924;
  assign n21196 = ~n25799 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n21195 = ~n25794 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n21611 = ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n21202 = ~n21198 | ~n21197;
  assign n21200 = ~n21233 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n21199 = ~n20952 | ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n21201 = ~n21200 | ~n21199;
  assign n21211 = ~n21202 & ~n21201;
  assign n21205 = ~n25782 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n21203 = ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n21209 = ~n21205 | ~n21204;
  assign n21615 = ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n21208 = ~n21207 | ~n21206;
  assign n21214 = ~n21253 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n21213 = ~n21212 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n21218 = ~n21214 | ~n21213;
  assign n21216 = ~n21247 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n21215 = ~n20339 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n21217 = ~n21216 | ~n21215;
  assign n21220 = ~n21321 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n21219 = ~n21256 | ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n21222 = ~n21220 | ~n21219;
  assign n21221 = ~n26137 & ~n26066;
  assign n21223 = ~n21222 & ~n21221;
  assign n21229 = ~n25799 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n21228 = ~n25794 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n21232 = n21229 & n21228;
  assign n21230 = ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n21237 = ~n21232 | ~n21231;
  assign n21233 = ~n26070;
  assign n21235 = ~n21233 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n21236 = ~n21235 | ~n21234;
  assign n21246 = ~n21237 & ~n21236;
  assign n21239 = ~n20952 | ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n22288 = ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n21238 = n22328 | n22288;
  assign n21244 = ~n21239 | ~n21238;
  assign n21240 = ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n21242 = n25822 | n21240;
  assign n21243 = ~n21242 | ~n21241;
  assign n21249 = ~n21247 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n21248 = ~n21321 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n21252 = ~n21249 | ~n21248;
  assign n21250 = ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n21251 = ~n26137 & ~n21250;
  assign n21255 = ~n21253 | ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n21254 = ~n21212 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n21261 = ~n21255 | ~n21254;
  assign n21259 = ~n21256 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n21258 = ~n21257 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n21260 = ~n21259 | ~n21258;
  assign n21262 = ~n21261 & ~n21260;
  assign n21264 = ~n21263 | ~n21262;
  assign n34783 = ~n21265 & ~n21264;
  assign n21267 = ~n25799 | ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n21266 = ~n25794 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n21270 = n21267 & n21266;
  assign n25821 = ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n21269 = n21019 | n25821;
  assign n21271 = ~n25782 | ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n21272 = ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n21273 = ~n26070 & ~n21272;
  assign n21283 = ~n21274 & ~n21273;
  assign n21277 = ~n20952 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n21275 = ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n21276 = n22328 | n21275;
  assign n21281 = ~n21277 | ~n21276;
  assign n21580 = ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n21279 = n25822 | n21580;
  assign n21280 = ~n21279 | ~n21278;
  assign n21282 = ~n21281 & ~n21280;
  assign n21298 = ~n21283 | ~n21282;
  assign n21285 = ~n21247 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n21284 = ~n21321 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n21288 = ~n21285 | ~n21284;
  assign n21286 = ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n21287 = ~n26137 & ~n21286;
  assign n21296 = ~n21288 & ~n21287;
  assign n21290 = ~n21253 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n21289 = ~n21212 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n21294 = ~n21290 | ~n21289;
  assign n21292 = ~n21256 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n21291 = ~n20339 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n21293 = ~n21292 | ~n21291;
  assign n21295 = ~n21294 & ~n21293;
  assign n21297 = ~n21296 | ~n21295;
  assign n21301 = ~n25782 | ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n21299 = ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n21302 = ~n21301 | ~n21300;
  assign n21304 = ~n21302 & ~n20363;
  assign n26136 = ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n21311 = ~n21304 | ~n21303;
  assign n21306 = ~n21247 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n21305 = ~n20339 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n21309 = ~n20952 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n21307 = ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n21308 = n22328 | n21307;
  assign n21310 = ~n20900 | ~n20898;
  assign n21329 = ~n21311 & ~n21310;
  assign n40816 = ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n21315 = n40469 | n40816;
  assign n40839 = ~n21313;
  assign n21314 = ~n40839 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n21319 = ~n21315 | ~n21314;
  assign n40838 = ~n26187;
  assign n21317 = ~n40838 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n21316 = ~n40820 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n21318 = ~n21317 | ~n21316;
  assign n21323 = ~n21321 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n21322 = ~n25794 | ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n21325 = ~n21212 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n21324 = ~n21256 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n21326 = ~n20896 | ~n20901;
  assign n21328 = ~n21327 & ~n21326;
  assign n25855 = n21329 & n21328;
  assign n30492 = ~n21934;
  assign n29786 = ~n30492 | ~n29331;
  assign n34035 = ~n25608 & ~n29786;
  assign n22114 = ~n21331 | ~n34035;
  assign n21959 = ~n21333 & ~n21332;
  assign n21335 = ~n21951 | ~n21959;
  assign n21334 = ~n21335;
  assign n21338 = ~n21943 | ~n21334;
  assign n21337 = ~n21942 & ~n21335;
  assign n21336 = ~n22120;
  assign n29821 = ~n21337 & ~n21336;
  assign n21339 = ~n21338 | ~n29821;
  assign n21343 = ~n21431 | ~n21339;
  assign n21340 = ~n26169 & ~n34001;
  assign n21341 = ~n21340 & ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n30489 = ~P2_FLUSH_REG_SCAN_IN & ~n21341;
  assign n21342 = ~P2_STATE2_REG_1__SCAN_IN | ~n30489;
  assign n22100 = ~n21343 | ~n21342;
  assign n30086 = ~n25608 & ~n22176;
  assign n34609 = ~P2_STATE2_REG_1__SCAN_IN & ~n37331;
  assign n29819 = ~P2_STATE2_REG_0__SCAN_IN | ~n34609;
  assign n34083 = ~n29819;
  assign n40434 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n40368 = ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n40109 = ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n21390 = ~n25608 | ~n34783;
  assign n21351 = n22088 & n35031;
  assign n21374 = ~n21779 | ~n34924;
  assign n22175 = ~n21390 & ~n21391;
  assign n33974 = ~n22175 | ~n27051;
  assign n21355 = ~n34924;
  assign n21356 = ~n21355 | ~n22088;
  assign n21359 = ~n21357 | ~n21356;
  assign n21358 = n25855 | n34783;
  assign n21360 = ~n21359 | ~n21358;
  assign n21934 = ~n25564;
  assign n26203 = ~n21934;
  assign n21363 = ~n21779 | ~n34783;
  assign n21364 = ~n21415 & ~n21365;
  assign n25610 = ~n22155 | ~n21364;
  assign n22132 = ~n33974 | ~n25610;
  assign n21366 = ~n21365;
  assign n22139 = ~n21366 | ~n34924;
  assign n21367 = n25855 | n21779;
  assign n21368 = ~n21367 | ~n35516;
  assign n29336 = ~n21369 & ~n22143;
  assign n25448 = ~n25485 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n21370 = ~n25448;
  assign n21403 = ~n21370 | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n25847 = ~n22370;
  assign n21371 = ~n25847 | ~n22088;
  assign n22103 = ~n21371 | ~n21374;
  assign n35016 = ~n22088;
  assign n22110 = ~n22370 | ~n35016;
  assign n21372 = ~n22110 | ~n40860;
  assign n22147 = ~n21373 | ~n35031;
  assign n21375 = ~n22088 | ~n25855;
  assign n22135 = ~n25693 | ~n21376;
  assign n21405 = ~n22147 | ~n22135;
  assign n22136 = ~n22370 | ~n25564;
  assign n21383 = ~n21405 | ~n21395;
  assign n25690 = ~n21376 | ~n34783;
  assign n21378 = ~P2_EBX_REG_0__SCAN_IN;
  assign n21381 = ~n25488 & ~n21378;
  assign n21431 = ~P2_STATE2_REG_1__SCAN_IN;
  assign n34078 = ~n34075 | ~n21431;
  assign n21379 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n21380 = ~n34078 | ~n21379;
  assign n21382 = ~n21381 & ~n21380;
  assign n21386 = n21383 & n21382;
  assign n21385 = ~n21965 | ~P2_REIP_REG_0__SCAN_IN;
  assign n21401 = ~n21386 | ~n21385;
  assign n21387 = ~n22370 | ~n35031;
  assign n21389 = ~n22155 | ~n21387;
  assign n25691 = ~n35516 | ~n25564;
  assign n21388 = ~n25691;
  assign n22142 = ~n21389 | ~n21388;
  assign n21393 = ~n21390;
  assign n21392 = ~n21391 | ~n25564;
  assign n21394 = ~n21393 | ~n21392;
  assign n21397 = ~n21394 | ~n25565;
  assign n21396 = ~n21395 | ~n35516;
  assign n21398 = ~n21397 | ~n21396;
  assign n21400 = ~n21407;
  assign n21402 = ~n21401 & ~n21400;
  assign n21406 = ~n21405 | ~n21404;
  assign n21412 = ~n21446 | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n25583 = ~n34924 & ~n34075;
  assign n30495 = ~n25583;
  assign n21410 = ~n25610 & ~n30495;
  assign n21408 = n34078 | n36439;
  assign n21409 = ~n25488 | ~n21408;
  assign n21411 = ~n21410 & ~n21409;
  assign n21463 = ~n21412 | ~n21411;
  assign n21413 = n34078 | n35860;
  assign n27016 = ~n22175 | ~n29331;
  assign n21414 = ~n29336;
  assign n21416 = ~n21415 & ~n22139;
  assign n34005 = n30005 | n21416;
  assign n21417 = ~n34005 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n21426 = ~n21418 | ~n21417;
  assign n21420 = ~n25485 | ~n20890;
  assign n21419 = ~n21965 | ~P2_REIP_REG_1__SCAN_IN;
  assign n21427 = ~n21420 | ~n21419;
  assign n21421 = ~P2_EBX_REG_1__SCAN_IN;
  assign n21422 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n21424 = ~n21427 & ~n21425;
  assign n21429 = ~n21426 & ~n21425;
  assign n21428 = ~n21427;
  assign n21430 = ~n21429 | ~n21428;
  assign n21434 = ~n21446 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n21432 = ~n34075 | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n21433 = n21432 & n21431;
  assign n21435 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n21440 = ~n21965 | ~P2_REIP_REG_2__SCAN_IN;
  assign n21436 = ~P2_EBX_REG_2__SCAN_IN;
  assign n21437 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n21445 = ~n21444 | ~n21443;
  assign n21449 = ~n21446 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n21448 = n34078 | n21447;
  assign n34831 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n21455 = ~n21965 | ~P2_REIP_REG_3__SCAN_IN;
  assign n21451 = ~P2_EBX_REG_3__SCAN_IN;
  assign n21453 = n25488 | n21451;
  assign n21452 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n21462 = ~n21461 | ~n21460;
  assign n21466 = ~n21463;
  assign n21465 = ~n21464;
  assign n21467 = ~n21466 | ~n21465;
  assign n21468 = ~n20647 & ~n21509;
  assign n36849 = ~n34839 | ~n21468;
  assign n21470 = ~n30599;
  assign n21472 = ~n21471;
  assign n21473 = ~n21498 & ~n34064;
  assign n35590 = ~n34839 | ~n21473;
  assign n21478 = ~n34839;
  assign n21477 = ~n21512;
  assign n35376 = ~n21520 & ~n38451;
  assign n21479 = ~n35376 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n21481 = n20647 & n21477;
  assign n34862 = ~n34839 | ~n21481;
  assign n21482 = ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n21486 = n34862 | n21482;
  assign n21483 = ~n21497 & ~n34064;
  assign n36500 = ~n34839 | ~n21483;
  assign n21484 = ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n21485 = n36500 | n21484;
  assign n21494 = ~n21486 | ~n21485;
  assign n21487 = ~n21498 & ~n35527;
  assign n36170 = ~n34839 | ~n21487;
  assign n21488 = ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n21492 = n36170 | n21488;
  assign n21489 = ~n21497 & ~n35527;
  assign n36075 = ~n34839 | ~n21489;
  assign n21490 = ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n21491 = n36075 | n21490;
  assign n21493 = ~n21492 | ~n21491;
  assign n21495 = ~n21494 & ~n21493;
  assign n21508 = ~n21496 | ~n21495;
  assign n36457 = ~n21519 & ~n34064;
  assign n21500 = ~n36457 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n37332 = ~n21501 & ~n34064;
  assign n21499 = ~n37332 | ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n21506 = n21500 & n21499;
  assign n36552 = ~n21501 & ~n35527;
  assign n21504 = ~n36552 | ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n21502 = ~n21509;
  assign n21503 = ~n35866 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n21507 = ~n21506 | ~n21505;
  assign n21526 = ~n21508 & ~n21507;
  assign n21510 = n20647 & n21502;
  assign n37718 = ~n34839 | ~n21510;
  assign n39591 = ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n21511 = n37718 | n39591;
  assign n21516 = ~n21511 | ~n40626;
  assign n21513 = ~n20647 & ~n21512;
  assign n35265 = ~n34839 | ~n21513;
  assign n21514 = ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n21515 = ~n35265 & ~n21514;
  assign n21518 = ~n21516 & ~n21515;
  assign n21517 = ~n34982 | ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n21524 = ~n21518 | ~n21517;
  assign n35843 = ~n21519 & ~n35527;
  assign n21522 = ~n35843 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n34805 = ~n21520 & ~n20647;
  assign n21521 = ~n34805 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n21523 = ~n21522 | ~n21521;
  assign n21525 = ~n21524 & ~n21523;
  assign n21562 = ~n21526 | ~n21525;
  assign n21528 = ~n20338 | ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n21527 = ~n26100 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n21532 = ~n21528 | ~n21527;
  assign n21530 = ~n22222 | ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n21529 = ~n26048 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n21531 = ~n21530 | ~n21529;
  assign n21541 = ~n21532 & ~n21531;
  assign n21534 = ~n26146 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n21533 = ~n25836 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n21539 = ~n21534 | ~n21533;
  assign n21537 = ~n26147 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n21536 = ~n25783 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n21538 = ~n21537 | ~n21536;
  assign n21540 = ~n21539 & ~n21538;
  assign n21559 = ~n21541 | ~n21540;
  assign n21543 = ~n26127 | ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n21542 = ~n21791 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n21548 = ~n21543 | ~n21542;
  assign n21546 = ~n20333 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n21545 = ~n25810 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n21547 = ~n21546 | ~n21545;
  assign n21557 = ~n21548 & ~n21547;
  assign n21551 = ~n21268 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n21550 = ~n25744 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n21555 = ~n21551 | ~n21550;
  assign n21553 = ~n26095 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n25827 = ~n25753;
  assign n21552 = ~n25827 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n21554 = ~n21553 | ~n21552;
  assign n21556 = ~n21555 & ~n21554;
  assign n21558 = ~n21557 | ~n21556;
  assign n21560 = ~n31893 | ~n30492;
  assign n21743 = n22361 | n21560;
  assign n22382 = ~n21745;
  assign n21561 = ~n21743 | ~n22382;
  assign n21564 = ~n37332 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n21563 = ~n35866 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n21567 = n21564 & n21563;
  assign n21566 = ~n35376 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n21565 = ~n34805 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n21588 = ~n21567 | ~n20903;
  assign n21570 = n35590 | n25821;
  assign n21568 = ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n21569 = n37718 | n21568;
  assign n21575 = ~n21570 | ~n21569;
  assign n21571 = ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n21573 = n36500 | n21571;
  assign n25818 = ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n21572 = n34862 | n25818;
  assign n21574 = ~n21573 | ~n21572;
  assign n21586 = ~n21575 & ~n21574;
  assign n21576 = ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n21579 = n35265 | n21576;
  assign n21577 = ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n21578 = n36170 | n21577;
  assign n21584 = ~n21579 | ~n21578;
  assign n25817 = ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n21582 = n36075 | n25817;
  assign n21581 = n36849 | n21580;
  assign n21583 = ~n21582 | ~n21581;
  assign n21585 = ~n21584 & ~n21583;
  assign n21587 = ~n21586 | ~n21585;
  assign n21596 = ~n21588 & ~n21587;
  assign n21590 = ~n34982 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n21589 = ~n35843 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n21594 = ~n21590 | ~n21589;
  assign n21592 = ~n36457 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n21591 = ~n36552 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n21593 = ~n21592 | ~n21591;
  assign n21595 = ~n21594 & ~n21593;
  assign n22359 = ~n21736;
  assign n21667 = ~n21754;
  assign n21598 = ~n34982 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n21597 = ~n35376 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n21602 = ~n21598 | ~n21597;
  assign n21600 = ~n36552 | ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n21599 = ~n34805 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n21601 = ~n21600 | ~n21599;
  assign n21603 = ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n21605 = n35265 | n21603;
  assign n40631 = ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n21604 = n36500 | n40631;
  assign n21610 = ~n21605 | ~n21604;
  assign n21606 = ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n21608 = n34862 | n21606;
  assign n21651 = ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n21607 = n37718 | n21651;
  assign n21609 = ~n21608 | ~n21607;
  assign n21621 = ~n21610 & ~n21609;
  assign n26065 = ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n21613 = n36170 | n26065;
  assign n21612 = n35590 | n21611;
  assign n21619 = ~n21613 | ~n21612;
  assign n21614 = ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n21617 = n36075 | n21614;
  assign n21616 = n36849 | n21615;
  assign n21618 = ~n21617 | ~n21616;
  assign n21620 = ~n21619 & ~n21618;
  assign n21622 = ~n21621 | ~n21620;
  assign n21631 = ~n21623 & ~n21622;
  assign n21625 = ~n35843 | ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n21624 = ~n36457 | ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n21629 = ~n21625 | ~n21624;
  assign n21627 = ~n37332 | ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n21626 = ~n35866 | ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n21628 = ~n21627 | ~n21626;
  assign n21630 = ~n21629 & ~n21628;
  assign n21665 = ~n21631 | ~n21630;
  assign n21633 = ~n26147 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n21632 = ~n25836 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n21637 = ~n21633 | ~n21632;
  assign n21635 = ~n26095 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n21634 = ~n22523 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n21636 = ~n21635 | ~n21634;
  assign n21645 = ~n21637 & ~n21636;
  assign n21639 = ~n26048 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n21638 = ~n25783 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n21643 = ~n21639 | ~n21638;
  assign n21641 = ~n26146 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n21640 = ~n20338 | ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n21642 = ~n21641 | ~n21640;
  assign n21644 = ~n21643 & ~n21642;
  assign n21663 = n21645 & n21644;
  assign n21647 = ~n25827 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n21646 = ~n25810 | ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n21650 = n21647 & n21646;
  assign n21649 = ~n21791 | ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n21655 = ~n21650 | ~n21649;
  assign n21653 = n22211 | n21651;
  assign n21652 = n22328 | n26066;
  assign n21654 = ~n21653 | ~n21652;
  assign n21661 = ~n21655 & ~n21654;
  assign n21657 = ~n26100 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n21656 = ~n25744 | ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n21659 = ~n21657 | ~n21656;
  assign n21658 = n20333 & P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n21660 = ~n21659 & ~n21658;
  assign n21662 = n21661 & n21660;
  assign n22408 = ~n21663 | ~n21662;
  assign n21664 = n22408 | n40626;
  assign n21669 = ~n35843 | ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n21668 = ~n34805 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n21673 = ~n21669 | ~n21668;
  assign n21671 = ~n34982 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n21670 = ~n36552 | ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n21672 = ~n21671 | ~n21670;
  assign n21676 = n35590 | n21674;
  assign n21675 = n36849 | n22207;
  assign n21682 = ~n21676 | ~n21675;
  assign n21677 = ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n21680 = n36075 | n21677;
  assign n21678 = ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n21679 = n34862 | n21678;
  assign n21681 = ~n21680 | ~n21679;
  assign n21693 = ~n21682 & ~n21681;
  assign n21683 = ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n21686 = n37718 | n21683;
  assign n21684 = ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n21685 = n36500 | n21684;
  assign n21691 = ~n21686 | ~n21685;
  assign n21687 = ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n21689 = n35265 | n21687;
  assign n40773 = ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n21688 = n36170 | n40773;
  assign n21690 = ~n21689 | ~n21688;
  assign n21692 = ~n21691 & ~n21690;
  assign n21694 = ~n21693 | ~n21692;
  assign n21703 = ~n21695 & ~n21694;
  assign n21697 = ~n35376 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n21696 = ~n35866 | ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n21701 = ~n21697 | ~n21696;
  assign n21699 = ~n36457 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n21698 = ~n37332 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n21700 = ~n21699 | ~n21698;
  assign n21702 = ~n21701 & ~n21700;
  assign n21758 = ~n21703 | ~n21702;
  assign n21704 = ~n21758;
  assign n21706 = ~n26147 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n21705 = ~n20338 | ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n21710 = ~n21706 | ~n21705;
  assign n21708 = ~n26095 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n21707 = ~n25836 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n21709 = ~n21708 | ~n21707;
  assign n21718 = ~n21710 & ~n21709;
  assign n21712 = ~n26146 | ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n21711 = ~n26100 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n21716 = ~n21712 | ~n21711;
  assign n21714 = ~n26048 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n21713 = ~n25744 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n21715 = ~n21714 | ~n21713;
  assign n21717 = ~n21716 & ~n21715;
  assign n21735 = n21718 & n21717;
  assign n21719 = ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n21723 = ~n22211 & ~n21719;
  assign n21721 = ~n25827 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n21720 = ~n25810 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n21722 = ~n21721 | ~n21720;
  assign n21727 = ~n21723 & ~n21722;
  assign n21725 = n26139 | n26136;
  assign n21724 = n22328 | n21299;
  assign n21726 = n21725 & n21724;
  assign n21733 = ~n21727 | ~n21726;
  assign n21731 = n20333 & P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n21729 = ~n21791 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n21728 = ~n25783 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n21730 = ~n21729 | ~n21728;
  assign n21732 = n21731 | n21730;
  assign n21734 = ~n21733 & ~n21732;
  assign n21765 = ~n21761 | ~n25478;
  assign n39141 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n21738 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN & ~n31893;
  assign n31887 = n22361 ^ n21738;
  assign n21741 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN | ~n31887;
  assign n25658 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n21739 = ~n25658 & ~n31893;
  assign n21740 = ~n21739 | ~n20505;
  assign n21742 = ~n21741 | ~n21740;
  assign n21747 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN | ~n21742;
  assign n31245 = n21435 ^ ~n21742;
  assign n21744 = ~n21743;
  assign n31244 = n21745 ^ ~n21744;
  assign n21746 = ~n31245 | ~n31244;
  assign n21748 = ~n21747 | ~n21746;
  assign n34717 = P2_INSTADDRPOINTER_REG_3__SCAN_IN ^ n21748;
  assign n21749 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN | ~n21748;
  assign n21752 = ~n21751 | ~n21750;
  assign n36591 = ~n21755 | ~n21843;
  assign n21757 = ~n36591 | ~n37823;
  assign n36592 = ~n21756 | ~n21842;
  assign n21760 = ~n21757 | ~n36592;
  assign n25965 = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n21763 = n21761 ^ ~n25440;
  assign n21764 = ~n21763 | ~n21762;
  assign n39136 = P2_INSTADDRPOINTER_REG_8__SCAN_IN ^ ~n21765;
  assign n26977 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n40398 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n40318 = ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n40409 = ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n40103 = ~n40398 & ~n40409;
  assign n40107 = ~n40103 | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n40384 = ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n40360 = ~n40107 & ~n40384;
  assign n40153 = ~n40360 | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n21767 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n40328 = ~n40153 & ~n21767;
  assign n22167 = ~n40328 | ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n22169 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n40573 = ~n22167 & ~n22169;
  assign n21768 = ~n40573;
  assign n21772 = P2_EBX_REG_0__SCAN_IN | P2_EBX_REG_1__SCAN_IN;
  assign n21775 = ~n21773 | ~n20337;
  assign n21774 = ~n34908 | ~P2_EBX_REG_2__SCAN_IN;
  assign n21778 = ~n21776 | ~n20337;
  assign n21777 = ~n34908 | ~P2_EBX_REG_3__SCAN_IN;
  assign n21822 = ~n21778 | ~n21777;
  assign n21782 = ~n21780 | ~n20337;
  assign n21781 = ~n34908 | ~P2_EBX_REG_4__SCAN_IN;
  assign n21838 = ~n21782 | ~n21781;
  assign n21784 = ~n22408 | ~n20337;
  assign n38471 = ~P2_EBX_REG_5__SCAN_IN;
  assign n21783 = ~n34908 | ~n38471;
  assign n21844 = ~n21784 | ~n21783;
  assign n21786 = ~n26146 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n21785 = ~n26127 | ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n21790 = ~n21786 | ~n21785;
  assign n21788 = ~n20333 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n21787 = ~n25744 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n21789 = ~n21788 | ~n21787;
  assign n21816 = ~n21790 & ~n21789;
  assign n21796 = ~n21648 & ~n21792;
  assign n21794 = ~n25827 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n21793 = ~n25810 | ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n21795 = ~n21794 | ~n21793;
  assign n21798 = ~n21796 & ~n21795;
  assign n21797 = ~n21268 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n21814 = ~n21798 | ~n21797;
  assign n21800 = ~n22523 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n21799 = ~n26048 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n21804 = ~n21800 | ~n21799;
  assign n21802 = ~n26095 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n21801 = ~n26147 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n21803 = ~n21802 | ~n21801;
  assign n21812 = ~n21804 & ~n21803;
  assign n21806 = ~n25836 | ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n21805 = ~n25783 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n21810 = ~n21806 | ~n21805;
  assign n21808 = ~n20338 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n21807 = ~n26100 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n21809 = ~n21808 | ~n21807;
  assign n21811 = ~n21810 & ~n21809;
  assign n21813 = ~n21812 | ~n21811;
  assign n21815 = ~n21814 & ~n21813;
  assign n22358 = ~n21816 | ~n21815;
  assign n21817 = ~n22358;
  assign n21819 = ~n21817 | ~n20337;
  assign n21818 = ~n34908 | ~P2_EBX_REG_6__SCAN_IN;
  assign n21852 = ~n21819 | ~n21818;
  assign n21821 = ~n25478 | ~n20337;
  assign n35557 = ~P2_EBX_REG_7__SCAN_IN;
  assign n21820 = ~n34908 | ~n35557;
  assign n21866 = ~n34908 | ~P2_EBX_REG_9__SCAN_IN;
  assign n21893 = ~n34908 | ~P2_EBX_REG_12__SCAN_IN;
  assign n21863 = n34908 & P2_EBX_REG_13__SCAN_IN;
  assign n21901 = n34908 & P2_EBX_REG_16__SCAN_IN;
  assign n21907 = n34908 & P2_EBX_REG_17__SCAN_IN;
  assign n21911 = ~n34908 | ~P2_EBX_REG_18__SCAN_IN;
  assign n21918 = n34908 & P2_EBX_REG_19__SCAN_IN;
  assign n21916 = n34908 & P2_EBX_REG_20__SCAN_IN;
  assign n21926 = n34908 & P2_EBX_REG_21__SCAN_IN;
  assign n25205 = ~n34908 | ~P2_EBX_REG_22__SCAN_IN;
  assign n37860 = n25206 ^ ~n20709;
  assign n25227 = ~n37860 | ~n25478;
  assign n21824 = ~n21823 | ~n21822;
  assign n37025 = ~n21840 | ~n21824;
  assign n21825 = ~P2_EBX_REG_1__SCAN_IN | ~P2_EBX_REG_0__SCAN_IN;
  assign n21826 = ~n20337 & ~n21825;
  assign n35534 = ~n21833 & ~n21826;
  assign n21831 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN | ~n35534;
  assign n31882 = P2_INSTADDRPOINTER_REG_1__SCAN_IN ^ n35534;
  assign n21829 = ~n21827 | ~n20337;
  assign n21828 = ~n34908 | ~P2_EBX_REG_0__SCAN_IN;
  assign n35510 = n21829 & n21828;
  assign n31881 = ~n35510 & ~n25658;
  assign n21830 = ~n31882 | ~n31881;
  assign n31242 = ~n21831 | ~n21830;
  assign n38436 = n21833 ^ ~n21832;
  assign n31243 = n21435 ^ ~n38436;
  assign n21835 = ~n31242 | ~n31243;
  assign n21834 = ~n38436 | ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n34712 = ~n21835 | ~n21834;
  assign n21837 = ~n21836 | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n21839 = ~n21838;
  assign n38663 = n21840 ^ ~n21839;
  assign n35084 = ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n35090 = n38663 ^ ~n35084;
  assign n21841 = ~n38663 | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n21843 = ~n21842;
  assign n21847 = ~n21843 | ~n25440;
  assign n21846 = n21845 | n21844;
  assign n38476 = ~n21853 | ~n21846;
  assign n21848 = ~n21847 | ~n38476;
  assign n21850 = ~n36597 | ~n36596;
  assign n21849 = ~n21848 | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n25973 = ~n21850 | ~n21849;
  assign n21854 = ~n21853 | ~n21852;
  assign n37882 = ~n21860 | ~n21854;
  assign n21855 = ~n37882;
  assign n21861 = ~n21860 | ~n21859;
  assign n35556 = ~n25475 | ~n21861;
  assign n38853 = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n38688 = n21878 ^ ~n20471;
  assign n21862 = ~n40409 | ~n40109;
  assign n21870 = ~n40118 | ~n21862;
  assign n21864 = ~n21896 | ~n21863;
  assign n38705 = ~n21880 | ~n21864;
  assign n40020 = ~n38705 & ~n25440;
  assign n40290 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n40012 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n21865 = ~n40290 | ~n40012;
  assign n40123 = ~n40020 | ~n21865;
  assign n21867 = n20468 | n21866;
  assign n37662 = ~n21888 | ~n21867;
  assign n39536 = ~n25440 & ~n37662;
  assign n39714 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n21868 = ~n39141 | ~n39714;
  assign n40025 = ~n39536 | ~n21868;
  assign n21869 = n40123 & n40025;
  assign n21877 = ~n21870 | ~n21869;
  assign n21874 = ~n21894;
  assign n21873 = ~n21872 | ~n21871;
  assign n37679 = ~n21874 | ~n21873;
  assign n40000 = ~n25440 & ~n37679;
  assign n21876 = ~n40000;
  assign n21875 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN & ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n40027 = ~n21876 & ~n21875;
  assign n21882 = ~n21878;
  assign n21881 = ~n21880 | ~n21879;
  assign n38765 = ~n21882 | ~n21881;
  assign n40125 = ~n38765 & ~n25440;
  assign n21884 = n40125 | P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n40021 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN & ~n40000;
  assign n21883 = ~n40021;
  assign n21890 = ~n21884 | ~n21883;
  assign n21887 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN & ~n39536;
  assign n39139 = ~n35556 | ~n38853;
  assign n37145 = n21885 ^ n25475;
  assign n39140 = ~n37145 | ~n25478;
  assign n39143 = ~n39141 | ~n39140;
  assign n21886 = ~n39139 | ~n39143;
  assign n26958 = ~n21887 & ~n21886;
  assign n38415 = n21889 ^ n21888;
  assign n26960 = ~n38415 | ~n25478;
  assign n39996 = ~n26977 | ~n26960;
  assign n40022 = ~n26958 | ~n39996;
  assign n21892 = n21890 | n40022;
  assign n21891 = ~n40118 & ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n21899 = n21892 | n21891;
  assign n21895 = n21894 | n21893;
  assign n38740 = ~n21896 | ~n21895;
  assign n40165 = ~n25440 & ~n38740;
  assign n21898 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN & ~n40165;
  assign n21897 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN & ~n40020;
  assign n40119 = n21898 | n21897;
  assign n21900 = ~n21899 & ~n40119;
  assign n21902 = ~n21901;
  assign n38723 = n20427 ^ ~n21902;
  assign n21905 = ~n38723 | ~n25478;
  assign n40221 = n21905 & n40384;
  assign n40222 = ~n21905 & ~n40384;
  assign n21908 = ~n21907;
  assign n37427 = n20460 ^ ~n21908;
  assign n21909 = ~n37427 | ~n25478;
  assign n21910 = n21909 | n40368;
  assign n40546 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n21912 = ~n21911;
  assign n34615 = n21913 ^ ~n21912;
  assign n40160 = n34615 & n25478;
  assign n21915 = ~n21914 | ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n21917 = ~n21921 | ~n21916;
  assign n35489 = ~n21927 | ~n21917;
  assign n21920 = ~n21919 | ~n21918;
  assign n35946 = ~n21921 | ~n21920;
  assign n21922 = ~n25478 | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n40209 = n35946 | n21922;
  assign n21923 = ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n21924 = n35946 | n25440;
  assign n40210 = ~n21924 | ~n40318;
  assign n21929 = ~n25206;
  assign n21928 = ~n21927 | ~n21926;
  assign n35678 = ~n21929 | ~n21928;
  assign n29793 = n29331 | n30492;
  assign n21938 = ~n29793 | ~n21936;
  assign n21937 = ~n22176 | ~n21951;
  assign n21941 = ~n21938 | ~n21937;
  assign n21940 = n29331 | n21939;
  assign n21956 = ~n21941 | ~n21940;
  assign n21948 = ~n21942;
  assign n21946 = ~n27052 | ~n21943;
  assign n21944 = ~n21943;
  assign n21945 = ~n30492 | ~n21944;
  assign n21947 = ~n21946 | ~n21945;
  assign n21950 = ~n21948 | ~n21947;
  assign n21953 = ~n21950 | ~n21949;
  assign n21952 = ~n30492 | ~n21951;
  assign n21954 = ~n21953 | ~n21952;
  assign n21955 = ~n21954 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n21958 = ~n21956 & ~n21955;
  assign n21957 = ~P2_STATE2_REG_0__SCAN_IN & ~n34046;
  assign n21961 = ~n21958 & ~n21957;
  assign n21960 = n31666 | n21959;
  assign n21963 = ~n21961 | ~n21960;
  assign n21962 = n22120 | n31666;
  assign n21967 = ~n25167 | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n21966 = ~n25486 | ~P2_REIP_REG_22__SCAN_IN;
  assign n21971 = ~n21967 | ~n21966;
  assign n21969 = ~n25182 | ~P2_EBX_REG_22__SCAN_IN;
  assign n21968 = ~P2_PHYADDRPOINTER_REG_22__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n21970 = ~n21969 | ~n21968;
  assign n25175 = ~n21971 & ~n21970;
  assign n21974 = ~n25167 | ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n21973 = ~n25486 | ~P2_REIP_REG_20__SCAN_IN;
  assign n21978 = ~n21974 | ~n21973;
  assign n21976 = ~n25182 | ~P2_EBX_REG_20__SCAN_IN;
  assign n21975 = ~P2_PHYADDRPOINTER_REG_20__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n21977 = ~n21976 | ~n21975;
  assign n35495 = ~n21978 & ~n21977;
  assign n21980 = ~n25167 | ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n21979 = ~n25486 | ~P2_REIP_REG_18__SCAN_IN;
  assign n21984 = ~n21980 | ~n21979;
  assign n21982 = ~n25182 | ~P2_EBX_REG_18__SCAN_IN;
  assign n21981 = ~P2_PHYADDRPOINTER_REG_18__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n21983 = ~n21982 | ~n21981;
  assign n34625 = ~n21984 & ~n21983;
  assign n21986 = ~n25167 | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n21985 = ~n25486 | ~P2_REIP_REG_16__SCAN_IN;
  assign n21990 = ~n21986 | ~n21985;
  assign n21988 = ~n25182 | ~P2_EBX_REG_16__SCAN_IN;
  assign n21987 = ~P2_PHYADDRPOINTER_REG_16__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n21989 = ~n21988 | ~n21987;
  assign n35581 = ~n21990 & ~n21989;
  assign n21992 = ~n25167 | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n21991 = ~n25486 | ~P2_REIP_REG_14__SCAN_IN;
  assign n21996 = ~n21992 | ~n21991;
  assign n21994 = ~n25182 | ~P2_EBX_REG_14__SCAN_IN;
  assign n21993 = ~P2_PHYADDRPOINTER_REG_14__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n21995 = ~n21994 | ~n21993;
  assign n34468 = ~n21996 & ~n21995;
  assign n21998 = ~n25167 | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n21997 = ~n25486 | ~P2_REIP_REG_12__SCAN_IN;
  assign n22002 = ~n21998 | ~n21997;
  assign n22000 = ~n25182 | ~P2_EBX_REG_12__SCAN_IN;
  assign n21999 = ~P2_PHYADDRPOINTER_REG_12__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22001 = ~n22000 | ~n21999;
  assign n33877 = ~n22002 & ~n22001;
  assign n22004 = ~n25167 | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n22003 = ~n25486 | ~P2_REIP_REG_10__SCAN_IN;
  assign n22008 = ~n22004 | ~n22003;
  assign n22006 = ~n25182 | ~P2_EBX_REG_10__SCAN_IN;
  assign n22005 = ~P2_PHYADDRPOINTER_REG_10__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22007 = ~n22006 | ~n22005;
  assign n26965 = ~n22008 & ~n22007;
  assign n22010 = ~n25167 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n22009 = ~n25486 | ~P2_REIP_REG_8__SCAN_IN;
  assign n22014 = ~n22010 | ~n22009;
  assign n22012 = ~n25182 | ~P2_EBX_REG_8__SCAN_IN;
  assign n22011 = ~P2_PHYADDRPOINTER_REG_8__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22013 = ~n22012 | ~n22011;
  assign n32243 = ~n22014 & ~n22013;
  assign n22016 = ~n25167 | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n22015 = ~n25486 | ~P2_REIP_REG_6__SCAN_IN;
  assign n22020 = ~n22016 | ~n22015;
  assign n22018 = ~n25182 | ~P2_EBX_REG_6__SCAN_IN;
  assign n22017 = ~P2_PHYADDRPOINTER_REG_6__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22019 = ~n22018 | ~n22017;
  assign n25969 = ~n22020 & ~n22019;
  assign n22022 = ~n25167 | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n22021 = ~n25486 | ~P2_REIP_REG_4__SCAN_IN;
  assign n22026 = ~n22022 | ~n22021;
  assign n22024 = ~n25182 | ~P2_EBX_REG_4__SCAN_IN;
  assign n22023 = ~P2_PHYADDRPOINTER_REG_4__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22025 = ~n22024 | ~n22023;
  assign n33542 = ~n22026 & ~n22025;
  assign n22028 = ~n22027;
  assign n37823 = ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n22032 = ~n25448 & ~n37823;
  assign n22030 = ~n25486 | ~P2_REIP_REG_5__SCAN_IN;
  assign n22029 = ~n25182 | ~P2_EBX_REG_5__SCAN_IN;
  assign n22031 = ~n22030 | ~n22029;
  assign n22034 = ~n22032 & ~n22031;
  assign n22033 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n34509 = ~n22034 | ~n22033;
  assign n22038 = ~n25448 & ~n38853;
  assign n22036 = ~n25486 | ~P2_REIP_REG_7__SCAN_IN;
  assign n22035 = ~n25182 | ~P2_EBX_REG_7__SCAN_IN;
  assign n22037 = ~n22036 | ~n22035;
  assign n22040 = ~n22038 & ~n22037;
  assign n22039 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n33550 = ~n22040 | ~n22039;
  assign n22046 = ~n25167 | ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n22044 = n25486 & P2_REIP_REG_9__SCAN_IN;
  assign n22042 = ~n25182 | ~P2_EBX_REG_9__SCAN_IN;
  assign n22041 = ~P2_PHYADDRPOINTER_REG_9__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22043 = ~n22042 | ~n22041;
  assign n22045 = ~n22044 & ~n22043;
  assign n32962 = ~n22046 | ~n22045;
  assign n40334 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n22052 = n25448 | n40334;
  assign n22050 = n25486 & P2_REIP_REG_11__SCAN_IN;
  assign n22048 = ~n25182 | ~P2_EBX_REG_11__SCAN_IN;
  assign n22047 = ~P2_PHYADDRPOINTER_REG_11__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22049 = ~n22048 | ~n22047;
  assign n22051 = ~n22050 & ~n22049;
  assign n33703 = ~n22052 | ~n22051;
  assign n22056 = ~n25448 & ~n40012;
  assign n22054 = ~n25486 | ~P2_REIP_REG_13__SCAN_IN;
  assign n22053 = ~n25182 | ~P2_EBX_REG_13__SCAN_IN;
  assign n22055 = ~n22054 | ~n22053;
  assign n22058 = ~n22056 & ~n22055;
  assign n22057 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n34232 = ~n22058 | ~n22057;
  assign n22064 = ~n25167 | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n22062 = n25486 & P2_REIP_REG_15__SCAN_IN;
  assign n22060 = ~n25182 | ~P2_EBX_REG_15__SCAN_IN;
  assign n22059 = ~P2_PHYADDRPOINTER_REG_15__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22061 = ~n22060 | ~n22059;
  assign n22063 = ~n22062 & ~n22061;
  assign n34777 = ~n22064 | ~n22063;
  assign n22068 = ~n25448 & ~n40368;
  assign n22066 = ~n25486 | ~P2_REIP_REG_17__SCAN_IN;
  assign n22065 = ~n25182 | ~P2_EBX_REG_17__SCAN_IN;
  assign n22067 = ~n22066 | ~n22065;
  assign n22070 = ~n22068 & ~n22067;
  assign n22069 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n36043 = ~n22070 | ~n22069;
  assign n22077 = ~n25167 | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n22071 = ~P2_REIP_REG_19__SCAN_IN;
  assign n22075 = ~n21972 & ~n22071;
  assign n22073 = ~n25182 | ~P2_EBX_REG_19__SCAN_IN;
  assign n22072 = ~P2_PHYADDRPOINTER_REG_19__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22074 = ~n22073 | ~n22072;
  assign n22076 = ~n22075 & ~n22074;
  assign n35951 = ~n22077 | ~n22076;
  assign n22084 = ~n25167 | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n22078 = ~P2_REIP_REG_21__SCAN_IN;
  assign n22082 = ~n21972 & ~n22078;
  assign n22080 = ~n25182 | ~P2_EBX_REG_21__SCAN_IN;
  assign n22079 = ~P2_PHYADDRPOINTER_REG_21__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n22081 = ~n22080 | ~n22079;
  assign n22083 = ~n22082 & ~n22081;
  assign n35683 = ~n22084 | ~n22083;
  assign n22089 = n35516 | n22088;
  assign n22118 = n22122 | n22089;
  assign n34073 = ~READY21_REG_SCAN_IN | ~READY12_REG_SCAN_IN;
  assign n25567 = ~n29821 | ~n34073;
  assign n27360 = ~P2_STATE_REG_1__SCAN_IN;
  assign n27446 = ~P2_STATE_REG_0__SCAN_IN & ~n27360;
  assign n27361 = ~P2_STATE_REG_2__SCAN_IN;
  assign n27839 = ~n27446 | ~n27361;
  assign n22090 = ~n27839;
  assign n27785 = ~n22090;
  assign n22091 = ~P2_STATE_REG_0__SCAN_IN & ~P2_STATE_REG_1__SCAN_IN;
  assign n27436 = ~P2_STATE_REG_2__SCAN_IN | ~n22091;
  assign n30125 = ~n27785 | ~n27436;
  assign n22092 = ~n30492 & ~n30125;
  assign n22093 = ~n22092 & ~n34783;
  assign n22096 = ~n22175 & ~n22093;
  assign n22094 = ~n34783 | ~n25564;
  assign n22095 = ~n22094 & ~n30125;
  assign n22097 = n22096 | n22095;
  assign n22102 = ~n25567 & ~n22097;
  assign n22098 = ~n25608;
  assign n22099 = ~n22098 | ~n40626;
  assign n22101 = ~n22100 & ~n22099;
  assign n22116 = ~n22102 & ~n22101;
  assign n22104 = ~n22360 & ~n29786;
  assign n22108 = ~n22104 & ~n22103;
  assign n22123 = ~n35016 | ~n30492;
  assign n22105 = ~n22123 | ~n35516;
  assign n22106 = ~n22105 | ~n40860;
  assign n22107 = ~n22106 | ~n34783;
  assign n22113 = ~n22108 | ~n22107;
  assign n22109 = ~n22153;
  assign n22111 = n22110 & n22109;
  assign n22112 = ~n29336 & ~n22111;
  assign n25574 = ~n22113 & ~n22112;
  assign n22115 = n22114 & n25574;
  assign n22117 = n22116 & n22115;
  assign n22125 = n22118 & n22117;
  assign n22119 = ~n35516 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n22121 = n22120 | n22119;
  assign n22124 = n27013 | n22123;
  assign n22126 = ~n22125 | ~n22124;
  assign n30818 = ~n29336 | ~n30492;
  assign n22131 = ~n30818;
  assign n22133 = n22132 | n22131;
  assign n39129 = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN | ~P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n25959 = ~P2_INSTADDRPOINTER_REG_4__SCAN_IN | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n25963 = ~n34831 & ~n25959;
  assign n22134 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN | ~n25963;
  assign n39715 = ~n39129 & ~n22134;
  assign n26975 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN | ~n39715;
  assign n40331 = ~n26977 & ~n26975;
  assign n22165 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN | ~n40331;
  assign n22159 = ~n22165;
  assign n34726 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n33171 = ~n34726 & ~n25658;
  assign n22156 = ~n33171;
  assign n22137 = ~n22135;
  assign n22138 = ~n22137 | ~n22136;
  assign n22140 = ~n22138 | ~n34783;
  assign n22141 = ~n22140 | ~n22139;
  assign n22149 = ~n22142 | ~n22141;
  assign n22144 = ~n22143;
  assign n22145 = ~n22144 | ~n25690;
  assign n30003 = ~n29793 | ~n29786;
  assign n22146 = ~n22145 | ~n30003;
  assign n22148 = ~n22147 | ~n22146;
  assign n25609 = ~n22149 & ~n22148;
  assign n22150 = ~n25608 & ~n29793;
  assign n22151 = ~n22150 & ~n25855;
  assign n22152 = ~n25609 | ~n22151;
  assign n33170 = ~n22152 | ~n22174;
  assign n33176 = ~n22156 & ~n33170;
  assign n22158 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN | ~n33176;
  assign n22154 = ~n22370 & ~n22153;
  assign n25617 = ~n22155 | ~n22154;
  assign n30075 = ~n25617 & ~n25691;
  assign n33158 = n22174 & n30075;
  assign n33156 = ~n21435 | ~n22156;
  assign n22157 = ~n33158 | ~n33156;
  assign n40332 = ~n22158 | ~n22157;
  assign n40152 = ~n22159 | ~n40332;
  assign n34065 = ~n22174 & ~n40691;
  assign n22161 = ~n33158;
  assign n40148 = ~n22161 | ~n33170;
  assign n33157 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN | ~n33171;
  assign n22163 = ~n40148 | ~n33157;
  assign n22162 = n33156 & n33170;
  assign n22164 = ~n22163 & ~n22162;
  assign n25962 = ~n34065 & ~n22164;
  assign n22166 = ~n22165 | ~n40148;
  assign n40173 = ~n25962 | ~n22166;
  assign n22180 = ~n22174;
  assign n25568 = ~n22175 | ~n27052;
  assign n22178 = ~n25568;
  assign n30078 = n25617 | n22176;
  assign n30073 = ~n29336 | ~n40626;
  assign n22177 = ~n30078 | ~n30073;
  assign n22179 = ~n22178 & ~n22177;
  assign n40710 = ~n22180 & ~n22179;
  assign n22185 = ~n22389 & ~n20831;
  assign n22183 = ~n25513 | ~P2_REIP_REG_22__SCAN_IN;
  assign n22182 = ~n25514 | ~P2_EAX_REG_22__SCAN_IN;
  assign n22184 = ~n22183 | ~n22182;
  assign n25281 = ~n22185 & ~n22184;
  assign n22187 = ~n25513 | ~P2_REIP_REG_20__SCAN_IN;
  assign n22186 = ~n25514 | ~P2_EAX_REG_20__SCAN_IN;
  assign n22189 = ~n22187 | ~n22186;
  assign n22188 = ~n22389 & ~n21923;
  assign n35502 = ~n22189 & ~n22188;
  assign n22191 = ~n25513 | ~P2_REIP_REG_18__SCAN_IN;
  assign n22190 = ~n25514 | ~P2_EAX_REG_18__SCAN_IN;
  assign n22193 = ~n22191 | ~n22190;
  assign n22192 = ~n22389 & ~n40546;
  assign n34623 = ~n22193 & ~n22192;
  assign n22196 = ~n25513 | ~P2_REIP_REG_16__SCAN_IN;
  assign n22195 = ~n25514 | ~P2_EAX_REG_16__SCAN_IN;
  assign n22198 = ~n22196 | ~n22195;
  assign n22197 = ~n22389 & ~n40384;
  assign n35359 = ~n22198 & ~n22197;
  assign n22200 = ~n25514 | ~P2_EAX_REG_14__SCAN_IN;
  assign n22199 = ~n25513 | ~P2_REIP_REG_14__SCAN_IN;
  assign n22239 = ~n22200 | ~n22199;
  assign n22237 = ~n22571 | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n22202 = ~n26127 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n22201 = ~n25810 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n22206 = ~n22202 | ~n22201;
  assign n22204 = ~n20333 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n22203 = ~n25827 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n22205 = ~n22204 | ~n22203;
  assign n22234 = ~n22206 & ~n22205;
  assign n22210 = ~n26132 & ~n22207;
  assign n22209 = ~n21648 & ~n22208;
  assign n22215 = ~n22210 & ~n22209;
  assign n22213 = ~n26137 & ~n40787;
  assign n36001 = ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n22212 = ~n22211 & ~n36001;
  assign n22214 = ~n22213 & ~n22212;
  assign n22232 = ~n22215 | ~n22214;
  assign n22217 = ~n26146 | ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n22216 = ~n20338 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n22221 = ~n22217 | ~n22216;
  assign n22219 = ~n22341 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n22218 = ~n25744 | ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n22220 = ~n22219 | ~n22218;
  assign n22230 = ~n22221 & ~n22220;
  assign n26139 = ~n22222;
  assign n22523 = ~n26139;
  assign n22224 = ~n22523 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n22223 = ~n20339 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n22228 = ~n22224 | ~n22223;
  assign n22226 = ~n26147 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n22225 = ~n25836 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n22227 = ~n22226 | ~n22225;
  assign n22229 = ~n22228 & ~n22227;
  assign n22231 = ~n22230 | ~n22229;
  assign n22233 = ~n22232 & ~n22231;
  assign n34463 = ~n22234 | ~n22233;
  assign n22235 = ~n25564 | ~n37335;
  assign n22236 = ~n34463 | ~n22420;
  assign n22238 = ~n22237 | ~n22236;
  assign n33656 = ~n22239 & ~n22238;
  assign n22274 = ~n25513 | ~P2_REIP_REG_12__SCAN_IN;
  assign n22241 = ~n20333 | ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n22240 = ~n25810 | ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n22245 = ~n22241 | ~n22240;
  assign n22243 = ~n26127 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n22242 = ~n21791 | ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n22244 = ~n22243 | ~n22242;
  assign n22272 = ~n22245 & ~n22244;
  assign n22249 = ~n26069 & ~n22246;
  assign n22248 = ~n25753 & ~n22247;
  assign n22254 = ~n22249 & ~n22248;
  assign n22252 = ~n26132 & ~n22250;
  assign n36056 = ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n22251 = ~n22211 & ~n36056;
  assign n22253 = ~n22252 & ~n22251;
  assign n22270 = ~n22254 | ~n22253;
  assign n22256 = ~n20338 | ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n22255 = ~n20339 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n22260 = ~n22256 | ~n22255;
  assign n22258 = ~n22523 | ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n22257 = ~n25744 | ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n22259 = ~n22258 | ~n22257;
  assign n22268 = ~n22260 & ~n22259;
  assign n22262 = ~n26095 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n22261 = ~n25836 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n22266 = ~n22262 | ~n22261;
  assign n22264 = ~n26146 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n22263 = ~n26147 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n22265 = ~n22264 | ~n22263;
  assign n22267 = ~n22266 & ~n22265;
  assign n22269 = ~n22268 | ~n22267;
  assign n22271 = ~n22270 & ~n22269;
  assign n33874 = ~n22272 | ~n22271;
  assign n22273 = ~n33874 | ~n22420;
  assign n22278 = ~n22274 | ~n22273;
  assign n22276 = ~n25514 | ~P2_EAX_REG_12__SCAN_IN;
  assign n22275 = ~n22571 | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n22277 = ~n22276 | ~n22275;
  assign n32110 = ~n22278 & ~n22277;
  assign n22312 = ~n25513 | ~P2_REIP_REG_10__SCAN_IN;
  assign n22280 = ~n26127 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n22279 = ~n25827 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n22284 = ~n22280 | ~n22279;
  assign n22282 = ~n20333 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n22281 = ~n25810 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n22283 = ~n22282 | ~n22281;
  assign n22310 = ~n22284 & ~n22283;
  assign n37448 = ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n22287 = ~n22285 & ~n37448;
  assign n39645 = ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n22286 = ~n26139 & ~n39645;
  assign n22292 = ~n22287 & ~n22286;
  assign n22290 = ~n21549 & ~n22288;
  assign n36226 = ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n22289 = ~n21535 & ~n36226;
  assign n22291 = ~n22290 & ~n22289;
  assign n22308 = ~n22292 | ~n22291;
  assign n22294 = ~n21268 | ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n22293 = ~n21791 | ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n22298 = ~n22294 | ~n22293;
  assign n22296 = ~n26147 | ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n22295 = ~n22341 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n22297 = ~n22296 | ~n22295;
  assign n22306 = ~n22298 & ~n22297;
  assign n22300 = ~n26095 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n22299 = ~n26100 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n22304 = ~n22300 | ~n22299;
  assign n22302 = ~n26146 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n22301 = ~n20338 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n22303 = ~n22302 | ~n22301;
  assign n22305 = ~n22304 & ~n22303;
  assign n22307 = ~n22306 | ~n22305;
  assign n22309 = ~n22308 & ~n22307;
  assign n33214 = ~n22310 | ~n22309;
  assign n22311 = ~n33214 | ~n22420;
  assign n22316 = ~n22312 | ~n22311;
  assign n22314 = ~n22571 | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n22313 = ~n25514 | ~P2_EAX_REG_10__SCAN_IN;
  assign n22315 = ~n22314 | ~n22313;
  assign n26983 = ~n22316 & ~n22315;
  assign n22353 = ~n25513 | ~P2_REIP_REG_8__SCAN_IN;
  assign n22318 = ~n20333 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n22317 = ~n25810 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n22322 = ~n22318 | ~n22317;
  assign n22320 = ~n25836 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n22319 = ~n25783 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n22321 = ~n22320 | ~n22319;
  assign n22351 = ~n22322 & ~n22321;
  assign n22326 = ~n21648 & ~n22323;
  assign n22325 = ~n25753 & ~n22324;
  assign n22332 = ~n22326 & ~n22325;
  assign n22330 = ~n22211 & ~n35840;
  assign n22327 = ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n22329 = ~n22328 & ~n22327;
  assign n22331 = ~n22330 & ~n22329;
  assign n22349 = ~n22332 | ~n22331;
  assign n22334 = ~n26095 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n22333 = ~n25744 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n22338 = ~n22334 | ~n22333;
  assign n22336 = ~n26147 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n22335 = ~n26100 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n22337 = ~n22336 | ~n22335;
  assign n22347 = ~n22338 & ~n22337;
  assign n22340 = ~n26146 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n22339 = ~n20338 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n22345 = ~n22340 | ~n22339;
  assign n22343 = ~n22523 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n22342 = ~n22341 | ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n22344 = ~n22343 | ~n22342;
  assign n22346 = ~n22345 & ~n22344;
  assign n22348 = ~n22347 | ~n22346;
  assign n22350 = ~n22349 & ~n22348;
  assign n32237 = ~n22351 | ~n22350;
  assign n22352 = ~n32237 | ~n22420;
  assign n22357 = ~n22353 | ~n22352;
  assign n22355 = ~n22571 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n22354 = ~n25514 | ~P2_EAX_REG_8__SCAN_IN;
  assign n22356 = ~n22355 | ~n22354;
  assign n30575 = ~n22357 & ~n22356;
  assign n22415 = ~n22358 | ~n22420;
  assign n22403 = ~n22420 | ~n22359;
  assign n30543 = ~n22360;
  assign n22363 = ~n30543 & ~P2_STATE2_REG_3__SCAN_IN;
  assign n22362 = ~n22361 & ~n22568;
  assign n22365 = ~n22363 & ~n22362;
  assign n22364 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_STATE2_REG_3__SCAN_IN;
  assign n22378 = ~n22365 | ~n22364;
  assign n22367 = ~n20354 & ~n34726;
  assign n27841 = ~P2_REIP_REG_1__SCAN_IN;
  assign n22366 = ~n25415 & ~n27841;
  assign n22381 = ~n22378 & ~n22379;
  assign n22369 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~P2_STATE2_REG_3__SCAN_IN;
  assign n22368 = ~n31893 | ~n22420;
  assign n30490 = ~n22369 | ~n22368;
  assign n22383 = ~n20354 & ~n22370;
  assign n22372 = n22383 | n22371;
  assign n30532 = ~n30490 & ~n22372;
  assign n22374 = ~n25513 | ~P2_REIP_REG_0__SCAN_IN;
  assign n22373 = ~n40626 | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n22377 = ~n22374 | ~n22373;
  assign n22375 = ~n25855 | ~P2_EAX_REG_0__SCAN_IN;
  assign n22376 = ~n22375 | ~n37335;
  assign n30531 = ~n22377 & ~n22376;
  assign n30481 = ~n30532 & ~n30531;
  assign n22387 = ~n22381 & ~n22380;
  assign n22384 = ~n22382 & ~n22568;
  assign n22386 = ~n22384 & ~n22383;
  assign n22385 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_STATE2_REG_3__SCAN_IN;
  assign n22388 = ~n22386 | ~n22385;
  assign n31195 = n22388 ^ ~n22387;
  assign n22391 = ~n22389 & ~n21435;
  assign n27840 = ~P2_REIP_REG_2__SCAN_IN;
  assign n22390 = ~n25415 & ~n27840;
  assign n22393 = ~n22391 & ~n22390;
  assign n22392 = ~n25514 | ~P2_EAX_REG_2__SCAN_IN;
  assign n31194 = ~n22393 | ~n22392;
  assign n22395 = ~n22571 | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n22394 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P2_STATE2_REG_3__SCAN_IN;
  assign n22400 = ~n22395 | ~n22394;
  assign n22398 = ~n25514 | ~P2_EAX_REG_3__SCAN_IN;
  assign n22397 = n22396 | n22568;
  assign n22399 = ~n22398 | ~n22397;
  assign n22402 = ~n22400 & ~n22399;
  assign n22401 = ~n25513 | ~P2_REIP_REG_3__SCAN_IN;
  assign n33202 = ~n22402 | ~n22401;
  assign n27493 = ~P2_REIP_REG_4__SCAN_IN;
  assign n22405 = ~n25415 & ~n27493;
  assign n22404 = ~n22389 & ~n35084;
  assign n22407 = ~n22405 & ~n22404;
  assign n22406 = ~n25514 | ~P2_EAX_REG_4__SCAN_IN;
  assign n35074 = ~n22407 | ~n22406;
  assign n22410 = ~n35075 | ~n35074;
  assign n22409 = ~n22420 | ~n22408;
  assign n27503 = ~P2_REIP_REG_5__SCAN_IN;
  assign n22412 = ~n25415 & ~n27503;
  assign n22411 = ~n22389 & ~n37823;
  assign n22414 = ~n22412 & ~n22411;
  assign n22413 = ~n25514 | ~P2_EAX_REG_5__SCAN_IN;
  assign n35071 = ~n22414 | ~n22413;
  assign n37878 = ~P2_REIP_REG_6__SCAN_IN;
  assign n22417 = ~n25415 & ~n37878;
  assign n22416 = ~n22389 & ~n25965;
  assign n22419 = ~n22417 & ~n22416;
  assign n22418 = ~n25514 | ~P2_EAX_REG_6__SCAN_IN;
  assign n25956 = ~n22419 | ~n22418;
  assign n22421 = ~n22420 | ~n25478;
  assign n30652 = ~n22422 | ~n22421;
  assign n38844 = ~P2_REIP_REG_7__SCAN_IN;
  assign n22424 = ~n25415 & ~n38844;
  assign n22423 = ~n22389 & ~n38853;
  assign n22426 = ~n22424 & ~n22423;
  assign n22425 = ~n25514 | ~P2_EAX_REG_7__SCAN_IN;
  assign n30651 = ~n22426 | ~n22425;
  assign n30574 = ~n30652 | ~n30651;
  assign n31116 = ~n30575 & ~n30574;
  assign n22428 = ~n25514 | ~P2_EAX_REG_9__SCAN_IN;
  assign n22427 = ~n25513 | ~P2_REIP_REG_9__SCAN_IN;
  assign n22460 = ~n22428 | ~n22427;
  assign n22430 = ~n26146 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n22429 = ~n25836 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n22434 = ~n22430 | ~n22429;
  assign n22432 = ~n26147 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n22431 = ~n20338 | ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n22433 = ~n22432 | ~n22431;
  assign n22442 = ~n22434 & ~n22433;
  assign n22436 = ~n22523 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n22435 = ~n26048 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n22440 = ~n22436 | ~n22435;
  assign n22438 = ~n26095 | ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n22437 = ~n25744 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n22439 = ~n22438 | ~n22437;
  assign n22441 = ~n22440 & ~n22439;
  assign n22458 = ~n22442 | ~n22441;
  assign n22444 = ~n26127 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n22443 = ~n25810 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n22448 = ~n22444 | ~n22443;
  assign n22446 = ~n20333 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n22445 = ~n21791 | ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n22447 = ~n22446 | ~n22445;
  assign n22456 = ~n22448 & ~n22447;
  assign n22450 = ~n21268 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n22449 = ~n25827 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n22454 = ~n22450 | ~n22449;
  assign n22452 = ~n26100 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n22451 = ~n20339 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n22453 = ~n22452 | ~n22451;
  assign n22455 = ~n22454 & ~n22453;
  assign n22457 = ~n22456 | ~n22455;
  assign n25737 = ~n22458 & ~n22457;
  assign n22459 = ~n25737 & ~n22568;
  assign n22462 = ~n22460 & ~n22459;
  assign n22461 = ~n22571 | ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n31115 = ~n22462 | ~n22461;
  assign n22464 = ~n25514 | ~P2_EAX_REG_11__SCAN_IN;
  assign n22463 = ~n25513 | ~P2_REIP_REG_11__SCAN_IN;
  assign n22496 = ~n22464 | ~n22463;
  assign n22466 = ~n26146 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n22465 = ~n20338 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n22470 = ~n22466 | ~n22465;
  assign n22468 = ~n26095 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n22467 = ~n26048 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n22469 = ~n22468 | ~n22467;
  assign n22478 = ~n22470 & ~n22469;
  assign n22472 = ~n26100 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n22471 = ~n25744 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n22476 = ~n22472 | ~n22471;
  assign n22474 = ~n26147 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n22473 = ~n22523 | ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n22475 = ~n22474 | ~n22473;
  assign n22477 = ~n22476 & ~n22475;
  assign n22494 = ~n22478 | ~n22477;
  assign n22480 = ~n21268 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n22479 = ~n26127 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n22484 = ~n22480 | ~n22479;
  assign n22482 = ~n20333 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n22481 = ~n25810 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n22483 = ~n22482 | ~n22481;
  assign n22492 = ~n22484 & ~n22483;
  assign n22486 = ~n21791 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n22485 = ~n25827 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n22490 = ~n22486 | ~n22485;
  assign n22488 = ~n25836 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n22487 = ~n20339 | ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n22489 = ~n22488 | ~n22487;
  assign n22491 = ~n22490 & ~n22489;
  assign n22493 = ~n22492 | ~n22491;
  assign n25739 = ~n22494 & ~n22493;
  assign n22495 = ~n25739 & ~n22568;
  assign n22498 = ~n22496 & ~n22495;
  assign n22497 = ~n22571 | ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n31874 = ~n22498 | ~n22497;
  assign n22500 = ~n22571 | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n22499 = ~n25513 | ~P2_REIP_REG_13__SCAN_IN;
  assign n22533 = ~n22500 | ~n22499;
  assign n22502 = ~n20338 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n22501 = ~n26100 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n22506 = ~n22502 | ~n22501;
  assign n22504 = ~n26095 | ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n22503 = ~n26048 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n22505 = ~n22504 | ~n22503;
  assign n22514 = ~n22506 & ~n22505;
  assign n22508 = ~n25744 | ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n22507 = ~n25783 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n22512 = ~n22508 | ~n22507;
  assign n22510 = ~n26146 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n22509 = ~n25836 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n22511 = ~n22510 | ~n22509;
  assign n22513 = ~n22512 & ~n22511;
  assign n22531 = ~n22514 | ~n22513;
  assign n22516 = ~n25827 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n22515 = ~n25810 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n22520 = ~n22516 | ~n22515;
  assign n22518 = ~n26127 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n22517 = ~n20333 | ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n22519 = ~n22518 | ~n22517;
  assign n22529 = ~n22520 & ~n22519;
  assign n22522 = ~n21268 | ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n22521 = ~n21791 | ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n22527 = ~n22522 | ~n22521;
  assign n22525 = ~n26147 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n22524 = ~n22523 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n22526 = ~n22525 | ~n22524;
  assign n22528 = ~n22527 & ~n22526;
  assign n22530 = ~n22529 | ~n22528;
  assign n25740 = ~n22531 & ~n22530;
  assign n22532 = ~n25740 & ~n22568;
  assign n22535 = ~n22533 & ~n22532;
  assign n22534 = ~n25514 | ~P2_EAX_REG_13__SCAN_IN;
  assign n33139 = ~n22535 | ~n22534;
  assign n22537 = ~n25514 | ~P2_EAX_REG_15__SCAN_IN;
  assign n22536 = ~n25513 | ~P2_REIP_REG_15__SCAN_IN;
  assign n22570 = ~n22537 | ~n22536;
  assign n22539 = ~n22523 | ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n22538 = ~n26048 | ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n22543 = ~n22539 | ~n22538;
  assign n22541 = ~n26146 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n22540 = ~n25783 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n22542 = ~n22541 | ~n22540;
  assign n22551 = ~n22543 & ~n22542;
  assign n22545 = ~n26147 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n22544 = ~n26100 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n22549 = ~n22545 | ~n22544;
  assign n22547 = ~n26095 | ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n22546 = ~n20338 | ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n22548 = ~n22547 | ~n22546;
  assign n22550 = ~n22549 & ~n22548;
  assign n22567 = ~n22551 | ~n22550;
  assign n22553 = ~n21791 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n22552 = ~n25827 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n22557 = ~n22553 | ~n22552;
  assign n22555 = ~n26127 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n22554 = ~n20333 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n22556 = ~n22555 | ~n22554;
  assign n22565 = ~n22557 & ~n22556;
  assign n22559 = ~n21268 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n22558 = ~n25836 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n22563 = ~n22559 | ~n22558;
  assign n22561 = ~n25744 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n22560 = ~n25810 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n22562 = ~n22561 | ~n22560;
  assign n22564 = ~n22563 & ~n22562;
  assign n22566 = ~n22565 | ~n22564;
  assign n25741 = ~n22567 & ~n22566;
  assign n22569 = ~n25741 & ~n22568;
  assign n22573 = ~n22570 & ~n22569;
  assign n22572 = ~n22571 | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n33606 = ~n22573 | ~n22572;
  assign n37425 = ~P2_REIP_REG_17__SCAN_IN;
  assign n22575 = ~n25415 & ~n37425;
  assign n22574 = ~n22389 & ~n40368;
  assign n22577 = ~n22575 & ~n22574;
  assign n22576 = ~n25514 | ~P2_EAX_REG_17__SCAN_IN;
  assign n35670 = ~n22577 | ~n22576;
  assign n22579 = ~n25415 & ~n22071;
  assign n22578 = ~n22389 & ~n40318;
  assign n22581 = ~n22579 & ~n22578;
  assign n22580 = ~n25514 | ~P2_EAX_REG_19__SCAN_IN;
  assign n25853 = ~n22581 | ~n22580;
  assign n22583 = ~n25415 & ~n22078;
  assign n22582 = ~n22389 & ~n40434;
  assign n22585 = ~n22583 & ~n22582;
  assign n22584 = ~n25514 | ~P2_EAX_REG_21__SCAN_IN;
  assign n35690 = ~n22585 | ~n22584;
  assign n25277 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n25272 = ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n25287 = ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n25301 = ~n25272 & ~n25287;
  assign n25169 = ~n25167 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n25168 = ~n25486 | ~P2_REIP_REG_24__SCAN_IN;
  assign n25173 = ~n25169 | ~n25168;
  assign n25171 = ~n25182 | ~P2_EBX_REG_24__SCAN_IN;
  assign n25170 = ~P2_PHYADDRPOINTER_REG_24__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n25172 = ~n25171 | ~n25170;
  assign n37917 = ~n25173 & ~n25172;
  assign n25282 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n25179 = ~n25448 & ~n25282;
  assign n25177 = ~n25486 | ~P2_REIP_REG_23__SCAN_IN;
  assign n25176 = ~n25182 | ~P2_EBX_REG_23__SCAN_IN;
  assign n25178 = ~n25177 | ~n25176;
  assign n25181 = ~n25179 & ~n25178;
  assign n25180 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n38249 = ~n25181 | ~n25180;
  assign n25186 = ~n25448 & ~n25287;
  assign n25184 = ~n25486 | ~P2_REIP_REG_25__SCAN_IN;
  assign n25183 = ~n25182 | ~P2_EBX_REG_25__SCAN_IN;
  assign n25185 = ~n25184 | ~n25183;
  assign n25188 = ~n25186 & ~n25185;
  assign n25187 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n38063 = ~n25188 | ~n25187;
  assign n25195 = n25448 | n25272;
  assign n25193 = ~n25486 | ~P2_REIP_REG_26__SCAN_IN;
  assign n25189 = ~P2_EBX_REG_26__SCAN_IN;
  assign n25191 = n25488 | n25189;
  assign n25190 = ~P2_PHYADDRPOINTER_REG_26__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n25192 = n25191 & n25190;
  assign n25194 = n25193 & n25192;
  assign n25256 = ~n25195 | ~n25194;
  assign n25220 = n34908 & P2_EBX_REG_23__SCAN_IN;
  assign n25217 = n34908 & P2_EBX_REG_24__SCAN_IN;
  assign n25213 = ~n34908 | ~P2_EBX_REG_25__SCAN_IN;
  assign n25207 = n34908 & P2_EBX_REG_26__SCAN_IN;
  assign n25208 = ~n25215 | ~n25207;
  assign n39014 = ~n25240 | ~n25208;
  assign n25211 = ~n25227 | ~n20831;
  assign n25210 = ~n40439 | ~n40434;
  assign n25214 = n25219 | n25213;
  assign n38069 = ~n25215 | ~n25214;
  assign n25216 = ~n38069 & ~n25440;
  assign n40877 = ~n25216 & ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n25228 = ~n37920 & ~n25440;
  assign n40879 = ~n25228 & ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n25223 = n40877 | n40879;
  assign n25221 = ~n25220;
  assign n38251 = n25222 ^ ~n25221;
  assign n25229 = ~n38251 | ~n25478;
  assign n40580 = n25229 & n25282;
  assign n25224 = ~n25223 & ~n40580;
  assign n25225 = ~n25478 | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n40878 = ~n38069 & ~n25225;
  assign n25226 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN & ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n40578 = ~n25227 & ~n25226;
  assign n25231 = n40878 | n40578;
  assign n40882 = ~n25228 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n40697 = ~n25282 & ~n25229;
  assign n40581 = ~n40697;
  assign n25230 = ~n40882 | ~n40581;
  assign n25232 = ~n25231 & ~n25230;
  assign n25245 = ~n25238 | ~n25237;
  assign n25239 = n34908 & P2_EBX_REG_27__SCAN_IN;
  assign n25241 = n25240 & n25239;
  assign n39272 = n25241 | n25332;
  assign n25242 = ~n39272;
  assign n25243 = ~n25478 | ~n25272;
  assign n25244 = n39272 | n25243;
  assign n25376 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n25255 = n25448 | n25376;
  assign n25253 = ~n25486 | ~P2_REIP_REG_27__SCAN_IN;
  assign n25249 = ~P2_EBX_REG_27__SCAN_IN;
  assign n25251 = n25488 | n25249;
  assign n25250 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n25252 = n25251 & n25250;
  assign n25254 = n25253 & n25252;
  assign n25346 = ~n25255 | ~n25254;
  assign n25269 = ~n25301;
  assign n25298 = ~n40573 | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n40713 = ~n40152 & ~n25298;
  assign n25318 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN | ~n40713;
  assign n25420 = ~n25269 & ~n25318;
  assign n25271 = ~n25513 | ~P2_REIP_REG_26__SCAN_IN;
  assign n25270 = ~n22371 | ~P2_EAX_REG_26__SCAN_IN;
  assign n25274 = ~n25271 | ~n25270;
  assign n25273 = ~n22389 & ~n25272;
  assign n25313 = ~n25274 & ~n25273;
  assign n25276 = ~n25513 | ~P2_REIP_REG_24__SCAN_IN;
  assign n25275 = ~n25514 | ~P2_EAX_REG_24__SCAN_IN;
  assign n25279 = ~n25276 | ~n25275;
  assign n25278 = ~n22389 & ~n25277;
  assign n37915 = ~n25279 & ~n25278;
  assign n40567 = ~P2_REIP_REG_23__SCAN_IN;
  assign n25284 = ~n25415 & ~n40567;
  assign n25283 = ~n22389 & ~n25282;
  assign n25286 = ~n25284 & ~n25283;
  assign n25285 = ~n25514 | ~P2_EAX_REG_23__SCAN_IN;
  assign n26214 = ~n25286 | ~n25285;
  assign n40869 = ~P2_REIP_REG_25__SCAN_IN;
  assign n25289 = ~n25415 & ~n40869;
  assign n25288 = ~n22389 & ~n25287;
  assign n25291 = ~n25289 & ~n25288;
  assign n25290 = ~n25514 | ~P2_EAX_REG_25__SCAN_IN;
  assign n38067 = ~n25291 | ~n25290;
  assign n27810 = ~P2_REIP_REG_27__SCAN_IN;
  assign n25293 = ~n25415 & ~n27810;
  assign n25292 = ~n22389 & ~n25376;
  assign n25295 = ~n25293 & ~n25292;
  assign n25294 = ~n22371 | ~P2_EAX_REG_27__SCAN_IN;
  assign n25363 = ~n25295 | ~n25294;
  assign n25422 = ~n34065 & ~n40148;
  assign n25299 = ~n25298 | ~n40148;
  assign n25300 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN | ~n25299;
  assign n40715 = ~n40173 & ~n25300;
  assign n40923 = ~n25422 & ~n40715;
  assign n25302 = ~n25301 & ~n25422;
  assign n25426 = ~n40923 & ~n25302;
  assign n25329 = ~n25478 | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n25331 = ~n34908 | ~P2_EBX_REG_28__SCAN_IN;
  assign n25385 = ~n25332 | ~n25331;
  assign n25333 = n25332 | n25331;
  assign n39749 = ~n25385 | ~n25333;
  assign n25338 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n25345 = n25448 | n25338;
  assign n25343 = ~n25486 | ~P2_REIP_REG_28__SCAN_IN;
  assign n25339 = ~P2_EBX_REG_28__SCAN_IN;
  assign n25341 = n25488 | n25339;
  assign n25340 = ~P2_PHYADDRPOINTER_REG_28__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n25342 = n25341 & n25340;
  assign n25344 = n25343 & n25342;
  assign n25400 = ~n25345 | ~n25344;
  assign n25360 = ~n25513 | ~P2_REIP_REG_28__SCAN_IN;
  assign n25359 = ~n22371 | ~P2_EAX_REG_28__SCAN_IN;
  assign n25362 = ~n25360 | ~n25359;
  assign n25361 = ~n22389 & ~n25338;
  assign n25414 = ~n25362 & ~n25361;
  assign n25413 = ~n25364 | ~n25363;
  assign n25421 = ~n25376 & ~n25338;
  assign n25424 = ~n25421 | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n25381 = ~n25478 | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n25382 = n39749 | n25381;
  assign n25390 = ~n25383 | ~n25382;
  assign n25388 = ~n25390;
  assign n25384 = n34908 & P2_EBX_REG_29__SCAN_IN;
  assign n25386 = ~n25385 | ~n25384;
  assign n39935 = ~n25472 | ~n25386;
  assign n25387 = ~n25389;
  assign n25442 = ~n25390 | ~n25389;
  assign n25523 = ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n25399 = n25448 | n25523;
  assign n25393 = ~P2_EBX_REG_29__SCAN_IN;
  assign n25395 = n25488 | n25393;
  assign n25394 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n25397 = n25395 & n25394;
  assign n25396 = ~n21965 | ~P2_REIP_REG_29__SCAN_IN;
  assign n25398 = n25397 & n25396;
  assign n25456 = ~n25399 | ~n25398;
  assign n25512 = ~n25414 & ~n25413;
  assign n27816 = ~P2_REIP_REG_29__SCAN_IN;
  assign n25417 = ~n25415 & ~n27816;
  assign n25416 = ~n22389 & ~n25523;
  assign n25419 = ~n25417 & ~n25416;
  assign n25418 = ~n22371 | ~P2_EAX_REG_29__SCAN_IN;
  assign n25511 = ~n25419 | ~n25418;
  assign n25522 = ~n25421 | ~n25420;
  assign n25423 = ~n25422;
  assign n25425 = ~n25424 | ~n25423;
  assign n25556 = ~n25426 | ~n25425;
  assign n25439 = n34908 & P2_EBX_REG_30__SCAN_IN;
  assign n27060 = n25472 ^ ~n25439;
  assign n25444 = ~n25442 | ~n25523;
  assign n25468 = ~n25444 | ~n25443;
  assign n25553 = ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n25455 = n25448 | n25553;
  assign n25453 = ~n25486 | ~P2_REIP_REG_30__SCAN_IN;
  assign n25449 = ~P2_EBX_REG_30__SCAN_IN;
  assign n25451 = n25488 | n25449;
  assign n25450 = ~P2_PHYADDRPOINTER_REG_30__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n25452 = n25451 & n25450;
  assign n25454 = n25453 & n25452;
  assign n25495 = ~n25455 | ~n25454;
  assign n25471 = ~n25468 & ~n20402;
  assign n25469 = ~n25478 | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n25470 = ~n27060 & ~n25469;
  assign n25481 = ~n25471 & ~n25470;
  assign n25474 = ~n25472;
  assign n25473 = ~n20337 & ~P2_EBX_REG_30__SCAN_IN;
  assign n25477 = ~n25474 | ~n25473;
  assign n25476 = ~n25475 | ~n20337;
  assign n39888 = ~n25477 | ~n25476;
  assign n25479 = ~n39888 | ~n25478;
  assign n25480 = n25479 ^ ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n25506 = n25481 ^ ~n25480;
  assign n25657 = ~P2_INSTADDRPOINTER_REG_31__SCAN_IN | ~P2_STATE2_REG_0__SCAN_IN;
  assign n25484 = ~n25657;
  assign n25494 = ~n25485 | ~n25484;
  assign n25492 = ~n25486 | ~P2_REIP_REG_31__SCAN_IN;
  assign n25487 = ~P2_EBX_REG_31__SCAN_IN;
  assign n25490 = n25488 | n25487;
  assign n25489 = ~P2_PHYADDRPOINTER_REG_31__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n25491 = n25490 & n25489;
  assign n25493 = n25492 & n25491;
  assign n25499 = ~n25494 | ~n25493;
  assign n25497 = ~n25495;
  assign n25498 = ~n25497 & ~n25496;
  assign n37757 = n25499 ^ ~n25498;
  assign n25528 = P2_INSTADDRPOINTER_REG_31__SCAN_IN ^ ~n25501;
  assign n25526 = ~P2_REIP_REG_31__SCAN_IN | ~n40691;
  assign n25532 = ~n25506 | ~n40931;
  assign n25508 = ~n25513 | ~P2_REIP_REG_30__SCAN_IN;
  assign n25507 = ~n22371 | ~P2_EAX_REG_30__SCAN_IN;
  assign n25510 = ~n25508 | ~n25507;
  assign n25509 = ~n22389 & ~n25553;
  assign n25552 = ~n25510 & ~n25509;
  assign n25551 = ~n25512 | ~n25511;
  assign n25521 = ~n25552 & ~n25551;
  assign n25516 = ~n25513 | ~P2_REIP_REG_31__SCAN_IN;
  assign n25515 = ~n25514 | ~P2_EAX_REG_31__SCAN_IN;
  assign n25519 = ~n25516 | ~n25515;
  assign n25517 = ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n25518 = ~n22389 & ~n25517;
  assign n25520 = ~n25519 & ~n25518;
  assign n39881 = n25521 ^ ~n25520;
  assign n25530 = ~n40710 | ~n39881;
  assign n25524 = P2_INSTADDRPOINTER_REG_31__SCAN_IN ^ ~n25553;
  assign n25554 = ~n25523 & ~n25522;
  assign n25525 = ~n37757;
  assign n25527 = ~n40929 | ~n25525;
  assign n25529 = ~P2_INSTADDRPOINTER_REG_31__SCAN_IN | ~n25556;
  assign P2_U3015_Lock = ~n25532 | ~n25531;
  assign n35860 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign input_0 = keyinput_0 ^ READY12_REG_SCAN_IN;
  assign input_1 = keyinput_1 ^ READY21_REG_SCAN_IN;
  assign AND_1 = input_0 & input_1;
  assign input_2 = keyinput_2 ^ ~P2_STATE_REG_2__SCAN_IN;
  assign OR_2 = input_2 | AND_1;
  assign input_3 = keyinput_3 ^ ~P2_STATE_REG_1__SCAN_IN;
  assign OR_3 = input_3 | OR_2;
  assign input_4 = keyinput_4 ^ P2_STATE_REG_0__SCAN_IN;
  assign AND_4 = input_4 & OR_3;
  assign input_5 = keyinput_5 ^ ~P2_STATE2_REG_3__SCAN_IN;
  assign OR_5 = input_5 | AND_4;
  assign input_6 = keyinput_6 ^ P2_STATE2_REG_2__SCAN_IN;
  assign OR_6 = input_6 | OR_5;
  assign input_7 = keyinput_7 ^ ~P2_STATE2_REG_1__SCAN_IN;
  assign AND_7 = input_7 & OR_6;
  assign input_8 = keyinput_8 ^ P2_STATE2_REG_0__SCAN_IN;
  assign OR_8 = input_8 | AND_7;
  assign input_9 = keyinput_9 ^ ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign AND_9 = input_9 & OR_8;
  assign input_10 = keyinput_10 ^ P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign OR_10 = input_10 | AND_9;
  assign input_11 = keyinput_11 ^ ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign OR_11 = input_11 | OR_10;
  assign input_12 = keyinput_12 ^ P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign AND_12 = input_12 & OR_11;
  assign input_13 = keyinput_13 ^ P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign AND_13 = input_13 & AND_12;
  assign input_14 = keyinput_14 ^ ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign AND_14 = input_14 & AND_13;
  assign input_15 = keyinput_15 ^ P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign AND_15 = input_15 & AND_14;
  assign input_16 = keyinput_16 ^ ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign AND_16 = input_16 & AND_15;
  assign input_17 = keyinput_17 ^ P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign AND_17 = input_17 & AND_16;
  assign input_18 = keyinput_18 ^ ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign OR_18 = input_18 | AND_17;
  assign input_19 = keyinput_19 ^ ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign AND_19 = input_19 & OR_18;
  assign input_20 = keyinput_20 ^ ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign AND_20 = input_20 & AND_19;
  assign input_21 = keyinput_21 ^ P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign AND_21 = input_21 & AND_20;
  assign input_22 = keyinput_22 ^ P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign AND_22 = input_22 & AND_21;
  assign input_23 = keyinput_23 ^ ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign OR_23 = input_23 | AND_22;
  assign input_24 = keyinput_24 ^ P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign AND_24 = input_24 & OR_23;
  assign input_25 = keyinput_25 ^ P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign OR_25 = input_25 | AND_24;
  assign input_26 = keyinput_26 ^ P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign OR_26 = input_26 | OR_25;
  assign input_27 = keyinput_27 ^ P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign AND_27 = input_27 & OR_26;
  assign input_28 = keyinput_28 ^ ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign OR_28 = input_28 | AND_27;
  assign input_29 = keyinput_29 ^ P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign OR_29 = input_29 | OR_28;
  assign input_30 = keyinput_30 ^ P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign OR_30 = input_30 | OR_29;
  assign input_31 = keyinput_31 ^ ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign AND_31 = input_31 & OR_30;
  assign input_32 = keyinput_32 ^ P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign OR_32 = input_32 | AND_31;
  assign input_33 = keyinput_33 ^ P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign AND_33 = input_33 & OR_32;
  assign input_34 = keyinput_34 ^ ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign AND_34 = input_34 & AND_33;
  assign input_35 = keyinput_35 ^ ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign OR_35 = input_35 | AND_34;
  assign input_36 = keyinput_36 ^ ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign AND_36 = input_36 & OR_35;
  assign input_37 = keyinput_37 ^ P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign AND_37 = input_37 & AND_36;
  assign input_38 = keyinput_38 ^ P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign OR_38 = input_38 | AND_37;
  assign input_39 = keyinput_39 ^ ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign OR_39 = input_39 | OR_38;
  assign input_40 = keyinput_40 ^ ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign OR_40 = input_40 | OR_39;
  assign input_41 = keyinput_41 ^ P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign OR_41 = input_41 | OR_40;
  assign input_42 = keyinput_42 ^ ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign OR_42 = input_42 | OR_41;
  assign input_43 = keyinput_43 ^ P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign OR_43 = input_43 | OR_42;
  assign input_44 = keyinput_44 ^ ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign OR_44 = input_44 | OR_43;
  assign input_45 = keyinput_45 ^ P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign OR_45 = input_45 | OR_44;
  assign input_46 = keyinput_46 ^ P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign OR_46 = input_46 | OR_45;
  assign input_47 = keyinput_47 ^ ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign OR_47 = input_47 | OR_46;
  assign input_48 = keyinput_48 ^ ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign OR_48 = input_48 | OR_47;
  assign input_49 = keyinput_49 ^ ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign AND_49 = input_49 & OR_48;
  assign input_50 = keyinput_50 ^ P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign AND_50 = input_50 & AND_49;
  assign input_51 = keyinput_51 ^ P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign AND_51 = input_51 & AND_50;
  assign input_52 = keyinput_52 ^ ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign OR_52 = input_52 | AND_51;
  assign input_53 = keyinput_53 ^ P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign OR_53 = input_53 | OR_52;
  assign input_54 = keyinput_54 ^ P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign AND_54 = input_54 & OR_53;
  assign input_55 = keyinput_55 ^ ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign OR_55 = input_55 | AND_54;
  assign input_56 = keyinput_56 ^ P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign AND_56 = input_56 & OR_55;
  assign input_57 = keyinput_57 ^ ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign OR_57 = input_57 | AND_56;
  assign input_58 = keyinput_58 ^ ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign AND_58 = input_58 & OR_57;
  assign input_59 = keyinput_59 ^ ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign AND_59 = input_59 & AND_58;
  assign input_60 = keyinput_60 ^ P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign AND_60 = input_60 & AND_59;
  assign input_61 = keyinput_61 ^ ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign AND_61 = input_61 & AND_60;
  assign input_62 = keyinput_62 ^ P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign OR_62 = input_62 | AND_61;
  assign input_63 = keyinput_63 ^ P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign AND_63 = input_63 & OR_62;
  assign input_64 = keyinput_64 ^ ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign AND_64 = input_64 & AND_63;
  assign input_65 = keyinput_65 ^ ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign OR_65 = input_65 | AND_64;
  assign input_66 = keyinput_66 ^ P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign AND_66 = input_66 & OR_65;
  assign input_67 = keyinput_67 ^ P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign AND_67 = input_67 & AND_66;
  assign input_68 = keyinput_68 ^ P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign AND_68 = input_68 & AND_67;
  assign input_69 = keyinput_69 ^ ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign AND_69 = input_69 & AND_68;
  assign input_70 = keyinput_70 ^ P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign AND_70 = input_70 & AND_69;
  assign input_71 = keyinput_71 ^ P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign OR_71 = input_71 | AND_70;
  assign input_72 = keyinput_72 ^ ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign AND_72 = input_72 & OR_71;
  assign input_73 = keyinput_73 ^ ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign OR_73 = input_73 | AND_72;
  assign input_74 = keyinput_74 ^ ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign OR_74 = input_74 | OR_73;
  assign input_75 = keyinput_75 ^ ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign AND_75 = input_75 & OR_74;
  assign input_76 = keyinput_76 ^ ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign OR_76 = input_76 | AND_75;
  assign input_77 = keyinput_77 ^ ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign AND_77 = input_77 & OR_76;
  assign input_78 = keyinput_78 ^ ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign AND_78 = input_78 & AND_77;
  assign input_79 = keyinput_79 ^ ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign AND_79 = input_79 & AND_78;
  assign input_80 = keyinput_80 ^ READY12_REG_SCAN_IN;
  assign input_81 = keyinput_81 ^ READY21_REG_SCAN_IN;
  assign AND_81 = input_80 & input_81;
  assign input_82 = keyinput_82 ^ P2_STATE_REG_2__SCAN_IN;
  assign OR_82 = input_82 | AND_81;
  assign input_83 = keyinput_83 ^ ~P2_STATE_REG_1__SCAN_IN;
  assign OR_83 = input_83 | OR_82;
  assign input_84 = keyinput_84 ^ P2_STATE_REG_0__SCAN_IN;
  assign AND_84 = input_84 & OR_83;
  assign input_85 = keyinput_85 ^ ~P2_STATE2_REG_3__SCAN_IN;
  assign OR_85 = input_85 | AND_84;
  assign input_86 = keyinput_86 ^ P2_STATE2_REG_2__SCAN_IN;
  assign OR_86 = input_86 | OR_85;
  assign input_87 = keyinput_87 ^ P2_STATE2_REG_1__SCAN_IN;
  assign AND_87 = input_87 & OR_86;
  assign input_88 = keyinput_88 ^ ~P2_STATE2_REG_0__SCAN_IN;
  assign OR_88 = input_88 | AND_87;
  assign input_89 = keyinput_89 ^ ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign AND_89 = input_89 & OR_88;
  assign input_90 = keyinput_90 ^ ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign OR_90 = input_90 | AND_89;
  assign input_91 = keyinput_91 ^ ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign OR_91 = input_91 | OR_90;
  assign input_92 = keyinput_92 ^ P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign AND_92 = input_92 & OR_91;
  assign input_93 = keyinput_93 ^ ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign AND_93 = input_93 & AND_92;
  assign input_94 = keyinput_94 ^ P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign AND_94 = input_94 & AND_93;
  assign input_95 = keyinput_95 ^ P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign AND_95 = input_95 & AND_94;
  assign input_96 = keyinput_96 ^ P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign AND_96 = input_96 & AND_95;
  assign input_97 = keyinput_97 ^ P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign AND_97 = input_97 & AND_96;
  assign input_98 = keyinput_98 ^ P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign OR_98 = input_98 | AND_97;
  assign input_99 = keyinput_99 ^ ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign AND_99 = input_99 & OR_98;
  assign input_100 = keyinput_100 ^ P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign AND_100 = input_100 & AND_99;
  assign input_101 = keyinput_101 ^ ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign AND_101 = input_101 & AND_100;
  assign input_102 = keyinput_102 ^ ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign AND_102 = input_102 & AND_101;
  assign input_103 = keyinput_103 ^ P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign OR_103 = input_103 | AND_102;
  assign input_104 = keyinput_104 ^ ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign AND_104 = input_104 & OR_103;
  assign input_105 = keyinput_105 ^ P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign OR_105 = input_105 | AND_104;
  assign input_106 = keyinput_106 ^ P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign OR_106 = input_106 | OR_105;
  assign input_107 = keyinput_107 ^ ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign AND_107 = input_107 & OR_106;
  assign input_108 = keyinput_108 ^ ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign OR_108 = input_108 | AND_107;
  assign input_109 = keyinput_109 ^ P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign OR_109 = input_109 | OR_108;
  assign input_110 = keyinput_110 ^ P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign OR_110 = input_110 | OR_109;
  assign input_111 = keyinput_111 ^ P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign AND_111 = input_111 & OR_110;
  assign input_112 = keyinput_112 ^ ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign OR_112 = input_112 | AND_111;
  assign input_113 = keyinput_113 ^ P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign AND_113 = input_113 & OR_112;
  assign input_114 = keyinput_114 ^ ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign AND_114 = input_114 & AND_113;
  assign input_115 = keyinput_115 ^ ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign OR_115 = input_115 | AND_114;
  assign input_116 = keyinput_116 ^ ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign AND_116 = input_116 & OR_115;
  assign input_117 = keyinput_117 ^ P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign AND_117 = input_117 & AND_116;
  assign input_118 = keyinput_118 ^ ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign OR_118 = input_118 | AND_117;
  assign input_119 = keyinput_119 ^ P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign OR_119 = input_119 | OR_118;
  assign input_120 = keyinput_120 ^ P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign OR_120 = input_120 | OR_119;
  assign input_121 = keyinput_121 ^ P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign OR_121 = input_121 | OR_120;
  assign input_122 = keyinput_122 ^ ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign OR_122 = input_122 | OR_121;
  assign input_123 = keyinput_123 ^ ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign OR_123 = input_123 | OR_122;
  assign input_124 = keyinput_124 ^ P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign OR_124 = input_124 | OR_123;
  assign input_125 = keyinput_125 ^ ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign OR_125 = input_125 | OR_124;
  assign input_126 = keyinput_126 ^ P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign OR_126 = input_126 | OR_125;
  assign input_127 = keyinput_127 ^ ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign OR_127 = input_127 | OR_126;
  assign input_128 = keyinput_128 ^ ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign OR_128 = input_128 | OR_127;
  assign input_129 = keyinput_129 ^ P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign AND_129 = input_129 & OR_128;
  assign input_130 = keyinput_130 ^ ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign AND_130 = input_130 & AND_129;
  assign input_131 = keyinput_131 ^ P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign AND_131 = input_131 & AND_130;
  assign input_132 = keyinput_132 ^ ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign OR_132 = input_132 | AND_131;
  assign input_133 = keyinput_133 ^ P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign OR_133 = input_133 | OR_132;
  assign input_134 = keyinput_134 ^ ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign AND_134 = input_134 & OR_133;
  assign input_135 = keyinput_135 ^ P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign OR_135 = input_135 | AND_134;
  assign input_136 = keyinput_136 ^ P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign AND_136 = input_136 & OR_135;
  assign input_137 = keyinput_137 ^ P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign OR_137 = input_137 | AND_136;
  assign input_138 = keyinput_138 ^ P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign AND_138 = input_138 & OR_137;
  assign input_139 = keyinput_139 ^ P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign AND_139 = input_139 & AND_138;
  assign input_140 = keyinput_140 ^ P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign AND_140 = input_140 & AND_139;
  assign input_141 = keyinput_141 ^ ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign AND_141 = input_141 & AND_140;
  assign input_142 = keyinput_142 ^ P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign OR_142 = input_142 | AND_141;
  assign input_143 = keyinput_143 ^ P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign AND_143 = input_143 & OR_142;
  assign input_144 = keyinput_144 ^ P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign AND_144 = input_144 & AND_143;
  assign input_145 = keyinput_145 ^ ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign OR_145 = input_145 | AND_144;
  assign input_146 = keyinput_146 ^ ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign AND_146 = input_146 & OR_145;
  assign input_147 = keyinput_147 ^ P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign AND_147 = input_147 & AND_146;
  assign input_148 = keyinput_148 ^ ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign AND_148 = input_148 & AND_147;
  assign input_149 = keyinput_149 ^ P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign AND_149 = input_149 & AND_148;
  assign input_150 = keyinput_150 ^ P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign AND_150 = input_150 & AND_149;
  assign input_151 = keyinput_151 ^ P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign OR_151 = input_151 | AND_150;
  assign input_152 = keyinput_152 ^ ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign AND_152 = input_152 & OR_151;
  assign input_153 = keyinput_153 ^ ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign OR_153 = input_153 | AND_152;
  assign input_154 = keyinput_154 ^ P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign OR_154 = input_154 | OR_153;
  assign input_155 = keyinput_155 ^ ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign AND_155 = input_155 & OR_154;
  assign input_156 = keyinput_156 ^ ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign OR_156 = input_156 | AND_155;
  assign input_157 = keyinput_157 ^ P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign AND_157 = input_157 & OR_156;
  assign input_158 = keyinput_158 ^ P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign AND_158 = input_158 & AND_157;
  assign input_159 = keyinput_159 ^ ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign AND_159 = input_159 & AND_158;
  assign AND_159_INV = ~AND_159;
  assign CASOP = AND_79 & AND_159_INV;
  assign P2_U3015 = P2_U3015_Lock ^ CASOP;
endmodule


